-------------------------------------------------------------------------------------------------------------
-- Extender
-- This unit recieves as input the immediate filed in the instruction(15-0). Depending on the value of the
-- control signal Unsigned_value it performs and unsigned sing-extension or a signed sign-extension(in two's
-- complement. The block is fully combinational.
-------------------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use work.globals.all;


-------------------------------------------------------------------------------------------------------------
-------------------------------------------------------------------------------------------------------------

entity extender is
	port (
		-- INPUTS
		immediate        : in std_logic_vector(15 downto 0);	  -- immediate filed (instruction 15 -0)
		unsigned_value   : in std_logic;			                  -- control signal generated by the CU
		-- OUTPUTS
		extended         : out std_logic_vector(31 downto 0)	  -- extended value
		);
end extender;


-------------------------------------------------------------------------------------------------------------
-------------------------------------------------------------------------------------------------------------

architecture behavioral of extender is

begin

	--------------------------------------------------
	-- Extend Process
	-- Type: Combinational
	-- Implemnents the
	-- sign-extensionl
	-- logic
	-----------------------i--------------------------
	extend_process:process(immediate, unsigned_value)
	begin
		if (unsigned_value = '1') then

			extended <= "0000000000000000" & immediate;

		else
			if (immediate(15) = '1') then

				extended(31 downto 16) <= (others => '1');
				extended(15 downto 0)  <= immediate;

			else

				extended(31 downto 16) <= (others => '0');
				extended(15 downto 0)  <= immediate;

			end if;
		end if;
	end process;

end behavioral;
