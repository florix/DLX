
module DLX ( clk, rst, iram_data, Data_out_fromRAM, addr_to_iram, read_op, 
        write_op, nibble, write_byte, Address_toRAM, Data_in );
  input [31:0] iram_data;
  input [31:0] Data_out_fromRAM;
  output [31:0] addr_to_iram;
  output [1:0] nibble;
  output [31:0] Address_toRAM;
  output [31:0] Data_in;
  input clk, rst;
  output read_op, write_op, write_byte;
  wire   addr_to_iram_29, addr_to_iram_28, addr_to_iram_27, addr_to_iram_26,
         addr_to_iram_25, addr_to_iram_24, addr_to_iram_23, addr_to_iram_22,
         addr_to_iram_21, addr_to_iram_20, addr_to_iram_19, addr_to_iram_18,
         addr_to_iram_17, addr_to_iram_16, addr_to_iram_15, addr_to_iram_14,
         addr_to_iram_13, addr_to_iram_12, addr_to_iram_11, addr_to_iram_10,
         addr_to_iram_9, addr_to_iram_8, addr_to_iram_7, addr_to_iram_6,
         addr_to_iram_5, addr_to_iram_4, addr_to_iram_3, addr_to_iram_2,
         addr_to_iram_1, addr_to_iram_0, write_byte_snps_wire, n9566, n8527,
         n8528, n8529, \u_DataPath/reg_write_i , \u_DataPath/jump_i ,
         \u_DataPath/u_fetch/pc1/N3 , \u_DataPath/u_ifidreg/N61 ,
         \u_DataPath/u_ifidreg/N59 , \u_DataPath/u_ifidreg/N57 ,
         \u_DataPath/u_decode_unit/reg_file0/N154 ,
         \u_DataPath/u_decode_unit/reg_file0/N153 ,
         \u_DataPath/u_decode_unit/reg_file0/N152 ,
         \u_DataPath/u_decode_unit/reg_file0/N151 ,
         \u_DataPath/u_decode_unit/reg_file0/N150 ,
         \u_DataPath/u_decode_unit/reg_file0/N149 ,
         \u_DataPath/u_decode_unit/reg_file0/N148 ,
         \u_DataPath/u_decode_unit/reg_file0/N147 ,
         \u_DataPath/u_decode_unit/reg_file0/N146 ,
         \u_DataPath/u_decode_unit/reg_file0/N145 ,
         \u_DataPath/u_decode_unit/reg_file0/N144 ,
         \u_DataPath/u_decode_unit/reg_file0/N143 ,
         \u_DataPath/u_decode_unit/reg_file0/N142 ,
         \u_DataPath/u_decode_unit/reg_file0/N141 ,
         \u_DataPath/u_decode_unit/reg_file0/N140 ,
         \u_DataPath/u_decode_unit/reg_file0/N139 ,
         \u_DataPath/u_decode_unit/reg_file0/N138 ,
         \u_DataPath/u_decode_unit/reg_file0/N137 ,
         \u_DataPath/u_decode_unit/reg_file0/N136 ,
         \u_DataPath/u_decode_unit/reg_file0/N135 ,
         \u_DataPath/u_decode_unit/reg_file0/N134 ,
         \u_DataPath/u_decode_unit/reg_file0/N133 ,
         \u_DataPath/u_decode_unit/reg_file0/N132 ,
         \u_DataPath/u_decode_unit/reg_file0/N131 ,
         \u_DataPath/u_decode_unit/reg_file0/N130 ,
         \u_DataPath/u_decode_unit/reg_file0/N129 ,
         \u_DataPath/u_decode_unit/reg_file0/N128 ,
         \u_DataPath/u_decode_unit/reg_file0/N127 ,
         \u_DataPath/u_decode_unit/reg_file0/N126 ,
         \u_DataPath/u_decode_unit/reg_file0/N125 ,
         \u_DataPath/u_decode_unit/reg_file0/N92 ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][0] ,
         \u_DataPath/u_idexreg/N16 , \u_DataPath/u_idexreg/N15 ,
         \u_DataPath/u_idexreg/N13 , \u_DataPath/u_idexreg/N12 ,
         \u_DataPath/u_idexreg/N10 , \u_DataPath/u_execute/ovf_i ,
         \u_DataPath/u_execute/A_inALU_i[26] ,
         \u_DataPath/u_execute/EXALU/N811 , \u_DataPath/u_execute/EXALU/N810 ,
         \u_DataPath/u_memwbreg/N74 , \u_DataPath/u_memwbreg/N73 ,
         \u_DataPath/u_memwbreg/N72 , \u_DataPath/u_memwbreg/N71 ,
         \u_DataPath/u_memwbreg/N70 , \u_DataPath/u_memwbreg/N45 , net3007,
         n1885, \lte_x_57/B[30] , \lte_x_57/B[29] , \lte_x_57/B[28] ,
         \lte_x_57/B[25] , \lte_x_57/B[15] , \lte_x_57/B[14] ,
         \lte_x_57/B[11] , \lte_x_57/B[10] , \lte_x_57/B[7] , \lte_x_57/B[6] ,
         \lte_x_57/B[4] , \lte_x_57/B[3] , \lte_x_57/B[2] , \sub_x_51/A[27] ,
         \sub_x_51/A[22] , \sub_x_51/A[21] , \sub_x_51/A[20] ,
         \sub_x_51/A[18] , \sub_x_51/A[16] , \sub_x_51/A[13] , \sub_x_51/A[8] ,
         \sub_x_51/A[5] , \add_x_50/A[23] , \add_x_50/A[19] , n2710, n2712,
         n2720, n2770, n2772, n2773, n2774, n2776, n2778, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3056, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3450, n3451,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3509, n3511, n3513, n3515, n3517,
         n3519, n3521, n3523, n3525, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3557, n3559, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3782, n3783, n3784, n3785, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
         n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
         n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
         n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4220,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
         n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
         n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
         n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
         n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
         n7647, n7648, n7649, n7650, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7672, n7673, n7674, n7675, n7676, n7677, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
         n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
         n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
         n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
         n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
         n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
         n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
         n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
         n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
         n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493,
         n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
         n8504, n8506, n8508, n8510, n8512, n8513, n8515, n8522, n8523, n8524,
         n8525, n8526, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
         n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
         n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687,
         n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
         n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
         n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
         n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
         n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
         n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
         n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
         n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
         n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
         n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
         n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
         n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
         n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
         n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
         n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
         n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
         n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
         n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
         n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
         n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
         n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
         n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
         n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
         n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
         n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
         n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
         n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
         n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
         n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407,
         n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417,
         n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
         n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
         n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
         n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
         n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467,
         n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477,
         n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487,
         n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497,
         n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507,
         n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
         n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
         n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9553, n9554, n9555, n9556, n9557, n9564, n9565;
  wire   [31:0] addr_to_iram;
  wire   [5:0] opcode_i;
  wire   [4:0] \u_DataPath/regfile_addr_out_towb_i ;
  wire   [31:0] \u_DataPath/from_alu_data_out_i ;
  wire   [31:0] \u_DataPath/from_mem_data_out_i ;
  wire   [4:0] \u_DataPath/RFaddr_out_memwb_i ;
  wire   [31:0] \u_DataPath/dataOut_exe_i ;
  wire   [2:0] \u_DataPath/cw_memwb_i ;
  wire   [31:0] \u_DataPath/mem_writedata_out_i ;
  wire   [10:0] \u_DataPath/cw_tomem_i ;
  wire   [31:0] \u_DataPath/toPC2_i ;
  wire   [10:0] \u_DataPath/cw_exmem_i ;
  wire   [4:0] \u_DataPath/rs_ex_i ;
  wire   [31:0] \u_DataPath/data_read_ex_2_i ;
  wire   [31:0] \u_DataPath/data_read_ex_1_i ;
  wire   [31:0] \u_DataPath/pc_4_to_ex_i ;
  wire   [21:0] \u_DataPath/cw_to_ex_i ;
  wire   [31:0] \u_DataPath/immediate_ext_dec_i ;
  wire   [31:0] \u_DataPath/pc4_to_idexreg_i ;
  wire   [31:0] \u_DataPath/jaddr_i ;
  wire   [4:0] \u_DataPath/idex_rt_i ;
  wire   [31:0] \u_DataPath/pc_4_i ;
  wire   [31:0] \u_DataPath/branch_target_i ;
  wire   [31:0] \u_DataPath/jump_address_i ;
  wire   [1:0] \u_DataPath/u_decode_unit/hdu_0/current_state ;
  wire   [31:0] \u_DataPath/u_execute/psw_status_i ;
  wire   [31:0] \u_DataPath/u_execute/link_value_i ;
  wire   [31:0] \u_DataPath/u_execute/resAdd1_i ;
  assign Address_toRAM[30] = 1'b0;
  assign Address_toRAM[31] = 1'b0;
  assign addr_to_iram[30] = 1'b0;
  assign addr_to_iram[31] = 1'b0;
  assign Address_toRAM[8] = n3441;
  assign Address_toRAM[12] = n3442;
  assign Data_in[31] = n3445;
  assign Data_in[28] = n3446;
  assign Data_in[30] = n3447;
  assign Data_in[29] = n3448;
  assign Data_in[9] = n3451;
  assign Address_toRAM[4] = n3506;
  assign Data_in[23] = n3507;
  assign Data_in[13] = n3509;
  assign Data_in[12] = n3511;
  assign Data_in[10] = n3513;
  assign Data_in[11] = n3515;
  assign Data_in[21] = n3517;
  assign Data_in[19] = n3519;
  assign Data_in[20] = n3521;
  assign Data_in[22] = n3523;
  assign Data_in[17] = n3525;
  assign Address_toRAM[11] = n3533;
  assign Address_toRAM[24] = n3535;
  assign Address_toRAM[6] = n3554;
  assign Data_in[14] = n3555;
  assign Data_in[18] = n3557;
  assign Data_in[15] = n3559;
  assign addr_to_iram[17] = n9506;
  assign addr_to_iram[22] = n9507;
  assign addr_to_iram[11] = n9508;
  assign addr_to_iram[13] = n9509;
  assign addr_to_iram[12] = n9510;
  assign addr_to_iram[16] = n9511;
  assign addr_to_iram[7] = n9512;
  assign addr_to_iram[9] = n9513;
  assign addr_to_iram[23] = n9514;
  assign addr_to_iram[10] = n9515;
  assign addr_to_iram[6] = n9516;
  assign addr_to_iram[8] = n9517;
  assign addr_to_iram[5] = n9518;
  assign addr_to_iram[4] = n9519;
  assign addr_to_iram[3] = n9520;
  assign addr_to_iram[2] = n9521;
  assign addr_to_iram[0] = n9522;
  assign addr_to_iram[1] = n9523;
  assign addr_to_iram[18] = n9524;
  assign addr_to_iram[20] = n9525;
  assign addr_to_iram[24] = n9526;
  assign addr_to_iram[14] = n9527;
  assign addr_to_iram[19] = n9528;
  assign addr_to_iram[21] = n9529;
  assign addr_to_iram[25] = n9530;
  assign addr_to_iram[15] = n9531;
  assign addr_to_iram[26] = n9532;
  assign addr_to_iram[27] = n9533;
  assign addr_to_iram[28] = n9534;
  assign addr_to_iram[29] = n9535;
  assign write_byte = n9536;

  HS65_LH_CNIVX3 U87 ( .A(rst), .Z(n1885) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7743), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7724), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7916), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7796), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7803), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7928), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7751), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7873), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7817), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7789), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7921), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7887), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7823), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7880), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7768), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7838), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7908), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7901), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7830), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7775), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7757), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7761), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7809), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7845), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7852), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7730), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7925), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7894), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7782), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7866), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7859), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7737), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7722), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7722), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7795), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7795), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7802), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7802), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7926), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7926), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7750), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7750), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7872), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7872), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7816), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7816), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7788), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7788), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7886), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7886), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7879), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7879), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7767), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7767), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7837), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7837), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7907), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7907), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7900), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7900), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7774), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7774), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7756), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7756), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7760), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7760), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7844), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7844), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7851), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7851), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7729), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7729), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7923), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7923), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7893), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7893), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7781), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7781), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7865), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7865), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7858), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7858), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7736), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7736), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7722), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7722), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7796), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7795), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7803), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7802), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7926), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7926), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7751), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7750), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7873), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7872), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7817), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7816), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7789), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7788), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7887), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7886), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7880), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7879), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7768), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7767), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7838), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7837), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7908), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7907), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7901), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7900), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7775), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7774), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7757), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7756), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7761), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7760), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7845), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7844), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7852), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7851), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7730), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7729), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7923), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7923), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7894), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7893), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7782), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7781), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7866), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7865), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7859), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7858), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7737), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7736), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7723), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7915), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7796), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7803), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7927), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7751), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7873), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7817), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7789), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7921), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7887), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7880), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7768), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7838), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7908), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7901), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7775), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7757), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7761), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7845), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7852), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7730), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7924), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7894), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7782), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7866), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7859), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7737), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7722), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7914), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7795), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7802), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7927), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7750), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7872), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7816), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7788), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7920), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7886), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7879), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7767), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7837), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7907), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7900), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7774), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7756), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7760), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7844), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7851), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7729), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7923), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7893), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7781), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7865), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7858), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7736), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][27] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_execute/EXALU/ovf_reg  ( .G(
        \u_DataPath/u_execute/EXALU/N810 ), .D(
        \u_DataPath/u_execute/EXALU/N811 ), .Q(\u_DataPath/u_execute/ovf_i )
         );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7744), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7723), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7915), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7795), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7802), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7927), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7750), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7872), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7816), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7788), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7920), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7886), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7824), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7879), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7767), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7837), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7907), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7900), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7831), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7774), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7756), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7760), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7810), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7844), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7851), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7729), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7924), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7893), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7781), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7865), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7858), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7736), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7743), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7916), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7921), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7823), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7830), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7809), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7745), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7744), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7914), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7914), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7920), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7920), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7824), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7825), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7831), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7832), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7810), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7811), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7744), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7824), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7831), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7810), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7745), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7722), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7914), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7795), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7802), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7926), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7750), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7872), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7816), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7788), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7920), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7886), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7825), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7879), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7767), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7837), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7907), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7900), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7832), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7774), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7756), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7760), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7811), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7844), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7851), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7729), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7923), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7893), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7781), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7865), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7858), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7736), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7745), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7722), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7914), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7796), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7803), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7926), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7751), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7873), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7817), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7789), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7921), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7887), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7825), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7880), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7768), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7838), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7908), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7901), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7832), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7775), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7757), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7761), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7811), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7845), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7852), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7730), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7923), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7894), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7782), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7866), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7859), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7737), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7745), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7744), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7723), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7915), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7795), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7802), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7927), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7750), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7872), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7816), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7788), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7920), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7886), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7824), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7825), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7879), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7767), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7837), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7907), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7900), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7831), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7832), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7774), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7756), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7760), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7810), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7811), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7844), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7851), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7729), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7924), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7893), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7781), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7865), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7858), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7736), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7744), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7723), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7914), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7914), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7915), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7797), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7804), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7927), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7752), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7874), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7818), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7790), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7922), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7888), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7824), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7881), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7769), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7839), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7909), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7902), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7831), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7776), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7758), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7762), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7810), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7846), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7853), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7731), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7924), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7895), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7783), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7867), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7860), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7738), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7744), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7745), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7921), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7920), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7825), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7824), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7832), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7831), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7811), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7810), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7744), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7744), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7745), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7745), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7722), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7722), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7723), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7914), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7914), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7915), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7795), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7795), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7795), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7802), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7802), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7802), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7926), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7926), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7927), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7750), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7750), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7750), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7872), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7872), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7872), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7816), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7816), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7816), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7788), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7788), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7788), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7920), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7920), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7920), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7886), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7886), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7886), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7825), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7824), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7825), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7824), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7879), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7879), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7879), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7767), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7767), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7767), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7837), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7837), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7837), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7907), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7907), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7907), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7900), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7900), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7900), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7832), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7831), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7832), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7831), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7774), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7774), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7774), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7756), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7756), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7756), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7760), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7760), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7760), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7811), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7810), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7811), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7810), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7844), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7844), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7844), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7851), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7851), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7851), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7729), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7729), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7729), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7923), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7923), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7924), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7893), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7893), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7893), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7781), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7781), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7781), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7865), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7865), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7865), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7858), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7858), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7858), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7736), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7736), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7736), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7744), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7722), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7914), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7795), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7802), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7926), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7750), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7872), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7816), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7788), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7920), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7886), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7824), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7879), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7767), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7837), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7907), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7900), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7831), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7774), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7756), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7760), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7810), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7844), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7851), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7729), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7923), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7893), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7781), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7865), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7858), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7736), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7745), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7722), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7914), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7796), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7803), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7926), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7751), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7873), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7817), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7789), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7921), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7887), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7825), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7880), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7768), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7838), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7908), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7901), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7832), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7775), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7757), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7761), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7811), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7845), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7852), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7730), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7923), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7894), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7782), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7866), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7859), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7737), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7744), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7722), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7914), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7795), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7802), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7926), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7750), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7872), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7816), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7788), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7920), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7886), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7824), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7879), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7767), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7837), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7907), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7900), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7831), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7774), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7756), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7760), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7810), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7844), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7851), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7729), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7923), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7893), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7781), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7865), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7858), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7736), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7743), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7724), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7723), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7723), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7915), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7915), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7796), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7797), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7796), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7803), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7804), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7803), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7928), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7926), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7927), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7751), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7752), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7751), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7873), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7874), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7873), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7817), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7818), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7817), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7789), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7790), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7789), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7922), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7921), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7887), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7888), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7887), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7823), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7880), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7881), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7880), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7768), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7769), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7768), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7838), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7839), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7838), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7908), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7909), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7908), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7901), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7902), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7901), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7830), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7775), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7776), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7775), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7757), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7758), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7757), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7761), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7762), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7761), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7809), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7845), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7846), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7845), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7852), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7853), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7852), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7730), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7731), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7730), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7925), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7924), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7924), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7894), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7895), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7894), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7782), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7783), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7782), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7866), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7867), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7866), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7859), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7860), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7859), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7737), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7738), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7737), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][27] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][31]  ( 
        .G(rst), .D(n7743), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][31] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][0]  ( 
        .G(rst), .D(n7723), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][0] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][1]  ( 
        .G(rst), .D(n7915), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][1] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][6]  ( 
        .G(rst), .D(n7796), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][6] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][18]  ( 
        .G(rst), .D(n7803), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][18] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][2]  ( 
        .G(rst), .D(n7927), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][2] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][17]  ( 
        .G(rst), .D(n7751), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][17] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][16]  ( 
        .G(rst), .D(n7873), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][16] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][20]  ( 
        .G(rst), .D(n7817), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][20] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][8]  ( 
        .G(rst), .D(n7789), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][8] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][4]  ( 
        .G(rst), .D(n7921), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][4] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][22]  ( 
        .G(rst), .D(n7887), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][22] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][28]  ( 
        .G(rst), .D(n7823), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][28] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][24]  ( 
        .G(rst), .D(n7880), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][24] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][9]  ( 
        .G(rst), .D(n7768), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][9] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][25]  ( 
        .G(rst), .D(n7838), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][25] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][5]  ( 
        .G(rst), .D(n7908), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][5] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][21]  ( 
        .G(rst), .D(n7901), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][21] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][29]  ( 
        .G(rst), .D(n7830), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][29] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][13]  ( 
        .G(rst), .D(n7775), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][13] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][7]  ( 
        .G(rst), .D(n7757), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][7] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][12]  ( 
        .G(rst), .D(n7761), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][12] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][30]  ( 
        .G(rst), .D(n7809), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][30] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][23]  ( 
        .G(rst), .D(n7845), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][23] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][26]  ( 
        .G(rst), .D(n7852), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][26] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][10]  ( 
        .G(rst), .D(n7730), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][10] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][3]  ( 
        .G(rst), .D(n7924), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][3] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][19]  ( 
        .G(rst), .D(n7894), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][19] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][11]  ( 
        .G(rst), .D(n7782), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][11] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][15]  ( 
        .G(rst), .D(n7866), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][15] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][14]  ( 
        .G(rst), .D(n7859), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][14] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][27]  ( 
        .G(rst), .D(n7737), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][27] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7743), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][31] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7724), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][0] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7916), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][1] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7797), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][6] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7804), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][18] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7928), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][2] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7752), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][17] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7874), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][16] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7818), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][20] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7790), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][8] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7922), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][4] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7888), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][22] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7823), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][28] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7881), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][24] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7769), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][9] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7839), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][25] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7909), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][5] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7902), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][21] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7830), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][29] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7776), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][13] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7758), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][7] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7762), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][12] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7809), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][30] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7846), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][23] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7853), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][26] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7731), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][10] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7925), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][3] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7895), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][19] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7783), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][11] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7867), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][15] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7860), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][14] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7738), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][27] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7744), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][31] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7724), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][0] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7916), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][1] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7797), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][6] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7804), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][18] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7928), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][2] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7752), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][17] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7874), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][16] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7818), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][20] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7790), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][8] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7922), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][4] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7888), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][22] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7824), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][28] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7881), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][24] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7769), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][9] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7839), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][25] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7909), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][5] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7902), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][21] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7831), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][29] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7776), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][13] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7758), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][7] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7762), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][12] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7810), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][30] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7846), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][23] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7853), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][26] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7731), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][10] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7925), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][3] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7895), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][19] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7783), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][11] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7867), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][15] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7860), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][14] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7738), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][27] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7744), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][31] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7824), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][28] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7831), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][29] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7810), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][30] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7743), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][31] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7921), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][4] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7823), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][28] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7830), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][29] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7809), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][30] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7743), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][31] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7723), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][0] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7916), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][1] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7915), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][1] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7797), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][6] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7804), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][18] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7927), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][2] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7752), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][17] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7874), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][16] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7818), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][20] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7790), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][8] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7922), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][4] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7888), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][22] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7823), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][28] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7881), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][24] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7769), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][9] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7839), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][25] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7909), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][5] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7902), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][21] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7830), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][29] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7776), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][13] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7758), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][7] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7762), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][12] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7809), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][30] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7846), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][23] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7853), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][26] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7731), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][10] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7924), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][3] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7895), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][19] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7783), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][11] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7867), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][15] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7860), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][14] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7738), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][27] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7915), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][1] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7743), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][31] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7921), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][4] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7823), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][28] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7830), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][29] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7809), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][30] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7743), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][31] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7743), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][31] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7723), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][0] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7915), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][1] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7796), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][6] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7803), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][18] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7927), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][2] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7751), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][17] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7873), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][16] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7817), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][20] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7789), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][8] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7922), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][4] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7921), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][4] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7887), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][22] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7823), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][28] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7823), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][28] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7880), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][24] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7768), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][9] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7838), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][25] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7908), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][5] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7901), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][21] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7830), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][29] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7830), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][29] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7775), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][13] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7757), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][7] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7761), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][12] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7809), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][30] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7809), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][30] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7845), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][23] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7852), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][26] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7730), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][10] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7924), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][3] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7894), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][19] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7782), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][11] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7866), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][15] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7859), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][14] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7737), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][27] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7916), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][1] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7724), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][0] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7916), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][1] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7797), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][6] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7804), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][18] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7928), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][2] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7752), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][17] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7874), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][16] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7818), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][20] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7790), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][8] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7922), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][4] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7888), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][22] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7881), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][24] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7769), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][9] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7839), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][25] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7909), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][5] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7902), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][21] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7776), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][13] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7758), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][7] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7762), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][12] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7846), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][23] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7853), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][26] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7731), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][10] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7925), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][3] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7895), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][19] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7783), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][11] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7867), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][15] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7860), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][14] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7738), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][27] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7723), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][0] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7796), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][6] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7803), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][18] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7927), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][2] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7751), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][17] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7873), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][16] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7817), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][20] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7789), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][8] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7887), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][22] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7880), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][24] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7768), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][9] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7838), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][25] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7908), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][5] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7901), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][21] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7775), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][13] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7757), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][7] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7761), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][12] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7845), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][23] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7852), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][26] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7730), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][10] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7924), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][3] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7894), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][19] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7782), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][11] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7866), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][15] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7859), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][14] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7737), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][27] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7743), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][31] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7724), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][0] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7724), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][0] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7916), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][1] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7796), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][6] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7796), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][6] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7803), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][18] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7803), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][18] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7928), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][2] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7928), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][2] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7751), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][17] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7751), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][17] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7873), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][16] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7873), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][16] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7817), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][20] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7817), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][20] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7789), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][8] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7789), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][8] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7921), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][4] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7887), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][22] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7887), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][22] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7823), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][28] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7880), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][24] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7880), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][24] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7768), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][9] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7768), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][9] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7838), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][25] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7838), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][25] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7908), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][5] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7908), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][5] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7901), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][21] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7901), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][21] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7830), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][29] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7775), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][13] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7775), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][13] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7757), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][7] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7757), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][7] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7761), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][12] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7761), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][12] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7809), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][30] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7845), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][23] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7845), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][23] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7852), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][26] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7852), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][26] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7730), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][10] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7730), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][10] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7925), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][3] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7925), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][3] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7894), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][19] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7894), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][19] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7782), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][11] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7782), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][11] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7866), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][15] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7866), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][15] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7859), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][14] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7859), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][14] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7737), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][27] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7737), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][27] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7724), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][0] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7797), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][6] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7804), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][18] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7928), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][2] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7752), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][17] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7874), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][16] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7818), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][20] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7790), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][8] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7888), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][22] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7881), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][24] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7769), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][9] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7839), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][25] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7909), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][5] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7902), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][21] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7776), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][13] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7758), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][7] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7762), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][12] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7846), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][23] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7853), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][26] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7731), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][10] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7925), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][3] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7895), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][19] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7783), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][11] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7867), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][15] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7860), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][14] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7738), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][27] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7743), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][31] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7723), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][0] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7915), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][1] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7797), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][6] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7804), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][18] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7927), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][2] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7752), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][17] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7874), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][16] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7818), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][20] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7790), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][8] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7922), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][4] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7888), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][22] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7823), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][28] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7881), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][24] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7769), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][9] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7839), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][25] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7909), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][5] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7902), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][21] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7830), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][29] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7776), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][13] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7758), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][7] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7762), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][12] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7809), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][30] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7846), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][23] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7853), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][26] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7731), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][10] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7924), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][3] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7895), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][19] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7783), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][11] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7867), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][15] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7860), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][14] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7738), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][27] ) );
  HS65_LH_BFX9 U3398 ( .A(n7302), .Z(n7701) );
  HS65_LH_BFX9 U3445 ( .A(n6267), .Z(n6908) );
  HS65_LH_BFX9 U3446 ( .A(n6976), .Z(n6726) );
  HS65_LH_BFX9 U3447 ( .A(n6977), .Z(n6727) );
  HS65_LH_BFX9 U3448 ( .A(n6975), .Z(n6725) );
  HS65_LH_BFX9 U3452 ( .A(n6265), .Z(n2801) );
  HS65_LH_BFX9 U3453 ( .A(n6346), .Z(n7001) );
  HS65_LH_BFX9 U3454 ( .A(n6985), .Z(n6909) );
  HS65_LH_NOR2X6 U3455 ( .A(n5963), .B(n5962), .Z(n2822) );
  HS65_LH_BFX9 U3456 ( .A(n6499), .Z(n6974) );
  HS65_LL_NOR2X6 U3460 ( .A(n5958), .B(n5952), .Z(n6113) );
  HS65_LH_NOR2AX3 U3461 ( .A(n9175), .B(n6478), .Z(n6486) );
  HS65_LH_NOR2X13 U3462 ( .A(n6184), .B(n6185), .Z(n6278) );
  HS65_LH_NOR2X6 U3463 ( .A(n6188), .B(n6187), .Z(n6348) );
  HS65_LH_AND2X4 U3465 ( .A(n9361), .B(n7307), .Z(n2849) );
  HS65_LH_NOR2X6 U3466 ( .A(n6186), .B(n6175), .Z(n6333) );
  HS65_LH_NOR2X6 U3467 ( .A(n5958), .B(n5950), .Z(n6108) );
  HS65_LH_NOR2X6 U3468 ( .A(n6182), .B(n6183), .Z(n6346) );
  HS65_LH_NOR2X6 U3469 ( .A(n5960), .B(n5963), .Z(n6131) );
  HS65_LH_NOR2X6 U3470 ( .A(n5963), .B(n5937), .Z(n6103) );
  HS65_LH_NOR2X6 U3471 ( .A(n6186), .B(n6162), .Z(n6258) );
  HS65_LH_NOR2X6 U3472 ( .A(n6182), .B(n6176), .Z(n6985) );
  HS65_LH_NOR2X6 U3473 ( .A(n6186), .B(n6176), .Z(n6338) );
  HS65_LH_NOR2X6 U3474 ( .A(n6188), .B(n6174), .Z(n6986) );
  HS65_LH_NOR2X6 U3475 ( .A(n5958), .B(n5951), .Z(n6111) );
  HS65_LH_NOR2X6 U3476 ( .A(n5958), .B(n5957), .Z(n6127) );
  HS65_LH_OR2X9 U3477 ( .A(\u_DataPath/jaddr_i [17]), .B(
        \u_DataPath/jaddr_i [16]), .Z(n5963) );
  HS65_LH_NAND2X7 U3478 ( .A(\u_DataPath/jaddr_i [16]), .B(
        \u_DataPath/jaddr_i [17]), .Z(n5958) );
  HS65_LL_AOI21X3 U3479 ( .A(n7327), .B(n4269), .C(n4268), .Z(n8350) );
  HS65_LH_NAND2X7 U3480 ( .A(n2816), .B(n6479), .Z(n6182) );
  HS65_LL_NOR2X2 U3481 ( .A(n4815), .B(n4814), .Z(n4816) );
  HS65_LH_AND2X4 U3483 ( .A(n2818), .B(\u_DataPath/jaddr_i [24]), .Z(n6163) );
  HS65_LH_AOI21X2 U3484 ( .A(n5517), .B(n4945), .C(n4387), .Z(n4388) );
  HS65_LH_AOI21X2 U3486 ( .A(n4925), .B(n4924), .C(n4923), .Z(n4939) );
  HS65_LH_AOI21X2 U3487 ( .A(n4667), .B(n4741), .C(n4666), .Z(n4668) );
  HS65_LH_AOI21X2 U3488 ( .A(n5255), .B(n5254), .C(n5253), .Z(n5256) );
  HS65_LH_IVX9 U3493 ( .A(n4305), .Z(n7325) );
  HS65_LH_OAI21X2 U3496 ( .A(n5212), .B(n5096), .C(n5214), .Z(n5099) );
  HS65_LH_AOI21X2 U3497 ( .A(n5393), .B(n5392), .C(n3960), .Z(n5237) );
  HS65_LL_AOI12X2 U3498 ( .A(n3905), .B(n4082), .C(n3904), .Z(n3906) );
  HS65_LL_NOR2AX3 U3503 ( .A(n3599), .B(n3598), .Z(n3600) );
  HS65_LH_NOR3X4 U3506 ( .A(\u_DataPath/cw_exmem_i [3]), .B(
        \u_DataPath/cw_exmem_i [6]), .C(n7210), .Z(n7211) );
  HS65_LH_IVX9 U3512 ( .A(n5196), .Z(n3204) );
  HS65_LH_IVX9 U3513 ( .A(\u_DataPath/jaddr_i [22]), .Z(n6479) );
  HS65_LH_IVX9 U3514 ( .A(n2817), .Z(n2818) );
  HS65_LH_IVX9 U3516 ( .A(n5312), .Z(n2790) );
  HS65_LH_IVX9 U3518 ( .A(\u_DataPath/jaddr_i [18]), .Z(n8016) );
  HS65_LH_AOI21X2 U3519 ( .A(n4796), .B(\lte_x_57/B[4] ), .C(n3475), .Z(n3478)
         );
  HS65_LL_NAND2AX4 U3520 ( .A(n4225), .B(n4750), .Z(n4150) );
  HS65_LH_BFX9 U3522 ( .A(\u_DataPath/jaddr_i [19]), .Z(n2804) );
  HS65_LL_NAND2X7 U3524 ( .A(n4433), .B(n4673), .Z(n5481) );
  HS65_LH_AOI21X2 U3526 ( .A(n5802), .B(n5741), .C(n5740), .Z(n5776) );
  HS65_LH_AOI21X2 U3527 ( .A(n5848), .B(n5737), .C(n5736), .Z(n5738) );
  HS65_LH_IVX18 U3530 ( .A(n3379), .Z(n5506) );
  HS65_LH_NOR2X6 U3533 ( .A(n4270), .B(n4023), .Z(n4238) );
  HS65_LH_IVX9 U3535 ( .A(n5529), .Z(n5192) );
  HS65_LH_AOI21X2 U3537 ( .A(n8736), .B(n9060), .C(n8722), .Z(n5646) );
  HS65_LH_AOI21X2 U3538 ( .A(n8891), .B(n8711), .C(n9296), .Z(n5633) );
  HS65_LH_AOI21X2 U3539 ( .A(n5647), .B(n5536), .C(n5535), .Z(n5537) );
  HS65_LH_IVX9 U3541 ( .A(\lte_x_57/B[28] ), .Z(n4901) );
  HS65_LH_IVX9 U3545 ( .A(n3039), .Z(n4032) );
  HS65_LH_IVX9 U3546 ( .A(\lte_x_57/B[10] ), .Z(n5385) );
  HS65_LH_IVX9 U3550 ( .A(n2774), .Z(n2780) );
  HS65_LH_AO112X9 U3552 ( .A(n8692), .B(n2712), .C(n3159), .D(n3158), .Z(n3160) );
  HS65_LH_NOR2X6 U3553 ( .A(n3173), .B(n2794), .Z(n8433) );
  HS65_LH_NAND2AX7 U3554 ( .A(n2922), .B(n2921), .Z(n4877) );
  HS65_LH_AOI21X2 U3557 ( .A(n9425), .B(n8733), .C(n8875), .Z(n7654) );
  HS65_LH_AOI21X2 U3558 ( .A(n2710), .B(n8695), .C(n3121), .Z(n3122) );
  HS65_LH_AOI21X2 U3559 ( .A(n8690), .B(n2710), .C(n3179), .Z(n3182) );
  HS65_LH_MUXI21X2 U3560 ( .D0(\u_DataPath/from_alu_data_out_i [31]), .D1(
        \u_DataPath/from_mem_data_out_i [31]), .S0(n3235), .Z(n8040) );
  HS65_LH_NOR2AX3 U3561 ( .A(\u_DataPath/from_alu_data_out_i [28]), .B(n3148), 
        .Z(n3115) );
  HS65_LH_CNIVX3 U3563 ( .A(n8160), .Z(n2785) );
  HS65_LL_IVX9 U3573 ( .A(n3048), .Z(n2781) );
  HS65_LH_AND2X4 U3574 ( .A(\u_DataPath/cw_memwb_i [2]), .B(n2907), .Z(n2912)
         );
  HS65_LLS_XOR2X3 U3575 ( .A(\u_DataPath/RFaddr_out_memwb_i [3]), .B(
        \u_DataPath/idex_rt_i [3]), .Z(n2770) );
  HS65_LL_NOR2AX25 U3586 ( .A(n9106), .B(n3568), .Z(Data_in[27]) );
  HS65_LL_NOR2AX25 U3591 ( .A(\u_DataPath/dataOut_exe_i [17]), .B(n3567), .Z(
        Address_toRAM[15]) );
  HS65_LH_NAND2X2 U3624 ( .A(\u_DataPath/pc_4_to_ex_i [9]), .B(
        \u_DataPath/pc_4_to_ex_i [8]), .Z(n6751) );
  HS65_LL_NAND2X2 U3626 ( .A(\add_x_50/A[23] ), .B(n5252), .Z(n4720) );
  HS65_LLS_XNOR2X3 U3628 ( .A(n4330), .B(n4346), .Z(n4958) );
  HS65_LH_NAND2X2 U3634 ( .A(\u_DataPath/pc_4_to_ex_i [13]), .B(
        \u_DataPath/pc_4_to_ex_i [12]), .Z(n6754) );
  HS65_LH_NOR2X2 U3640 ( .A(n8508), .B(\u_DataPath/pc_4_to_ex_i [12]), .Z(
        n5789) );
  HS65_LH_CNIVX3 U3646 ( .A(n2811), .Z(n2812) );
  HS65_LH_CNIVX3 U3649 ( .A(n5883), .Z(n5836) );
  HS65_LH_NOR2X2 U3651 ( .A(n5832), .B(n5835), .Z(n5795) );
  HS65_LH_OAI21X3 U3656 ( .A(n5913), .B(n5910), .C(n5912), .Z(n5734) );
  HS65_LL_OAI21X2 U3657 ( .A(n4563), .B(n4659), .C(n4282), .Z(n4301) );
  HS65_LH_NOR2X2 U3659 ( .A(n7965), .B(n7391), .Z(n7611) );
  HS65_LH_CNIVX3 U3660 ( .A(n5867), .Z(n5757) );
  HS65_LH_NOR2X2 U3661 ( .A(n8526), .B(\u_DataPath/pc_4_to_ex_i [26]), .Z(
        n5562) );
  HS65_LH_NOR2X2 U3662 ( .A(n8504), .B(\u_DataPath/pc_4_to_ex_i [14]), .Z(
        n5570) );
  HS65_LH_NAND2X2 U3663 ( .A(n8525), .B(\u_DataPath/pc_4_to_ex_i [9]), .Z(
        n5690) );
  HS65_LH_CNIVX3 U3664 ( .A(\u_DataPath/cw_tomem_i [6]), .Z(n3431) );
  HS65_LH_NAND2X2 U3665 ( .A(n7365), .B(n7379), .Z(n7374) );
  HS65_LH_CNIVX3 U3667 ( .A(\u_DataPath/dataOut_exe_i [9]), .Z(n3034) );
  HS65_LH_CNIVX3 U3674 ( .A(\u_DataPath/pc_4_to_ex_i [25]), .Z(n7636) );
  HS65_LH_NOR2X2 U3676 ( .A(n7435), .B(n7616), .Z(n7621) );
  HS65_LL_NOR2X2 U3677 ( .A(n4443), .B(n4442), .Z(n4453) );
  HS65_LH_CNIVX3 U3678 ( .A(\u_DataPath/from_alu_data_out_i [2]), .Z(n2971) );
  HS65_LH_NAND2X2 U3680 ( .A(n8498), .B(\u_DataPath/u_execute/link_value_i [1]), .Z(n5863) );
  HS65_LH_NAND2X2 U3685 ( .A(n8523), .B(\u_DataPath/pc_4_to_ex_i [6]), .Z(
        n5698) );
  HS65_LHS_XNOR2X3 U3686 ( .A(\u_DataPath/cw_tomem_i [3]), .B(n3431), .Z(n3432) );
  HS65_LH_OAI21X3 U3687 ( .A(n8688), .B(n8766), .C(n8023), .Z(n7999) );
  HS65_LH_CNIVX3 U3688 ( .A(addr_to_iram_28), .Z(n7407) );
  HS65_LH_CNIVX3 U3689 ( .A(n7377), .Z(n7452) );
  HS65_LH_IVX18 U3693 ( .A(n3054), .Z(n2793) );
  HS65_LH_MUXI21X5 U3696 ( .D0(n7675), .D1(n2927), .S0(n3235), .Z(n8066) );
  HS65_LH_NAND2X2 U3700 ( .A(n8500), .B(\u_DataPath/u_execute/link_value_i [0]), .Z(n5865) );
  HS65_LH_NAND2X2 U3702 ( .A(n8441), .B(n7302), .Z(n8320) );
  HS65_LH_NOR2X2 U3703 ( .A(opcode_i[4]), .B(n7333), .Z(n7403) );
  HS65_LH_NAND2X2 U3704 ( .A(n6748), .B(\u_DataPath/cw_tomem_i [0]), .Z(n8131)
         );
  HS65_LH_NOR2X2 U3706 ( .A(\u_DataPath/cw_tomem_i [3]), .B(
        \u_DataPath/cw_tomem_i [6]), .Z(n3429) );
  HS65_LH_CNIVX3 U3707 ( .A(n3443), .Z(n3444) );
  HS65_LHS_XNOR2X3 U3709 ( .A(n7357), .B(n7385), .Z(\u_DataPath/pc_4_i [14])
         );
  HS65_LH_NOR2X2 U3710 ( .A(n9080), .B(rst), .Z(n7943) );
  HS65_LH_OR3ABCX9 U3712 ( .A(n9184), .B(n8007), .C(n9170), .Z(n8004) );
  HS65_LH_AOI22X1 U3713 ( .A(\sub_x_51/A[18] ), .B(n7679), .C(n7681), .D(
        \u_DataPath/u_execute/resAdd1_i [18]), .Z(n8146) );
  HS65_LH_NOR2X6 U3715 ( .A(n9398), .B(n2794), .Z(n8403) );
  HS65_LH_CNIVX3 U3716 ( .A(n7780), .Z(n7784) );
  HS65_LH_CNIVX3 U3717 ( .A(n7660), .Z(n8298) );
  HS65_LH_CNIVX3 U3718 ( .A(n7773), .Z(n7777) );
  HS65_LH_CNIVX3 U3719 ( .A(n7878), .Z(n7882) );
  HS65_LH_CNIVX3 U3720 ( .A(n7815), .Z(n7819) );
  HS65_LH_OAI21X3 U3724 ( .A(n8222), .B(n8456), .C(n8223), .Z(n8308) );
  HS65_LH_NAND2X2 U3725 ( .A(n3443), .B(n2805), .Z(n8267) );
  HS65_LH_BFX9 U3726 ( .A(n8316), .Z(n7696) );
  HS65_LH_NAND2X2 U3727 ( .A(n8789), .B(n7950), .Z(n7947) );
  HS65_LH_CNIVX3 U3728 ( .A(n8131), .Z(n6749) );
  HS65_LH_CNIVX3 U3729 ( .A(n8084), .Z(\u_DataPath/pc4_to_idexreg_i [26]) );
  HS65_LH_CNIVX3 U3733 ( .A(n8132), .Z(\u_DataPath/jump_address_i [29]) );
  HS65_LH_OAI22X1 U3734 ( .A(n6861), .B(n7861), .C(n7716), .D(n8060), .Z(
        \u_DataPath/data_read_ex_2_i [14]) );
  HS65_LH_OAI22X1 U3737 ( .A(n6861), .B(n7840), .C(n7716), .D(n8058), .Z(
        \u_DataPath/data_read_ex_2_i [25]) );
  HS65_LH_OAI22X1 U3738 ( .A(n7719), .B(n7889), .C(n7718), .D(n8272), .Z(
        \u_DataPath/data_read_ex_2_i [22]) );
  HS65_LH_OAI22X1 U3740 ( .A(n7701), .B(n7805), .C(n7699), .D(n8243), .Z(
        \u_DataPath/data_read_ex_1_i [18]) );
  HS65_LH_NOR2X2 U3741 ( .A(n9389), .B(rst), .Z(n8522) );
  HS65_LH_CNIVX3 U3742 ( .A(n7935), .Z(n8508) );
  HS65_LH_NOR3X1 U3743 ( .A(n8807), .B(n9063), .C(n7956), .Z(
        \u_DataPath/u_idexreg/N13 ) );
  HS65_LH_CNIVX3 U3744 ( .A(n8101), .Z(\u_DataPath/pc4_to_idexreg_i [15]) );
  HS65_LH_CNIVX3 U3745 ( .A(n8135), .Z(\u_DataPath/branch_target_i [27]) );
  HS65_LH_CNIVX3 U3746 ( .A(n8172), .Z(\u_DataPath/branch_target_i [10]) );
  HS65_LL_OR2X18 U3748 ( .A(n9366), .B(n2800), .Z(n2772) );
  HS65_LL_OAI12X5 U3751 ( .A(n3271), .B(n3455), .C(n3270), .Z(n4692) );
  HS65_LL_OAI21X6 U3752 ( .A(n9142), .B(n8357), .C(n7658), .Z(n7657) );
  HS65_LL_NOR2X6 U3756 ( .A(\u_DataPath/RFaddr_out_memwb_i [4]), .B(
        \u_DataPath/RFaddr_out_memwb_i [2]), .Z(n2880) );
  HS65_LLS_XNOR2X6 U3757 ( .A(\u_DataPath/idex_rt_i [3]), .B(n8028), .Z(n2914)
         );
  HS65_LL_OA12X4 U3759 ( .A(n5160), .B(n5159), .C(n5158), .Z(n2850) );
  HS65_LL_NOR2X2 U3761 ( .A(n3812), .B(n3811), .Z(n3813) );
  HS65_LL_AOI12X2 U3768 ( .A(n3911), .B(n4829), .C(n3910), .Z(n3912) );
  HS65_LL_IVX2 U3774 ( .A(n4746), .Z(n3331) );
  HS65_LL_NAND2X2 U3777 ( .A(n5498), .B(n3128), .Z(n3643) );
  HS65_LL_NAND2AX7 U3778 ( .A(n3153), .B(n3152), .Z(n4383) );
  HS65_LL_IVX2 U3788 ( .A(n3787), .Z(n3790) );
  HS65_LL_AOI12X2 U3789 ( .A(\sub_x_51/A[21] ), .B(n4208), .C(n3714), .Z(n3787) );
  HS65_LL_NAND2X2 U3793 ( .A(n3883), .B(n4090), .Z(n3615) );
  HS65_LLS_XNOR2X3 U3795 ( .A(n4582), .B(n4581), .Z(n4583) );
  HS65_LL_NOR2X5 U3796 ( .A(n4658), .B(n3397), .Z(n4514) );
  HS65_LL_AOI22X1 U3800 ( .A(n4667), .B(n4789), .C(n4829), .D(n3696), .Z(n3697) );
  HS65_LL_AO12X9 U3807 ( .A(n3036), .B(n7329), .C(n2836), .Z(n5079) );
  HS65_LL_AOI12X2 U3808 ( .A(\lte_x_57/B[2] ), .B(n3742), .C(n3319), .Z(n3917)
         );
  HS65_LL_MUX21I1X6 U3819 ( .D0(n8447), .D1(n8730), .S0(n3174), .Z(n5190) );
  HS65_LL_NAND2AX7 U3824 ( .A(n3147), .B(n3146), .Z(n3993) );
  HS65_LL_IVX2 U3826 ( .A(n3925), .Z(n2784) );
  HS65_LL_NAND3X5 U3836 ( .A(n4116), .B(n4115), .C(n4114), .Z(n4831) );
  HS65_LL_MUXI21X2 U3837 ( .D0(\u_DataPath/from_alu_data_out_i [10]), .D1(
        \u_DataPath/from_mem_data_out_i [10]), .S0(n3235), .Z(n8160) );
  HS65_LL_NAND2X7 U3840 ( .A(n4433), .B(n3326), .Z(n5499) );
  HS65_LL_MUX21I1X6 U3841 ( .D0(n8448), .D1(n8730), .S0(n3174), .Z(n3106) );
  HS65_LL_NAND2X2 U3849 ( .A(n4647), .B(n4639), .Z(n4649) );
  HS65_LL_AOI21X2 U3855 ( .A(n4433), .B(n4045), .C(n3413), .Z(n3414) );
  HS65_LL_AOI21X4 U3856 ( .A(n9269), .B(n7664), .C(n7657), .Z(n7663) );
  HS65_LL_OAI12X3 U3857 ( .A(n7668), .B(n8356), .C(n7667), .Z(n7666) );
  HS65_LL_NAND2X4 U3858 ( .A(n8315), .B(n8327), .Z(n7661) );
  HS65_LH_OAI21X6 U3860 ( .A(n9044), .B(n8654), .C(n8255), .Z(
        \u_DataPath/dataOut_exe_i [25]) );
  HS65_LH_IVX9 U3861 ( .A(n8678), .Z(\u_DataPath/dataOut_exe_i [15]) );
  HS65_LL_AOI22X3 U3863 ( .A(\u_DataPath/u_execute/link_value_i [13]), .B(
        n7694), .C(n8315), .D(n8348), .Z(n8161) );
  HS65_LL_OAI12X3 U3864 ( .A(n9044), .B(n8779), .C(n8592), .Z(
        \u_DataPath/dataOut_exe_i [17]) );
  HS65_LL_AOI22X3 U3866 ( .A(\u_DataPath/u_execute/link_value_i [15]), .B(
        n7694), .C(n8315), .D(n8345), .Z(n8299) );
  HS65_LH_IVX9 U3867 ( .A(n3658), .Z(n3663) );
  HS65_LL_NOR2AX3 U3868 ( .A(n5478), .B(n5477), .Z(n5526) );
  HS65_LH_IVX9 U3875 ( .A(n8218), .Z(\u_DataPath/dataOut_exe_i [7]) );
  HS65_LL_AOI22X3 U3878 ( .A(\u_DataPath/u_execute/link_value_i [7]), .B(n7695), .C(n8315), .D(n8344), .Z(n8218) );
  HS65_LL_NOR2X2 U3882 ( .A(n4678), .B(n4677), .Z(n4699) );
  HS65_LL_NOR2X2 U3885 ( .A(n4744), .B(n4562), .Z(n3461) );
  HS65_LL_NAND2X2 U3895 ( .A(n5470), .B(n5469), .Z(n5471) );
  HS65_LH_NOR2X2 U3897 ( .A(n4653), .B(n4031), .Z(n3409) );
  HS65_LL_OAI22X1 U3916 ( .A(n4564), .B(n4563), .C(n4665), .D(n4562), .Z(n4565) );
  HS65_LH_CB4I1X9 U3918 ( .A(n5388), .B(n5034), .C(n5428), .D(n5033), .Z(n2837) );
  HS65_LL_NAND2X2 U3924 ( .A(n4671), .B(n4843), .Z(n4220) );
  HS65_LL_NOR3X1 U3931 ( .A(n2789), .B(n4147), .C(n4146), .Z(n4167) );
  HS65_LL_NAND2X2 U3941 ( .A(n4595), .B(n3201), .Z(n3203) );
  HS65_LH_OAI112X3 U3943 ( .A(n5390), .B(n5389), .C(n5388), .D(n5387), .Z(
        n5401) );
  HS65_LH_OA12X9 U3944 ( .A(n4690), .B(n4689), .C(n4688), .Z(n2835) );
  HS65_LH_NAND2X2 U3958 ( .A(n3248), .B(n4375), .Z(n3542) );
  HS65_LH_NAND3X3 U3974 ( .A(\lte_x_57/B[30] ), .B(n5446), .C(n2790), .Z(n4009) );
  HS65_LL_NOR2X2 U3976 ( .A(n3676), .B(n3673), .Z(n3261) );
  HS65_LL_NOR2X2 U3992 ( .A(\lte_x_57/B[3] ), .B(n2995), .Z(n4765) );
  HS65_LH_NOR2X5 U4003 ( .A(n5077), .B(n4203), .Z(n5372) );
  HS65_LH_NAND2X4 U4007 ( .A(\lte_x_57/B[3] ), .B(n3251), .Z(n4801) );
  HS65_LH_NAND2X4 U4019 ( .A(\lte_x_57/B[15] ), .B(n5496), .Z(n3402) );
  HS65_LH_NOR2X3 U4024 ( .A(n3951), .B(n5089), .Z(n5333) );
  HS65_LH_NAND2X7 U4028 ( .A(n4680), .B(n4679), .Z(n4697) );
  HS65_LH_NAND2X4 U4029 ( .A(\lte_x_57/B[11] ), .B(n5498), .Z(n3460) );
  HS65_LH_NOR2X3 U4032 ( .A(\lte_x_57/B[30] ), .B(n2790), .Z(n5146) );
  HS65_LL_AOI22X1 U4041 ( .A(\add_x_50/A[23] ), .B(n3826), .C(n2792), .D(
        \sub_x_51/A[20] ), .Z(n3345) );
  HS65_LH_NAND2X7 U4043 ( .A(n8401), .B(n3020), .Z(n3021) );
  HS65_LL_NAND2X4 U4046 ( .A(\lte_x_57/B[7] ), .B(n4208), .Z(n4315) );
  HS65_LL_NOR2X2 U4047 ( .A(n7321), .B(n5148), .Z(n5266) );
  HS65_LL_NAND2X4 U4048 ( .A(\lte_x_57/B[7] ), .B(n4346), .Z(n4338) );
  HS65_LH_OAI22X3 U4051 ( .A(n7302), .B(n7725), .C(n7698), .D(n8059), .Z(
        \u_DataPath/data_read_ex_1_i [0]) );
  HS65_LH_OAI22X3 U4052 ( .A(n7302), .B(n8298), .C(n7698), .D(n8057), .Z(
        \u_DataPath/data_read_ex_1_i [3]) );
  HS65_LH_AOI22X3 U4053 ( .A(\lte_x_57/B[6] ), .B(n7679), .C(n7681), .D(
        \u_DataPath/u_execute/resAdd1_i [6]), .Z(n8176) );
  HS65_LH_OAI22X3 U4056 ( .A(n7302), .B(n8282), .C(n7698), .D(n8056), .Z(
        \u_DataPath/data_read_ex_1_i [2]) );
  HS65_LH_OAI22X3 U4057 ( .A(n7302), .B(n7896), .C(n7698), .D(n8198), .Z(
        \u_DataPath/data_read_ex_1_i [19]) );
  HS65_LH_OAI22X4 U4058 ( .A(n6861), .B(n8055), .C(n7716), .D(n8018), .Z(
        \u_DataPath/data_read_ex_2_i [4]) );
  HS65_LH_OAI22X3 U4059 ( .A(n7302), .B(n7739), .C(n7698), .D(n8207), .Z(
        \u_DataPath/data_read_ex_1_i [27]) );
  HS65_LH_OAI22X3 U4060 ( .A(n7302), .B(n7875), .C(n7698), .D(n8188), .Z(
        \u_DataPath/data_read_ex_1_i [16]) );
  HS65_LH_OAI22X3 U4061 ( .A(n7302), .B(n8055), .C(n7698), .D(n8054), .Z(
        \u_DataPath/data_read_ex_1_i [4]) );
  HS65_LH_OAI22X3 U4062 ( .A(n7302), .B(n7917), .C(n7698), .D(n8050), .Z(
        \u_DataPath/data_read_ex_1_i [1]) );
  HS65_LH_OAI22X3 U4063 ( .A(n7302), .B(n7784), .C(n7699), .D(n8217), .Z(
        \u_DataPath/data_read_ex_1_i [11]) );
  HS65_LH_OAI22X3 U4064 ( .A(n7302), .B(n7882), .C(n7698), .D(n8189), .Z(
        \u_DataPath/data_read_ex_1_i [24]) );
  HS65_LH_OAI22X3 U4065 ( .A(n7302), .B(n7847), .C(n7699), .D(n8211), .Z(
        \u_DataPath/data_read_ex_1_i [23]) );
  HS65_LH_OAI22X3 U4066 ( .A(n7302), .B(n7753), .C(n7698), .D(n8194), .Z(
        \u_DataPath/data_read_ex_1_i [17]) );
  HS65_LH_OAI211X4 U4067 ( .A(n8318), .B(n8302), .C(n8167), .D(n7696), .Z(
        \u_DataPath/from_mem_data_out_i [13]) );
  HS65_LH_IVX7 U4068 ( .A(n8081), .Z(\u_DataPath/pc4_to_idexreg_i [28]) );
  HS65_LH_OAI211X4 U4069 ( .A(n8231), .B(n8302), .C(n8230), .D(n7696), .Z(
        \u_DataPath/from_mem_data_out_i [8]) );
  HS65_LH_OAI211X4 U4070 ( .A(n8302), .B(n8260), .C(n8259), .D(n7696), .Z(
        \u_DataPath/from_mem_data_out_i [9]) );
  HS65_LH_OAI211X4 U4071 ( .A(n8250), .B(n8302), .C(n8234), .D(n7696), .Z(
        \u_DataPath/from_mem_data_out_i [10]) );
  HS65_LL_NOR3X1 U4073 ( .A(n3174), .B(n8682), .C(n2772), .Z(n3095) );
  HS65_LH_OAI211X4 U4074 ( .A(n8216), .B(n8302), .C(n8215), .D(n7696), .Z(
        \u_DataPath/from_mem_data_out_i [11]) );
  HS65_LH_OAI211X4 U4075 ( .A(n8294), .B(n8302), .C(n8239), .D(n7696), .Z(
        \u_DataPath/from_mem_data_out_i [12]) );
  HS65_LH_OAI211X4 U4076 ( .A(n8288), .B(n8302), .C(n8253), .D(n7696), .Z(
        \u_DataPath/from_mem_data_out_i [14]) );
  HS65_LH_OAI211X4 U4078 ( .A(n8311), .B(n8302), .C(n8301), .D(n7696), .Z(
        \u_DataPath/from_mem_data_out_i [15]) );
  HS65_LH_CNIVX3 U4080 ( .A(n8073), .Z(\u_DataPath/cw_to_ex_i [20]) );
  HS65_LH_AOI22X4 U4083 ( .A(n3128), .B(n7679), .C(n7681), .D(
        \u_DataPath/u_execute/resAdd1_i [17]), .Z(n8147) );
  HS65_LH_IVX4 U4085 ( .A(n7946), .Z(\u_DataPath/cw_to_ex_i [15]) );
  HS65_LH_CNIVX3 U4086 ( .A(n8359), .Z(\u_DataPath/cw_exmem_i [0]) );
  HS65_LH_NOR2X3 U4087 ( .A(n9418), .B(n8359), .Z(\u_DataPath/cw_to_ex_i [19])
         );
  HS65_LH_NOR2X2 U4088 ( .A(n8882), .B(n7947), .Z(\u_DataPath/cw_exmem_i [6])
         );
  HS65_LH_AO22X9 U4089 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][26] ), .B(n9156), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][26] ), .D(
        n9475), .Z(n6936) );
  HS65_LL_NOR3X2 U4093 ( .A(n8165), .B(nibble[0]), .C(n8222), .Z(n8306) );
  HS65_LH_OAI112X3 U4095 ( .A(n8407), .B(n2794), .C(n8406), .D(n8441), .Z(
        n8408) );
  HS65_LH_NAND2X4 U4096 ( .A(n9303), .B(n7950), .Z(n8359) );
  HS65_LH_NOR2X6 U4097 ( .A(n3142), .B(n2794), .Z(n8430) );
  HS65_LH_AOI22X3 U4098 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][2] ), .B(n9226), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][2] ), .D(n9193), .Z(n6230) );
  HS65_LH_AO22X9 U4099 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][4] ), .B(n9251), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][4] ), .D(
        n9155), .Z(n6427) );
  HS65_LH_AO22X9 U4102 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][13] ), .B(n9156), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][13] ), .D(
        n9475), .Z(n6402) );
  HS65_LH_AO22X9 U4103 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][14] ), .B(n9156), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][14] ), .D(
        n9475), .Z(n6867) );
  HS65_LH_AO22X9 U4104 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][21] ), .B(n9156), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][21] ), .D(
        n9475), .Z(n6382) );
  HS65_LH_NAND2X5 U4108 ( .A(n1885), .B(n8958), .Z(n8101) );
  HS65_LH_NAND2X5 U4109 ( .A(n1885), .B(n9145), .Z(n8103) );
  HS65_LH_IVX9 U4110 ( .A(n7705), .Z(n7704) );
  HS65_LH_NOR2X5 U4111 ( .A(n8666), .B(n3149), .Z(n3126) );
  HS65_LH_NAND2X5 U4112 ( .A(n1885), .B(n8960), .Z(n8095) );
  HS65_LH_NAND2X5 U4113 ( .A(n1885), .B(n8962), .Z(n8093) );
  HS65_LH_NAND2X5 U4114 ( .A(n1885), .B(n9017), .Z(n8090) );
  HS65_LH_NAND2X2 U4115 ( .A(n1885), .B(n8460), .Z(\u_DataPath/u_fetch/pc1/N3 ) );
  HS65_LH_NAND2X5 U4118 ( .A(n1885), .B(n8959), .Z(n8105) );
  HS65_LH_AOI21X2 U4119 ( .A(n8751), .B(n2798), .C(n3119), .Z(n3120) );
  HS65_LH_IVX4 U4120 ( .A(n8112), .Z(\u_DataPath/pc4_to_idexreg_i [8]) );
  HS65_LH_IVX4 U4123 ( .A(n8114), .Z(\u_DataPath/pc4_to_idexreg_i [7]) );
  HS65_LH_NOR2X5 U4124 ( .A(\u_DataPath/dataOut_exe_i [20]), .B(n3178), .Z(
        n3172) );
  HS65_LH_IVX4 U4126 ( .A(n8109), .Z(\u_DataPath/pc4_to_idexreg_i [10]) );
  HS65_LH_NOR2X5 U4127 ( .A(\u_DataPath/dataOut_exe_i [17]), .B(n3178), .Z(
        n3127) );
  HS65_LH_NOR2X5 U4132 ( .A(n9125), .B(n3178), .Z(n3098) );
  HS65_LH_NOR2X5 U4133 ( .A(\u_DataPath/dataOut_exe_i [23]), .B(n3178), .Z(
        n3159) );
  HS65_LH_NAND2X4 U4136 ( .A(n1885), .B(n9074), .Z(n8109) );
  HS65_LH_NAND2X4 U4137 ( .A(n1885), .B(n8953), .Z(n8114) );
  HS65_LH_NAND2X4 U4147 ( .A(n9382), .B(n2800), .Z(n8395) );
  HS65_LH_NAND2X4 U4151 ( .A(n9459), .B(n2800), .Z(n8396) );
  HS65_LH_NOR2X2 U4152 ( .A(\u_DataPath/dataOut_exe_i [12]), .B(n9012), .Z(
        n3053) );
  HS65_LH_NAND2X4 U4153 ( .A(addr_to_iram_8), .B(n7461), .Z(n7462) );
  HS65_LH_OAI21X3 U4154 ( .A(n2819), .B(n7613), .C(n7612), .Z(n7992) );
  HS65_LH_NOR2X2 U4155 ( .A(n9541), .B(n9012), .Z(n2937) );
  HS65_LH_NAND2X4 U4156 ( .A(n3130), .B(n2800), .Z(n8425) );
  HS65_LH_CNIVX3 U4157 ( .A(n8118), .Z(\u_DataPath/pc4_to_idexreg_i [4]) );
  HS65_LH_IVX4 U4159 ( .A(n3563), .Z(n8458) );
  HS65_LH_NOR2X3 U4160 ( .A(n7710), .B(n7654), .Z(n8483) );
  HS65_LH_NOR2X3 U4161 ( .A(n7710), .B(n8751), .Z(n8485) );
  HS65_LHS_XOR2X3 U4163 ( .A(n7460), .B(n7459), .Z(\u_DataPath/pc_4_i [5]) );
  HS65_LH_NOR2X2 U4164 ( .A(n7711), .B(n8278), .Z(n8462) );
  HS65_LH_NAND2X2 U4165 ( .A(n1885), .B(n8936), .Z(n8118) );
  HS65_LL_NAND2X4 U4166 ( .A(n2892), .B(n2914), .Z(n2899) );
  HS65_LH_NOR2X5 U4169 ( .A(n7344), .B(n7446), .Z(n7464) );
  HS65_LH_NOR2X3 U4172 ( .A(n7710), .B(n8719), .Z(n8494) );
  HS65_LH_NOR2X2 U4174 ( .A(n7711), .B(n8721), .Z(n8487) );
  HS65_LH_NOR2X2 U4175 ( .A(n7710), .B(n8695), .Z(n8486) );
  HS65_LH_NOR2X2 U4176 ( .A(n7712), .B(n8692), .Z(n8488) );
  HS65_LLS_XNOR2X3 U4177 ( .A(n2864), .B(n7014), .Z(n2866) );
  HS65_LH_NAND2X4 U4178 ( .A(addr_to_iram_2), .B(n7458), .Z(n7459) );
  HS65_LH_NOR2X2 U4179 ( .A(n7711), .B(n8697), .Z(n8493) );
  HS65_LH_NOR2X2 U4180 ( .A(n7711), .B(n8717), .Z(n8495) );
  HS65_LL_NAND2X2 U4181 ( .A(n3437), .B(n3436), .Z(n3443) );
  HS65_LL_NOR2X6 U4182 ( .A(n2882), .B(n2903), .Z(n2883) );
  HS65_LH_NAND2X2 U4183 ( .A(n1885), .B(n8997), .Z(n8120) );
  HS65_LH_NOR2X2 U4184 ( .A(n7711), .B(n8696), .Z(n8471) );
  HS65_LH_NOR2X3 U4185 ( .A(n7712), .B(n8698), .Z(n8478) );
  HS65_LH_NOR2X2 U4186 ( .A(n7710), .B(n8691), .Z(n8484) );
  HS65_LH_NOR2X2 U4187 ( .A(n7711), .B(n8699), .Z(n8476) );
  HS65_LH_NOR2X6 U4188 ( .A(n5745), .B(n5777), .Z(n5747) );
  HS65_LH_NOR2X2 U4191 ( .A(n8245), .B(n7711), .Z(n8481) );
  HS65_LH_CNIVX3 U4192 ( .A(n7379), .Z(n7380) );
  HS65_LH_NOR2X2 U4193 ( .A(n7710), .B(n8701), .Z(n8491) );
  HS65_LH_CNIVX3 U4194 ( .A(n5827), .Z(n5828) );
  HS65_LH_NOR2X2 U4195 ( .A(n7712), .B(n8693), .Z(n8492) );
  HS65_LHS_XNOR2X3 U4197 ( .A(n7416), .B(n7618), .Z(
        \u_DataPath/u_execute/link_value_i [4]) );
  HS65_LH_NOR2X2 U4198 ( .A(n7710), .B(n8718), .Z(n8482) );
  HS65_LH_NOR2X2 U4199 ( .A(n7711), .B(n8709), .Z(n8480) );
  HS65_LH_NOR2X2 U4200 ( .A(n7712), .B(n8724), .Z(n8479) );
  HS65_LH_NOR2X2 U4201 ( .A(n7712), .B(n8694), .Z(n8473) );
  HS65_LH_NOR2X2 U4202 ( .A(n7712), .B(n8690), .Z(n8496) );
  HS65_LL_NOR3X1 U4204 ( .A(n9445), .B(n8752), .C(n8154), .Z(n8314) );
  HS65_LH_IVX7 U4205 ( .A(n7942), .Z(n8506) );
  HS65_LH_IVX7 U4206 ( .A(n7939), .Z(n8510) );
  HS65_LH_IVX7 U4207 ( .A(n7938), .Z(n8504) );
  HS65_LH_IVX7 U4208 ( .A(n8063), .Z(n8469) );
  HS65_LH_IVX7 U4209 ( .A(n8074), .Z(n8525) );
  HS65_LH_IVX7 U4210 ( .A(n8075), .Z(n8524) );
  HS65_LH_IVX7 U4211 ( .A(n8065), .Z(n8474) );
  HS65_LH_IVX7 U4212 ( .A(n8076), .Z(n8523) );
  HS65_LL_NAND3X5 U4216 ( .A(n2879), .B(n2878), .C(n2877), .Z(n2882) );
  HS65_LH_IVX7 U4218 ( .A(n7964), .Z(n7398) );
  HS65_LH_NOR2X5 U4223 ( .A(n9419), .B(rst), .Z(n8500) );
  HS65_LH_NAND2X5 U4224 ( .A(n5667), .B(n5532), .Z(n5556) );
  HS65_LH_NOR2X5 U4225 ( .A(n9420), .B(rst), .Z(n8498) );
  HS65_LH_NAND2X2 U4226 ( .A(n1885), .B(n8872), .Z(n8182) );
  HS65_LH_CNIVX3 U4227 ( .A(n7384), .Z(n7386) );
  HS65_LH_NOR2X5 U4228 ( .A(n9311), .B(rst), .Z(n8466) );
  HS65_LH_NAND2AX4 U4229 ( .A(n7714), .B(n8815), .Z(n7942) );
  HS65_LH_NAND2AX4 U4230 ( .A(n7714), .B(n8803), .Z(n7935) );
  HS65_LH_NAND2AX4 U4231 ( .A(n7714), .B(n8809), .Z(n7939) );
  HS65_LH_NAND2AX4 U4232 ( .A(n7714), .B(n8808), .Z(n7938) );
  HS65_LH_IVX35 U4233 ( .A(n7650), .Z(n3148) );
  HS65_LH_IVX4 U4234 ( .A(addr_to_iram_9), .Z(n7463) );
  HS65_LH_IVX4 U4235 ( .A(addr_to_iram_11), .Z(n7363) );
  HS65_LH_IVX4 U4236 ( .A(n5619), .Z(n5680) );
  HS65_LH_IVX4 U4237 ( .A(n5685), .Z(n5597) );
  HS65_LH_IVX4 U4238 ( .A(addr_to_iram_7), .Z(n7466) );
  HS65_LH_CNIVX3 U4239 ( .A(addr_to_iram_8), .Z(n7343) );
  HS65_LH_NAND2X4 U4240 ( .A(n5867), .B(n5866), .Z(n5869) );
  HS65_LH_CNIVX3 U4241 ( .A(addr_to_iram_6), .Z(n7345) );
  HS65_LH_IVX4 U4242 ( .A(addr_to_iram_13), .Z(n7359) );
  HS65_LH_IVX4 U4243 ( .A(addr_to_iram_19), .Z(n7472) );
  HS65_LH_IVX4 U4244 ( .A(addr_to_iram_15), .Z(n7388) );
  HS65_LH_IVX7 U4245 ( .A(\u_DataPath/immediate_ext_dec_i [2]), .Z(n8030) );
  HS65_LH_IVX4 U4246 ( .A(addr_to_iram_18), .Z(n7383) );
  HS65_LH_IVX4 U4247 ( .A(\u_DataPath/immediate_ext_dec_i [1]), .Z(n8053) );
  HS65_LH_IVX4 U4248 ( .A(addr_to_iram_24), .Z(n7378) );
  HS65_LH_IVX7 U4249 ( .A(\u_DataPath/immediate_ext_dec_i [0]), .Z(n8051) );
  HS65_LH_CNIVX3 U4250 ( .A(addr_to_iram_2), .Z(n7331) );
  HS65_LH_CNIVX3 U4251 ( .A(addr_to_iram_3), .Z(n7460) );
  HS65_LH_IVX7 U4252 ( .A(addr_to_iram_4), .Z(n7447) );
  HS65_LH_CNIVX3 U4253 ( .A(addr_to_iram_5), .Z(n7339) );
  HS65_LH_CNIVX3 U4254 ( .A(opcode_i[0]), .Z(n8321) );
  HS65_LL_NAND2X4 U4255 ( .A(n3434), .B(n3438), .Z(n7351) );
  HS65_LH_IVX4 U4256 ( .A(n5603), .Z(n5604) );
  HS65_LH_NAND2X4 U4257 ( .A(opcode_i[3]), .B(opcode_i[4]), .Z(n7391) );
  HS65_LH_CNIVX3 U4258 ( .A(n7421), .Z(n7424) );
  HS65_LL_CNIVX21 U4259 ( .A(n7650), .Z(n3235) );
  HS65_LH_IVX4 U4260 ( .A(addr_to_iram_17), .Z(n7373) );
  HS65_LH_IVX7 U4261 ( .A(addr_to_iram_26), .Z(n7390) );
  HS65_LH_CNIVX3 U4262 ( .A(n5704), .Z(n5654) );
  HS65_LH_CNIVX3 U4263 ( .A(n5854), .Z(n5906) );
  HS65_LH_NOR2X5 U4264 ( .A(n8512), .B(\u_DataPath/pc_4_to_ex_i [15]), .Z(
        n5770) );
  HS65_LH_NOR2X3 U4265 ( .A(n8498), .B(\u_DataPath/u_execute/link_value_i [1]), 
        .Z(n5861) );
  HS65_LH_NOR2X5 U4266 ( .A(n8510), .B(\u_DataPath/pc_4_to_ex_i [13]), .Z(
        n5808) );
  HS65_LH_NOR2X5 U4267 ( .A(n8467), .B(\u_DataPath/pc_4_to_ex_i [4]), .Z(n5854) );
  HS65_LH_IVX9 U4268 ( .A(\u_DataPath/data_read_ex_2_i [1]), .Z(n2958) );
  HS65_LH_OR2X4 U4269 ( .A(n8515), .B(\u_DataPath/pc_4_to_ex_i [30]), .Z(n5866) );
  HS65_LH_NOR2X5 U4270 ( .A(n8506), .B(\u_DataPath/pc_4_to_ex_i [11]), .Z(
        n5797) );
  HS65_LH_IVX4 U4271 ( .A(\u_DataPath/pc_4_to_ex_i [28]), .Z(n7308) );
  HS65_LH_NOR2X5 U4272 ( .A(n8525), .B(\u_DataPath/pc_4_to_ex_i [9]), .Z(n5890) );
  HS65_LH_NOR2X3 U4273 ( .A(\u_DataPath/rs_ex_i [2]), .B(
        \u_DataPath/pc_4_to_ex_i [23]), .Z(n5839) );
  HS65_LH_NAND2X5 U4274 ( .A(n8522), .B(\u_DataPath/pc_4_to_ex_i [5]), .Z(
        n5853) );
  HS65_LH_NAND2X7 U4275 ( .A(n8524), .B(\u_DataPath/pc_4_to_ex_i [8]), .Z(
        n5691) );
  HS65_LH_NOR2X5 U4276 ( .A(n8523), .B(\u_DataPath/pc_4_to_ex_i [6]), .Z(n5903) );
  HS65_LH_NOR2X3 U4277 ( .A(n8515), .B(\u_DataPath/pc_4_to_ex_i [25]), .Z(
        n5784) );
  HS65_LH_NOR2X5 U4278 ( .A(n8474), .B(\u_DataPath/pc_4_to_ex_i [7]), .Z(n5898) );
  HS65_LH_NOR2X3 U4279 ( .A(n8526), .B(\u_DataPath/pc_4_to_ex_i [24]), .Z(
        n5581) );
  HS65_LH_IVX4 U4280 ( .A(\u_DataPath/idex_rt_i [0]), .Z(n7204) );
  HS65_LH_NOR2X3 U4281 ( .A(n8526), .B(\u_DataPath/pc_4_to_ex_i [22]), .Z(
        n5638) );
  HS65_LH_NOR2X5 U4282 ( .A(\u_DataPath/idex_rt_i [1]), .B(
        \u_DataPath/pc_4_to_ex_i [17]), .Z(n5832) );
  HS65_LH_NAND2X7 U4283 ( .A(\u_DataPath/idex_rt_i [3]), .B(
        \u_DataPath/pc_4_to_ex_i [19]), .Z(n5876) );
  HS65_LH_NOR2X6 U4284 ( .A(n8506), .B(\u_DataPath/pc_4_to_ex_i [11]), .Z(
        n5589) );
  HS65_LH_NOR2X6 U4287 ( .A(n8510), .B(\u_DataPath/pc_4_to_ex_i [13]), .Z(
        n5600) );
  HS65_LH_IVX9 U4288 ( .A(\u_DataPath/data_read_ex_2_i [10]), .Z(n3016) );
  HS65_LH_IVX7 U4289 ( .A(\u_DataPath/dataOut_exe_i [4]), .Z(n2947) );
  HS65_LH_IVX4 U4290 ( .A(\u_DataPath/pc_4_to_ex_i [16]), .Z(n7642) );
  HS65_LH_IVX9 U4291 ( .A(\u_DataPath/data_read_ex_2_i [17]), .Z(n3129) );
  HS65_LH_NAND2X2 U4292 ( .A(\u_DataPath/u_execute/ovf_i ), .B(n1885), .Z(
        n8042) );
  HS65_LL_NAND2X4 U4293 ( .A(n7662), .B(n7661), .Z(
        \u_DataPath/dataOut_exe_i [24]) );
  HS65_LL_NAND2X4 U4294 ( .A(n8315), .B(n8326), .Z(n7655) );
  HS65_LL_OAI12X3 U4295 ( .A(n9044), .B(n8755), .C(n8595), .Z(
        \u_DataPath/dataOut_exe_i [21]) );
  HS65_LL_OAI12X3 U4299 ( .A(n9044), .B(n8745), .C(n8249), .Z(
        \u_DataPath/dataOut_exe_i [26]) );
  HS65_LL_AOI22X3 U4300 ( .A(n8952), .B(n7694), .C(n8315), .D(n8322), .Z(n8246) );
  HS65_LL_AOI22X3 U4303 ( .A(\u_DataPath/u_execute/link_value_i [14]), .B(
        n7694), .C(n8315), .D(n8346), .Z(n8252) );
  HS65_LL_AOI22X3 U4306 ( .A(\u_DataPath/u_execute/link_value_i [12]), .B(
        n7694), .C(n8315), .D(n8349), .Z(n8238) );
  HS65_LL_AOI12X2 U4311 ( .A(n2837), .B(n5056), .C(n5055), .Z(n5057) );
  HS65_LL_AOI12X2 U4314 ( .A(n3659), .B(n4732), .C(n4449), .Z(n4450) );
  HS65_LL_OAI22X1 U4316 ( .A(n9505), .B(n4305), .C(n4812), .D(n4430), .Z(n3817) );
  HS65_LL_OAI112X1 U4318 ( .A(n4738), .B(n4483), .C(n4482), .D(n4481), .Z(
        n4484) );
  HS65_LLS_XOR2X3 U4320 ( .A(n4274), .B(n4273), .Z(n4307) );
  HS65_LL_NAND2X2 U4327 ( .A(n4411), .B(n4410), .Z(n4421) );
  HS65_LH_NAND2X4 U4332 ( .A(n4551), .B(n4639), .Z(n3376) );
  HS65_LH_OAI12X3 U4335 ( .A(n3392), .B(n4564), .C(n3391), .Z(n3393) );
  HS65_LL_NAND3X2 U4342 ( .A(n3857), .B(n3856), .C(n4844), .Z(n3858) );
  HS65_LH_OAI21X3 U4358 ( .A(n4014), .B(n4013), .C(n4012), .Z(n4015) );
  HS65_LH_AOI21X2 U4360 ( .A(n5011), .B(n4011), .C(n4010), .Z(n4012) );
  HS65_LH_IVX7 U4372 ( .A(n8128), .Z(\u_DataPath/jump_address_i [31]) );
  HS65_LL_NOR2X2 U4392 ( .A(n4275), .B(n4046), .Z(n4259) );
  HS65_LL_NOR2X3 U4394 ( .A(\sub_x_51/A[20] ), .B(n3192), .Z(n5184) );
  HS65_LH_IVX9 U4395 ( .A(n3320), .Z(n4789) );
  HS65_LL_AOI12X2 U4401 ( .A(\lte_x_57/B[28] ), .B(n3742), .C(n3327), .Z(n4325) );
  HS65_LH_IVX4 U4403 ( .A(n5456), .Z(n5457) );
  HS65_LL_NAND2X7 U4413 ( .A(n5092), .B(n2995), .Z(n4613) );
  HS65_LH_NOR2X5 U4419 ( .A(n5386), .B(n5385), .Z(n5375) );
  HS65_LL_NAND2X2 U4429 ( .A(n4211), .B(n4210), .Z(n4838) );
  HS65_LH_IVX4 U4431 ( .A(n3416), .Z(n3417) );
  HS65_LH_IVX4 U4439 ( .A(n5350), .Z(n5404) );
  HS65_LH_OAI21X3 U4441 ( .A(n2825), .B(n3322), .C(n3625), .Z(n3690) );
  HS65_LH_NOR2X2 U4446 ( .A(rst), .B(n7676), .Z(
        \u_DataPath/mem_writedata_out_i [24]) );
  HS65_LH_NAND2X4 U4450 ( .A(\lte_x_57/B[4] ), .B(n3742), .Z(n4778) );
  HS65_LH_NOR2X6 U4459 ( .A(\lte_x_57/B[28] ), .B(n2791), .Z(n4541) );
  HS65_LH_IVX18 U4460 ( .A(n7321), .Z(n7317) );
  HS65_LH_OAI22X3 U4471 ( .A(n6861), .B(n7917), .C(n7716), .D(n8052), .Z(
        \u_DataPath/data_read_ex_2_i [1]) );
  HS65_LH_OAI22X3 U4472 ( .A(n6861), .B(n7875), .C(n7716), .D(n8069), .Z(
        \u_DataPath/data_read_ex_2_i [16]) );
  HS65_LH_OAI22X3 U4473 ( .A(n6861), .B(n7882), .C(n7716), .D(n8068), .Z(
        \u_DataPath/data_read_ex_2_i [24]) );
  HS65_LH_OAI22X3 U4474 ( .A(n6861), .B(n7777), .C(n7716), .D(n8153), .Z(
        \u_DataPath/data_read_ex_2_i [13]) );
  HS65_LH_OAI22X3 U4475 ( .A(n6861), .B(n7805), .C(n7716), .D(n8061), .Z(
        \u_DataPath/data_read_ex_2_i [18]) );
  HS65_LL_OAI12X5 U4477 ( .A(n3044), .B(n8418), .C(n3043), .Z(n5084) );
  HS65_LH_NOR2X2 U4478 ( .A(rst), .B(n8447), .Z(
        \u_DataPath/mem_writedata_out_i [26]) );
  HS65_LL_AOI12X4 U4480 ( .A(n3090), .B(n8451), .C(n3984), .Z(n7321) );
  HS65_LH_NOR2X2 U4481 ( .A(rst), .B(n2773), .Z(
        \u_DataPath/mem_writedata_out_i [29]) );
  HS65_LH_NAND2X7 U4482 ( .A(n9409), .B(n2797), .Z(n8401) );
  HS65_LH_NOR2X2 U4483 ( .A(rst), .B(n8450), .Z(
        \u_DataPath/mem_writedata_out_i [30]) );
  HS65_LH_NOR2X2 U4484 ( .A(rst), .B(n8449), .Z(
        \u_DataPath/mem_writedata_out_i [28]) );
  HS65_LH_NOR2X6 U4485 ( .A(n2968), .B(n5497), .Z(n3775) );
  HS65_LH_NOR2X5 U4487 ( .A(n8683), .B(n2772), .Z(n8415) );
  HS65_LL_OR2X9 U4488 ( .A(n4870), .B(n9538), .Z(n2830) );
  HS65_LH_NOR2X5 U4489 ( .A(n8638), .B(n2772), .Z(n8418) );
  HS65_LH_IVX7 U4490 ( .A(n8098), .Z(\u_DataPath/pc4_to_idexreg_i [17]) );
  HS65_LH_IVX18 U4491 ( .A(n4383), .Z(\sub_x_51/A[18] ) );
  HS65_LH_AO22X4 U4494 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][30] ), .B(n9254), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][30] ), .D(
        n9064), .Z(n7531) );
  HS65_LH_AO22X9 U4496 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][0] ), .B(n9251), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][0] ), .D(
        n9155), .Z(n6207) );
  HS65_LL_MX41X4 U4500 ( .D0(n8770), .S0(n9478), .D1(n8623), .S1(n9492), .D2(
        n9499), .S2(n8767), .D3(n9081), .S3(n9485), .Z(
        \u_DataPath/from_mem_data_out_i [2]) );
  HS65_LH_NOR2X2 U4503 ( .A(n9418), .B(n7947), .Z(\u_DataPath/u_idexreg/N12 )
         );
  HS65_LH_NOR3X1 U4505 ( .A(n8452), .B(rst), .C(n8451), .Z(n8453) );
  HS65_LH_AO22X9 U4507 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][27] ), .B(n9251), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][27] ), .D(
        n9155), .Z(n6319) );
  HS65_LH_AOI22X3 U4512 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][10] ), .B(n9255), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][10] ), .D(
        n9116), .Z(n6706) );
  HS65_LH_AOI22X3 U4513 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][11] ), .B(n9259), 
        .C(n9256), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][11] ), .Z(n6810)
         );
  HS65_LH_AOI22X3 U4514 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][6] ), .B(n9255), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][6] ), .D(
        n9116), .Z(n6730) );
  HS65_LH_AO22X9 U4518 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][22] ), .B(n9258), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][22] ), .D(
        n9065), .Z(n7180) );
  HS65_LH_AO22X9 U4519 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][15] ), .B(n9153), 
        .C(n9253), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][15] ), .Z(n7263)
         );
  HS65_LH_AOI22X3 U4521 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][8] ), .B(n9255), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][8] ), .D(
        n9116), .Z(n6646) );
  HS65_LH_AOI22X3 U4522 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][15] ), .B(n9248), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][15] ), .D(
        n9163), .Z(n6896) );
  HS65_LH_AOI22X3 U4526 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][12] ), .B(n9255), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][12] ), .D(
        n9116), .Z(n6686) );
  HS65_LH_AOI22X3 U4527 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][15] ), .B(n9159), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][15] ), .D(
        n9265), .Z(n7271) );
  HS65_LL_NAND2X5 U4529 ( .A(n8166), .B(n8219), .Z(n8316) );
  HS65_LH_NOR2X5 U4531 ( .A(n8636), .B(n3181), .Z(n2922) );
  HS65_LL_OAI12X3 U4533 ( .A(n3139), .B(n3137), .C(n3136), .Z(n3138) );
  HS65_LH_AO22X9 U4535 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][2] ), .B(n9251), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][2] ), .D(
        n9155), .Z(n6227) );
  HS65_LH_AO22X9 U4536 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][4] ), .B(n9156), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][4] ), .D(
        n9475), .Z(n6422) );
  HS65_LH_AOI22X3 U4537 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][4] ), .B(n9226), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][4] ), .D(n9193), .Z(n6430) );
  HS65_LL_NAND3X3 U4539 ( .A(n9071), .B(n8046), .C(n8186), .Z(n8223) );
  HS65_LH_NAND2AX4 U4542 ( .A(iram_data[30]), .B(n7706), .Z(opcode_i[4]) );
  HS65_LL_NAND2X2 U4543 ( .A(n2943), .B(n2712), .Z(n2944) );
  HS65_LH_NAND2X7 U4544 ( .A(n9352), .B(n7305), .Z(n7627) );
  HS65_LL_AOI12X4 U4545 ( .A(\u_DataPath/dataOut_exe_i [0]), .B(n8454), .C(
        n8044), .Z(n8186) );
  HS65_LH_NAND2X7 U4546 ( .A(n7693), .B(\u_DataPath/u_execute/link_value_i [9]), .Z(n8258) );
  HS65_LH_IVX7 U4549 ( .A(n8178), .Z(\u_DataPath/branch_target_i [4]) );
  HS65_LH_NAND2X2 U4551 ( .A(n8441), .B(n8396), .Z(n8398) );
  HS65_LH_NAND2X5 U4552 ( .A(n1885), .B(n9014), .Z(n8112) );
  HS65_LH_NOR2X3 U4553 ( .A(n7374), .B(n7452), .Z(n7371) );
  HS65_LH_IVX7 U4555 ( .A(n8361), .Z(n7709) );
  HS65_LH_NAND2X2 U4558 ( .A(\u_DataPath/dataOut_exe_i [26]), .B(n3107), .Z(
        n3111) );
  HS65_LHS_XOR2X3 U4559 ( .A(n9232), .B(n9403), .Z(
        \u_DataPath/u_execute/link_value_i [18]) );
  HS65_LH_NAND2X7 U4560 ( .A(n7693), .B(\u_DataPath/u_execute/link_value_i [8]), .Z(n8229) );
  HS65_LH_NOR2X3 U4561 ( .A(n8734), .B(n9012), .Z(n3038) );
  HS65_LH_NAND2X4 U4563 ( .A(n8664), .B(n2800), .Z(n8389) );
  HS65_LH_IVX7 U4565 ( .A(n7439), .Z(n7639) );
  HS65_LH_NOR2X3 U4568 ( .A(n7711), .B(n8741), .Z(n8489) );
  HS65_LL_NOR2X5 U4571 ( .A(n6184), .B(n6162), .Z(n6259) );
  HS65_LH_NAND2X5 U4572 ( .A(n1885), .B(n8771), .Z(n8226) );
  HS65_LL_NAND2X5 U4573 ( .A(n3553), .B(n3563), .Z(n3566) );
  HS65_LL_NOR2X5 U4574 ( .A(n2874), .B(n2873), .Z(n2887) );
  HS65_LH_IVX7 U4575 ( .A(n8066), .Z(n2931) );
  HS65_LH_IVX4 U4577 ( .A(n8228), .Z(n3029) );
  HS65_LH_NOR2X2 U4579 ( .A(n7710), .B(n8263), .Z(n8497) );
  HS65_LH_NAND2X7 U4580 ( .A(\u_DataPath/reg_write_i ), .B(n2915), .Z(n2894)
         );
  HS65_LH_IVX9 U4581 ( .A(n8693), .Z(n3139) );
  HS65_LHS_XNOR2X3 U4584 ( .A(n9011), .B(n5916), .Z(
        \u_DataPath/u_execute/resAdd1_i [3]) );
  HS65_LH_NOR2X2 U4585 ( .A(n7710), .B(n8774), .Z(n8472) );
  HS65_LH_CNIVX3 U4586 ( .A(n8120), .Z(\u_DataPath/pc4_to_idexreg_i [3]) );
  HS65_LH_NOR2X2 U4587 ( .A(n7711), .B(n8769), .Z(n8470) );
  HS65_LH_NOR2X2 U4589 ( .A(n7711), .B(n8157), .Z(n8499) );
  HS65_LH_NOR2X2 U4590 ( .A(n7711), .B(n8700), .Z(n8490) );
  HS65_LH_IVX4 U4591 ( .A(n8213), .Z(n3007) );
  HS65_LH_NOR2X3 U4592 ( .A(n7710), .B(n8702), .Z(n8477) );
  HS65_LL_NOR2X5 U4593 ( .A(n5961), .B(n5960), .Z(n7587) );
  HS65_LL_NAND2X5 U4595 ( .A(\u_DataPath/jaddr_i [18]), .B(n5944), .Z(n5952)
         );
  HS65_LH_CNIVX3 U4597 ( .A(n7352), .Z(n7353) );
  HS65_LH_CNIVX3 U4598 ( .A(n5632), .Z(n5635) );
  HS65_LH_NOR2X5 U4599 ( .A(n9236), .B(rst), .Z(\u_DataPath/idex_rt_i [3]) );
  HS65_LH_CNIVX3 U4600 ( .A(n5826), .Z(n5829) );
  HS65_LH_CNIVX3 U4602 ( .A(n8182), .Z(\u_DataPath/branch_target_i [0]) );
  HS65_LH_IVX4 U4603 ( .A(n7417), .Z(n7616) );
  HS65_LH_NAND2X4 U4605 ( .A(opcode_i[2]), .B(n7933), .Z(n7930) );
  HS65_LL_NAND2X5 U4606 ( .A(\u_DataPath/cw_memwb_i [2]), .B(n2881), .Z(n2903)
         );
  HS65_LH_CNIVX3 U4607 ( .A(n7415), .Z(n7618) );
  HS65_LH_IVX4 U4610 ( .A(n5571), .Z(n5577) );
  HS65_LH_IVX4 U4611 ( .A(n5575), .Z(n5576) );
  HS65_LL_NAND3X3 U4612 ( .A(n2812), .B(\u_DataPath/jaddr_i [24]), .C(n2817), 
        .Z(n6175) );
  HS65_LH_CNIVX3 U4613 ( .A(n5593), .Z(n5596) );
  HS65_LH_NOR3X3 U4614 ( .A(n9351), .B(n9146), .C(rst), .Z(n8183) );
  HS65_LL_NAND3X3 U4615 ( .A(n2804), .B(n8017), .C(n8016), .Z(n5960) );
  HS65_LL_NAND2X5 U4616 ( .A(\u_DataPath/jaddr_i [17]), .B(n5935), .Z(n5959)
         );
  HS65_LL_NAND2X5 U4617 ( .A(\u_DataPath/jaddr_i [16]), .B(n5936), .Z(n5961)
         );
  HS65_LH_NOR2X6 U4618 ( .A(n7337), .B(n7336), .Z(n7342) );
  HS65_LH_CNIVX3 U4619 ( .A(n7337), .Z(n7458) );
  HS65_LH_NAND2AX4 U4620 ( .A(n7714), .B(n8791), .Z(n8065) );
  HS65_LH_NAND2AX4 U4621 ( .A(n7714), .B(n8793), .Z(n8074) );
  HS65_LH_NAND2AX4 U4622 ( .A(n7714), .B(n8790), .Z(n8075) );
  HS65_LH_NAND2AX4 U4623 ( .A(n7714), .B(n8792), .Z(n8063) );
  HS65_LH_NAND2AX4 U4624 ( .A(n7714), .B(n8814), .Z(n8076) );
  HS65_LH_NOR2X2 U4625 ( .A(n7710), .B(n9171), .Z(\u_DataPath/cw_tomem_i [4])
         );
  HS65_LH_NAND2AX4 U4626 ( .A(n7714), .B(n9080), .Z(n7936) );
  HS65_LH_NAND2X4 U4627 ( .A(n8466), .B(\u_DataPath/pc_4_to_ex_i [3]), .Z(
        n5709) );
  HS65_LH_IVX4 U4628 ( .A(n5773), .Z(n5870) );
  HS65_LH_NOR2X6 U4629 ( .A(n5650), .B(n5653), .Z(n5648) );
  HS65_LH_NOR2X3 U4631 ( .A(n8156), .B(rst), .Z(n8463) );
  HS65_LH_NAND2X2 U4632 ( .A(n1885), .B(n8547), .Z(n8125) );
  HS65_LH_NAND2X2 U4633 ( .A(n1885), .B(n8546), .Z(n8123) );
  HS65_LH_IVX4 U4634 ( .A(n5570), .Z(n5676) );
  HS65_LH_CNIVX3 U4635 ( .A(\u_DataPath/immediate_ext_dec_i [5]), .Z(n8077) );
  HS65_LH_IVX4 U4636 ( .A(n5835), .Z(n5882) );
  HS65_LH_CNIVX3 U4637 ( .A(addr_to_iram_0), .Z(\u_DataPath/pc_4_i [2]) );
  HS65_LH_IVX4 U4638 ( .A(n5586), .Z(n5606) );
  HS65_LH_CNIVX3 U4639 ( .A(addr_to_iram_1), .Z(n7330) );
  HS65_LH_NAND2X5 U4640 ( .A(n5673), .B(n5672), .Z(n5675) );
  HS65_LH_CNIVX3 U4641 ( .A(n5669), .Z(n5532) );
  HS65_LL_NAND2X5 U4642 ( .A(\u_DataPath/jaddr_i [22]), .B(n2815), .Z(n6188)
         );
  HS65_LH_NOR2X2 U4643 ( .A(n9228), .B(rst), .Z(\u_DataPath/u_memwbreg/N74 )
         );
  HS65_LH_NOR2X2 U4644 ( .A(n9219), .B(rst), .Z(\u_DataPath/u_memwbreg/N71 )
         );
  HS65_LH_IVX9 U4645 ( .A(n2815), .Z(n2816) );
  HS65_LH_IVX9 U4646 ( .A(\u_DataPath/jaddr_i [20]), .Z(n8017) );
  HS65_LH_NOR2X2 U4648 ( .A(n9218), .B(rst), .Z(\u_DataPath/u_memwbreg/N72 )
         );
  HS65_LH_NOR2X2 U4649 ( .A(n9220), .B(rst), .Z(\u_DataPath/u_memwbreg/N70 )
         );
  HS65_LH_NAND2X4 U4650 ( .A(n8522), .B(\u_DataPath/pc_4_to_ex_i [5]), .Z(
        n5652) );
  HS65_LH_NAND2X4 U4651 ( .A(n8467), .B(\u_DataPath/pc_4_to_ex_i [4]), .Z(
        n5704) );
  HS65_LH_CNIVX3 U4652 ( .A(\u_DataPath/pc_4_to_ex_i [17]), .Z(n7426) );
  HS65_LH_IVX4 U4653 ( .A(\u_DataPath/dataOut_exe_i [8]), .Z(n3027) );
  HS65_LH_CNIVX3 U4654 ( .A(\u_DataPath/pc_4_to_ex_i [2]), .Z(
        \u_DataPath/u_execute/link_value_i [2]) );
  HS65_LH_NAND2X5 U4655 ( .A(\u_DataPath/pc_4_to_ex_i [17]), .B(
        \u_DataPath/pc_4_to_ex_i [16]), .Z(n6753) );
  HS65_LH_NAND2X5 U4656 ( .A(n8474), .B(\u_DataPath/pc_4_to_ex_i [7]), .Z(
        n5697) );
  HS65_LH_NAND2X4 U4658 ( .A(n8500), .B(\u_DataPath/u_execute/link_value_i [0]), .Z(n5664) );
  HS65_LH_CNIVX3 U4659 ( .A(\u_DataPath/pc_4_to_ex_i [4]), .Z(n7416) );
  HS65_LH_NAND2X5 U4662 ( .A(\u_DataPath/idex_rt_i [2]), .B(
        \u_DataPath/pc_4_to_ex_i [18]), .Z(n5877) );
  HS65_LH_CNIVX3 U4663 ( .A(\u_DataPath/pc_4_to_ex_i [14]), .Z(n7438) );
  HS65_LH_NOR2X6 U4664 ( .A(n8512), .B(\u_DataPath/pc_4_to_ex_i [15]), .Z(
        n5567) );
  HS65_LL_OAI12X3 U4673 ( .A(n9044), .B(n8756), .C(n8283), .Z(
        \u_DataPath/dataOut_exe_i [22]) );
  HS65_LL_OAI12X3 U4674 ( .A(n9044), .B(n8765), .C(n8588), .Z(
        \u_DataPath/dataOut_exe_i [31]) );
  HS65_LL_OAI12X3 U4677 ( .A(n9044), .B(n8746), .C(n8241), .Z(
        \u_DataPath/dataOut_exe_i [18]) );
  HS65_LL_NAND2X4 U4678 ( .A(n3711), .B(n3710), .Z(n8353) );
  HS65_LL_OAI12X3 U4679 ( .A(n8310), .B(n8347), .C(n8229), .Z(
        \u_DataPath/dataOut_exe_i [8]) );
  HS65_LL_OAI112X1 U4691 ( .A(n4695), .B(n4694), .C(n2835), .D(n4693), .Z(
        n4696) );
  HS65_LL_AO12X4 U4694 ( .A(n4723), .B(n4732), .C(n4729), .Z(n3456) );
  HS65_LL_IVX2 U4701 ( .A(n4996), .Z(n5175) );
  HS65_LH_NOR2AX3 U4703 ( .A(n5486), .B(n4813), .Z(n4814) );
  HS65_LH_NAND2X4 U4707 ( .A(n4080), .B(n3905), .Z(n3907) );
  HS65_LL_AOI22X1 U4711 ( .A(n4667), .B(n4831), .C(n4851), .D(n4294), .Z(n4252) );
  HS65_LH_AOI21X2 U4714 ( .A(n5505), .B(n4780), .C(n4779), .Z(n4788) );
  HS65_LHS_XNOR2X6 U4725 ( .A(n3681), .B(n3680), .Z(n3709) );
  HS65_LL_NOR3X1 U4735 ( .A(n5211), .B(n4147), .C(n4146), .Z(n3873) );
  HS65_LH_NAND2X4 U4741 ( .A(n4743), .B(n4466), .Z(n4470) );
  HS65_LH_IVX9 U4749 ( .A(n3865), .Z(n4281) );
  HS65_LH_NAND2X4 U4750 ( .A(n5426), .B(n4237), .Z(n4243) );
  HS65_LH_IVX7 U4754 ( .A(n4682), .Z(n4414) );
  HS65_LH_NOR2X3 U4759 ( .A(n5341), .B(n5342), .Z(n5418) );
  HS65_LH_IVX9 U4760 ( .A(n4292), .Z(n5505) );
  HS65_LL_AOI21X2 U4761 ( .A(n3900), .B(n3263), .C(n3262), .Z(n3264) );
  HS65_LH_NAND2X7 U4767 ( .A(n4325), .B(n4324), .Z(n3696) );
  HS65_LL_CNIVX3 U4768 ( .A(n3636), .Z(n3157) );
  HS65_LL_NAND3X2 U4777 ( .A(n5051), .B(n5027), .C(n4912), .Z(n4906) );
  HS65_LH_IVX9 U4784 ( .A(n5132), .Z(n4551) );
  HS65_LH_AOI21X2 U4785 ( .A(n4257), .B(n4260), .C(n3677), .Z(n3678) );
  HS65_LH_NAND2X7 U4793 ( .A(n5455), .B(n5453), .Z(n5281) );
  HS65_LH_OAI21X3 U4807 ( .A(n2788), .B(n4846), .C(n4621), .Z(n3910) );
  HS65_LH_NOR2X6 U4809 ( .A(n3297), .B(n3296), .Z(n4111) );
  HS65_LL_NOR2X2 U4810 ( .A(n4804), .B(n4799), .Z(n3253) );
  HS65_LH_NAND2X7 U4811 ( .A(n5354), .B(n5388), .Z(n5373) );
  HS65_LH_NOR2X6 U4819 ( .A(n4283), .B(n5201), .Z(n5335) );
  HS65_LH_NAND2X7 U4820 ( .A(n3629), .B(n3628), .Z(n3923) );
  HS65_LH_NAND2X7 U4821 ( .A(n3103), .B(n3106), .Z(n5455) );
  HS65_LH_NOR2X6 U4827 ( .A(n3978), .B(n3977), .Z(n5255) );
  HS65_LL_IVX9 U4834 ( .A(n3251), .Z(n2995) );
  HS65_LH_IVX9 U4835 ( .A(n5436), .Z(n5444) );
  HS65_LL_IVX7 U4839 ( .A(n5067), .Z(n3200) );
  HS65_LH_IVX9 U4840 ( .A(n3330), .Z(n4324) );
  HS65_LH_NOR2X5 U4841 ( .A(\lte_x_57/B[3] ), .B(n3251), .Z(n4799) );
  HS65_LH_NAND2X7 U4842 ( .A(n2780), .B(n5508), .Z(n5490) );
  HS65_LH_OAI12X3 U4847 ( .A(n3901), .B(n3896), .C(n3898), .Z(n3262) );
  HS65_LL_NOR2X3 U4849 ( .A(\lte_x_57/B[7] ), .B(n5207), .Z(n4347) );
  HS65_LH_AOI22X1 U4852 ( .A(n5192), .B(n3826), .C(n2796), .D(\sub_x_51/A[22] ), .Z(n3829) );
  HS65_LL_NOR2X3 U4853 ( .A(\sub_x_51/A[5] ), .B(n2787), .Z(n3765) );
  HS65_LL_NOR2X3 U4860 ( .A(n4718), .B(n4727), .Z(n3269) );
  HS65_LL_AOI13X2 U4861 ( .A(n3379), .B(n4653), .C(n4652), .D(n5148), .Z(n4654) );
  HS65_LH_IVX9 U4863 ( .A(n5011), .Z(n5437) );
  HS65_LH_NAND2X7 U4865 ( .A(n5072), .B(n5016), .Z(n5452) );
  HS65_LL_NOR2X3 U4866 ( .A(n7317), .B(n3239), .Z(n5014) );
  HS65_LH_NOR2X5 U4868 ( .A(n5393), .B(n2829), .Z(n3341) );
  HS65_LH_IVX9 U4870 ( .A(n8141), .Z(\u_DataPath/jump_address_i [21]) );
  HS65_LH_NAND2X7 U4873 ( .A(n8431), .B(n3143), .Z(n3144) );
  HS65_LH_OA12X4 U4874 ( .A(n8657), .B(n7646), .C(n8453), .Z(
        \u_DataPath/mem_writedata_out_i [31]) );
  HS65_LH_NAND2X4 U4878 ( .A(\lte_x_57/B[25] ), .B(n4796), .Z(n3407) );
  HS65_LH_CBI4I1X3 U4879 ( .A(n2802), .B(n5252), .C(n5506), .D(
        \add_x_50/A[23] ), .Z(n4751) );
  HS65_LH_NAND2X7 U4881 ( .A(n4901), .B(n4902), .Z(n5453) );
  HS65_LH_IVX9 U4882 ( .A(n8171), .Z(\u_DataPath/jump_address_i [11]) );
  HS65_LL_NAND2X4 U4883 ( .A(n3160), .B(n5252), .Z(n5284) );
  HS65_LH_NOR2X6 U4884 ( .A(n4032), .B(n2829), .Z(n3860) );
  HS65_LH_NAND2X5 U4885 ( .A(\lte_x_57/B[14] ), .B(n2792), .Z(n3682) );
  HS65_LH_IVX9 U4887 ( .A(n5084), .Z(n2788) );
  HS65_LH_IVX9 U4888 ( .A(n8143), .Z(\u_DataPath/jump_address_i [20]) );
  HS65_LL_NAND2X4 U4889 ( .A(n2793), .B(n4208), .Z(n3851) );
  HS65_LH_NAND2X4 U4892 ( .A(\u_DataPath/u_execute/A_inALU_i[26] ), .B(n2792), 
        .Z(n3628) );
  HS65_LH_OA12X4 U4894 ( .A(n8682), .B(n7646), .C(n8446), .Z(
        \u_DataPath/mem_writedata_out_i [25]) );
  HS65_LH_OAI22X4 U4895 ( .A(n7302), .B(n7903), .C(n7698), .D(n8203), .Z(
        \u_DataPath/data_read_ex_1_i [21]) );
  HS65_LH_OAI22X4 U4896 ( .A(n6861), .B(n7746), .C(n7716), .D(n8039), .Z(
        \u_DataPath/data_read_ex_2_i [31]) );
  HS65_LH_OAI22X4 U4897 ( .A(n7302), .B(n7777), .C(n7698), .D(n8168), .Z(
        \u_DataPath/data_read_ex_1_i [13]) );
  HS65_LH_AOI22X6 U4898 ( .A(\sub_x_51/A[20] ), .B(n7679), .C(n7681), .D(
        \u_DataPath/u_execute/resAdd1_i [20]), .Z(n8143) );
  HS65_LH_AOI22X6 U4900 ( .A(\sub_x_51/A[21] ), .B(n7679), .C(n7681), .D(
        \u_DataPath/u_execute/resAdd1_i [21]), .Z(n8141) );
  HS65_LH_AOI22X6 U4901 ( .A(\lte_x_57/B[11] ), .B(n7679), .C(n7681), .D(
        \u_DataPath/u_execute/resAdd1_i [11]), .Z(n8171) );
  HS65_LH_IVX9 U4902 ( .A(n8136), .Z(\u_DataPath/jump_address_i [25]) );
  HS65_LH_NOR2X2 U4904 ( .A(rst), .B(n8448), .Z(
        \u_DataPath/mem_writedata_out_i [27]) );
  HS65_LH_IVX9 U4905 ( .A(n8169), .Z(\u_DataPath/jump_address_i [13]) );
  HS65_LL_OAI12X6 U4907 ( .A(n8415), .B(n3051), .C(n3050), .Z(n5392) );
  HS65_LH_NAND2X7 U4911 ( .A(n9291), .B(n2797), .Z(n8394) );
  HS65_LL_OAI12X3 U4912 ( .A(n9149), .B(n5565), .C(n9026), .Z(n5721) );
  HS65_LH_NOR2X5 U4916 ( .A(n8681), .B(n2772), .Z(n8439) );
  HS65_LL_IVX7 U4917 ( .A(\lte_x_57/B[14] ), .Z(n5393) );
  HS65_LH_AOI22X6 U4921 ( .A(\lte_x_57/B[25] ), .B(n7680), .C(n7682), .D(
        \u_DataPath/u_execute/resAdd1_i [25]), .Z(n8136) );
  HS65_LL_OAI21X2 U4922 ( .A(n8651), .B(n2772), .C(n3120), .Z(n8449) );
  HS65_LH_AOI22X6 U4923 ( .A(\sub_x_51/A[13] ), .B(n7679), .C(n7681), .D(
        \u_DataPath/u_execute/resAdd1_i [13]), .Z(n8169) );
  HS65_LL_IVX7 U4924 ( .A(\lte_x_57/B[30] ), .Z(n5311) );
  HS65_LHS_XNOR2X3 U4926 ( .A(n9215), .B(n7303), .Z(
        \u_DataPath/u_execute/link_value_i [26]) );
  HS65_LH_CNIVX3 U4927 ( .A(\u_DataPath/u_idexreg/N15 ), .Z(n8024) );
  HS65_LH_CNIVX3 U4928 ( .A(\u_DataPath/u_idexreg/N16 ), .Z(n8025) );
  HS65_LH_AO22X9 U4930 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][26] ), .B(n9254), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][26] ), .D(
        n9244), .Z(n6795) );
  HS65_LH_IVX9 U4933 ( .A(n7947), .Z(n7948) );
  HS65_LL_NOR2X6 U4934 ( .A(n2985), .B(n2984), .Z(\lte_x_57/B[3] ) );
  HS65_LL_AO112X4 U4935 ( .A(n8699), .B(n2710), .C(n3053), .D(n3052), .Z(n3054) );
  HS65_LL_NOR2X6 U4937 ( .A(n3047), .B(n3046), .Z(\lte_x_57/B[14] ) );
  HS65_LL_NOR2X3 U4940 ( .A(n7606), .B(n7605), .Z(n7456) );
  HS65_LH_AOI22X3 U4942 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][21] ), .B(n9247), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][21] ), .D(
        n9227), .Z(n6002) );
  HS65_LH_AO22X4 U4944 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][10] ), .B(n9258), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][10] ), .D(
        n9245), .Z(n7040) );
  HS65_LH_AOI22X3 U4949 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][17] ), .B(n9248), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][17] ), .D(
        n9240), .Z(n6369) );
  HS65_LH_AOI22X3 U4950 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][21] ), .B(n9248), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][21] ), .D(
        n9240), .Z(n6389) );
  HS65_LH_AOI22X3 U4951 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][17] ), .B(n9247), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][17] ), .D(
        n9227), .Z(n5953) );
  HS65_LH_AOI22X3 U4952 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][15] ), .B(n8851), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][15] ), .D(
        n9264), .Z(n6892) );
  HS65_LH_AO22X4 U4954 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][31] ), .B(n9199), 
        .C(n9158), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][31] ), .Z(n7496)
         );
  HS65_LH_AO22X4 U4955 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][14] ), .B(n9258), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][14] ), .D(
        n9245), .Z(n6084) );
  HS65_LH_AO22X9 U4956 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][9] ), .B(n9254), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][9] ), .D(
        n9244), .Z(n7070) );
  HS65_LH_AOI22X3 U4960 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][16] ), .B(n9246), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][16] ), .D(
        n9067), .Z(n6177) );
  HS65_LH_AO22X9 U4964 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][12] ), .B(n9206), 
        .C(n9205), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][12] ), .Z(n7137)
         );
  HS65_LH_AO22X9 U4965 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][12] ), .B(n9204), 
        .C(n9203), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][12] ), .Z(n7136)
         );
  HS65_LH_AOI22X3 U4966 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][19] ), .B(n9259), 
        .C(n9256), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][19] ), .Z(n6770)
         );
  HS65_LH_AO22X4 U4967 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][19] ), .B(n9258), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][19] ), .D(
        n9245), .Z(n6765) );
  HS65_LH_AOI22X3 U4970 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][5] ), .B(n9159), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][5] ), .D(n9265), .Z(n7089) );
  HS65_LH_AO22X9 U4972 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][5] ), .B(n9254), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][5] ), .D(
        n9244), .Z(n7090) );
  HS65_LH_AOI22X3 U4973 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][14] ), .B(n9188), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][14] ), .D(
        n9190), .Z(n6868) );
  HS65_LH_AOI22X3 U4974 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][13] ), .B(n8950), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][13] ), .D(
        n9471), .Z(n6404) );
  HS65_LH_AO22X9 U4975 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][27] ), .B(n9187), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][27] ), .D(
        n8852), .Z(n6313) );
  HS65_LH_AOI22X3 U4980 ( .A(n7679), .B(\sub_x_51/A[8] ), .C(n7681), .D(
        \u_DataPath/u_execute/resAdd1_i [8]), .Z(n8174) );
  HS65_LH_IVX7 U4986 ( .A(n8087), .Z(\u_DataPath/pc4_to_idexreg_i [24]) );
  HS65_LH_IVX7 U4987 ( .A(n8090), .Z(\u_DataPath/pc4_to_idexreg_i [22]) );
  HS65_LH_IVX7 U4988 ( .A(n8093), .Z(\u_DataPath/pc4_to_idexreg_i [20]) );
  HS65_LH_IVX7 U4989 ( .A(n8095), .Z(\u_DataPath/pc4_to_idexreg_i [19]) );
  HS65_LH_IVX7 U4990 ( .A(n8105), .Z(\u_DataPath/pc4_to_idexreg_i [13]) );
  HS65_LH_IVX7 U4993 ( .A(n8513), .Z(n8363) );
  HS65_LH_NOR2X6 U4994 ( .A(n2924), .B(n2794), .Z(n8387) );
  HS65_LH_NOR2X5 U4995 ( .A(n8672), .B(n3181), .Z(n3101) );
  HS65_LH_NOR2X6 U4996 ( .A(n3139), .B(n2794), .Z(n8421) );
  HS65_LH_NOR2X6 U4997 ( .A(n3131), .B(n2794), .Z(n8423) );
  HS65_LH_AOI22X3 U4999 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][4] ), .B(n9248), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][4] ), .D(
        n9240), .Z(n6429) );
  HS65_LH_AOI22X3 U5000 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][4] ), .B(n8851), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][4] ), .D(n9264), .Z(n6426) );
  HS65_LH_AOI22X3 U5003 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][2] ), .B(n9248), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][2] ), .D(
        n9240), .Z(n6229) );
  HS65_LH_AOI211X2 U5004 ( .A(n8721), .B(n2798), .C(n8444), .D(rst), .Z(n8446)
         );
  HS65_LH_NOR2X5 U5010 ( .A(n8677), .B(n3149), .Z(n2953) );
  HS65_LH_AOI21X2 U5011 ( .A(n8741), .B(n2798), .C(n3113), .Z(n3114) );
  HS65_LL_IVX4 U5018 ( .A(n3214), .Z(n2904) );
  HS65_LHS_XOR2X3 U5019 ( .A(n8912), .B(n5790), .Z(
        \u_DataPath/u_execute/resAdd1_i [12]) );
  HS65_LL_OAI12X3 U5020 ( .A(n9126), .B(n5641), .C(n9032), .Z(n5725) );
  HS65_LH_NOR2X5 U5022 ( .A(n3174), .B(n8426), .Z(n3154) );
  HS65_LH_BFX9 U5027 ( .A(n7709), .Z(n7705) );
  HS65_LHS_XNOR2X3 U5028 ( .A(n9290), .B(n7441), .Z(
        \u_DataPath/u_execute/link_value_i [20]) );
  HS65_LH_NOR2X2 U5031 ( .A(rst), .B(n2820), .Z(
        \u_DataPath/u_decode_unit/hdu_0/current_state [1]) );
  HS65_LH_IVX7 U5035 ( .A(n8179), .Z(\u_DataPath/branch_target_i [3]) );
  HS65_LH_NAND2X7 U5037 ( .A(n7693), .B(
        \u_DataPath/u_execute/link_value_i [10]), .Z(n8233) );
  HS65_LL_OAI12X3 U5038 ( .A(n5550), .B(n5611), .C(n5549), .Z(n5717) );
  HS65_LH_NAND2X7 U5039 ( .A(n7693), .B(n9381), .Z(n8286) );
  HS65_LH_BFX18 U5040 ( .A(n6111), .Z(n7516) );
  HS65_LL_NOR2X2 U5041 ( .A(n3174), .B(n8414), .Z(n3049) );
  HS65_LL_AOI21X2 U5043 ( .A(n8934), .B(n5572), .C(n5545), .Z(n5611) );
  HS65_LL_NOR2X6 U5044 ( .A(n2917), .B(n2916), .Z(n2988) );
  HS65_LH_BFX18 U5045 ( .A(n6127), .Z(n7586) );
  HS65_LL_NAND3X5 U5046 ( .A(n2888), .B(n2889), .C(n2887), .Z(n2885) );
  HS65_LL_NOR2X5 U5050 ( .A(n5961), .B(n5957), .Z(n6119) );
  HS65_LL_NOR2X5 U5051 ( .A(n5958), .B(n5962), .Z(n6120) );
  HS65_LL_NOR2X5 U5052 ( .A(n5959), .B(n5937), .Z(n6101) );
  HS65_LHS_XOR2X3 U5053 ( .A(n7447), .B(n7446), .Z(\u_DataPath/pc_4_i [6]) );
  HS65_LL_NOR2X5 U5054 ( .A(n5961), .B(n5937), .Z(n6100) );
  HS65_LL_NOR2X5 U5055 ( .A(n7422), .B(n6756), .Z(n7439) );
  HS65_LL_NOR2X5 U5056 ( .A(n5961), .B(n5962), .Z(n6128) );
  HS65_LH_NAND2X5 U5057 ( .A(n1885), .B(n8159), .Z(n8282) );
  HS65_LL_NOR2X5 U5058 ( .A(n5958), .B(n5937), .Z(n6102) );
  HS65_LL_NOR2X5 U5059 ( .A(n5963), .B(n5951), .Z(n7588) );
  HS65_LH_NAND2X4 U5060 ( .A(n8158), .B(n1885), .Z(n8055) );
  HS65_LL_IVX4 U5062 ( .A(n8041), .Z(n2960) );
  HS65_LL_NOR2X5 U5063 ( .A(n2866), .B(n8041), .Z(n2888) );
  HS65_LH_IVX4 U5066 ( .A(n7342), .Z(n7446) );
  HS65_LH_NAND3X5 U5067 ( .A(\u_DataPath/cw_tomem_i [5]), .B(n3438), .C(n7352), 
        .Z(n2805) );
  HS65_LH_NAND2X7 U5068 ( .A(n7417), .B(n6752), .Z(n7422) );
  HS65_LL_NAND4ABX6 U5069 ( .A(n2903), .B(n2770), .C(n2908), .D(n2902), .Z(
        n3048) );
  HS65_LH_IVX9 U5070 ( .A(n3219), .Z(n3220) );
  HS65_LH_NAND2X7 U5071 ( .A(n2811), .B(n6163), .Z(n6162) );
  HS65_LH_CNIVX3 U5073 ( .A(n8082), .Z(\u_DataPath/pc_4_to_ex_i [28]) );
  HS65_LH_IVX4 U5074 ( .A(n8036), .Z(n8512) );
  HS65_LH_CNIVX3 U5075 ( .A(n8106), .Z(\u_DataPath/pc_4_to_ex_i [13]) );
  HS65_LH_CNIVX3 U5076 ( .A(n8107), .Z(\u_DataPath/pc_4_to_ex_i [12]) );
  HS65_LH_CNIVX3 U5077 ( .A(n8108), .Z(\u_DataPath/pc_4_to_ex_i [11]) );
  HS65_LH_CNIVX3 U5078 ( .A(n8110), .Z(\u_DataPath/pc_4_to_ex_i [10]) );
  HS65_LH_CNIVX3 U5079 ( .A(n8111), .Z(\u_DataPath/pc_4_to_ex_i [9]) );
  HS65_LH_CNIVX3 U5080 ( .A(n8113), .Z(\u_DataPath/pc_4_to_ex_i [8]) );
  HS65_LH_CNIVX3 U5081 ( .A(n8115), .Z(\u_DataPath/pc_4_to_ex_i [7]) );
  HS65_LH_CNIVX3 U5082 ( .A(n8116), .Z(\u_DataPath/pc_4_to_ex_i [6]) );
  HS65_LH_CNIVX3 U5083 ( .A(n8080), .Z(\u_DataPath/pc_4_to_ex_i [29]) );
  HS65_LH_CNIVX3 U5084 ( .A(n8083), .Z(\u_DataPath/pc_4_to_ex_i [27]) );
  HS65_LH_CNIVX3 U5085 ( .A(n8079), .Z(\u_DataPath/pc_4_to_ex_i [30]) );
  HS65_LH_CNIVX3 U5086 ( .A(n8185), .Z(\u_DataPath/pc_4_to_ex_i [31]) );
  HS65_LH_CNIVX3 U5087 ( .A(n8085), .Z(\u_DataPath/pc_4_to_ex_i [26]) );
  HS65_LH_CNIVX3 U5088 ( .A(n8086), .Z(\u_DataPath/pc_4_to_ex_i [25]) );
  HS65_LH_CNIVX3 U5089 ( .A(n8088), .Z(\u_DataPath/pc_4_to_ex_i [24]) );
  HS65_LH_CNIVX3 U5090 ( .A(n8089), .Z(\u_DataPath/pc_4_to_ex_i [23]) );
  HS65_LH_CNIVX3 U5091 ( .A(n8091), .Z(\u_DataPath/pc_4_to_ex_i [22]) );
  HS65_LH_CNIVX3 U5092 ( .A(n8129), .Z(\u_DataPath/jump_i ) );
  HS65_LH_CNIVX3 U5093 ( .A(n8360), .Z(\u_DataPath/cw_tomem_i [0]) );
  HS65_LH_CNIVX3 U5094 ( .A(n8092), .Z(\u_DataPath/pc_4_to_ex_i [21]) );
  HS65_LH_CNIVX3 U5095 ( .A(n8032), .Z(\u_DataPath/cw_tomem_i [8]) );
  HS65_LH_CNIVX3 U5096 ( .A(n8033), .Z(\u_DataPath/cw_tomem_i [6]) );
  HS65_LH_CNIVX3 U5097 ( .A(n8094), .Z(\u_DataPath/pc_4_to_ex_i [20]) );
  HS65_LH_CNIVX3 U5098 ( .A(n8117), .Z(\u_DataPath/pc_4_to_ex_i [5]) );
  HS65_LH_CNIVX3 U5099 ( .A(n8096), .Z(\u_DataPath/pc_4_to_ex_i [19]) );
  HS65_LH_CNIVX3 U5100 ( .A(n8097), .Z(\u_DataPath/pc_4_to_ex_i [18]) );
  HS65_LH_CNIVX3 U5101 ( .A(n8099), .Z(\u_DataPath/pc_4_to_ex_i [17]) );
  HS65_LH_CNIVX3 U5102 ( .A(n8100), .Z(\u_DataPath/pc_4_to_ex_i [16]) );
  HS65_LH_CNIVX3 U5103 ( .A(n8048), .Z(\u_DataPath/cw_memwb_i [0]) );
  HS65_LH_CNIVX3 U5104 ( .A(n8102), .Z(\u_DataPath/pc_4_to_ex_i [15]) );
  HS65_LH_CNIVX3 U5105 ( .A(n8104), .Z(\u_DataPath/pc_4_to_ex_i [14]) );
  HS65_LH_CNIVX3 U5106 ( .A(n8124), .Z(\u_DataPath/u_execute/link_value_i [1])
         );
  HS65_LH_CNIVX3 U5107 ( .A(n8121), .Z(\u_DataPath/pc_4_to_ex_i [3]) );
  HS65_LH_NAND2X4 U5108 ( .A(n5876), .B(n5875), .Z(n5881) );
  HS65_LL_NOR2X3 U5109 ( .A(n2901), .B(n2900), .Z(n2902) );
  HS65_LL_NAND2X7 U5110 ( .A(n2871), .B(n7672), .Z(n7014) );
  HS65_LH_AOI12X6 U5111 ( .A(n5794), .B(n5749), .C(n5748), .Z(n5827) );
  HS65_LH_IVX7 U5112 ( .A(n5778), .Z(n5779) );
  HS65_LH_NAND2X5 U5114 ( .A(n8280), .B(n8310), .Z(n7667) );
  HS65_LL_NAND2X7 U5116 ( .A(n2816), .B(\u_DataPath/jaddr_i [22]), .Z(n6186)
         );
  HS65_LH_NAND2X4 U5117 ( .A(n5569), .B(n5568), .Z(n5580) );
  HS65_LL_NAND2X2 U5118 ( .A(n3184), .B(n9429), .Z(n3033) );
  HS65_LH_NOR2X6 U5119 ( .A(\u_DataPath/immediate_ext_dec_i [1]), .B(n8051), 
        .Z(n7990) );
  HS65_LH_NAND2X4 U5120 ( .A(n5697), .B(n5696), .Z(n5702) );
  HS65_LH_IVX7 U5121 ( .A(n7412), .Z(n7413) );
  HS65_LL_NAND3X5 U5122 ( .A(\u_DataPath/jaddr_i [20]), .B(n2804), .C(n8016), 
        .Z(n5950) );
  HS65_LH_NAND2X7 U5123 ( .A(opcode_i[3]), .B(n7965), .Z(n7333) );
  HS65_LH_NOR2X6 U5124 ( .A(n7360), .B(n7355), .Z(n7368) );
  HS65_LH_CNIVX3 U5125 ( .A(n8123), .Z(\u_DataPath/pc4_to_idexreg_i [1]) );
  HS65_LH_CNIVX3 U5127 ( .A(n8125), .Z(\u_DataPath/pc4_to_idexreg_i [0]) );
  HS65_LH_NOR2X2 U5128 ( .A(n7710), .B(n9285), .Z(\u_DataPath/cw_tomem_i [5])
         );
  HS65_LH_IVX9 U5129 ( .A(\u_DataPath/jaddr_i [16]), .Z(n5935) );
  HS65_LH_NOR2X6 U5130 ( .A(n5616), .B(n5619), .Z(n5626) );
  HS65_LH_NOR2X6 U5131 ( .A(n6751), .B(n7435), .Z(n6752) );
  HS65_LH_IVX4 U5132 ( .A(n5789), .Z(n5814) );
  HS65_LL_NAND2X2 U5134 ( .A(n2905), .B(n2907), .Z(n2900) );
  HS65_LL_IVX2 U5135 ( .A(n2906), .Z(n2901) );
  HS65_LH_IVX4 U5136 ( .A(n5592), .Z(n5684) );
  HS65_LH_NOR2X5 U5137 ( .A(n8466), .B(\u_DataPath/pc_4_to_ex_i [3]), .Z(n5910) );
  HS65_LH_NOR2X2 U5138 ( .A(n9268), .B(rst), .Z(\u_DataPath/u_memwbreg/N45 )
         );
  HS65_LH_IVX7 U5139 ( .A(\u_DataPath/data_read_ex_1_i [24]), .Z(n3096) );
  HS65_LH_NOR3X3 U5140 ( .A(\u_DataPath/cw_to_ex_i [17]), .B(
        \u_DataPath/cw_exmem_i [9]), .C(\u_DataPath/cw_to_ex_i [15]), .Z(n8155) );
  HS65_LH_CNIVX3 U5141 ( .A(\u_DataPath/pc_4_to_ex_i [6]), .Z(n7617) );
  HS65_LH_IVX9 U5142 ( .A(\u_DataPath/idex_rt_i [1]), .Z(n2893) );
  HS65_LH_NAND2X4 U5143 ( .A(n8498), .B(\u_DataPath/u_execute/link_value_i [1]), .Z(n5662) );
  HS65_LH_NAND2X4 U5144 ( .A(n8465), .B(\u_DataPath/pc_4_to_ex_i [2]), .Z(
        n5710) );
  HS65_LH_IVX7 U5145 ( .A(n8526), .Z(n3981) );
  HS65_LH_NOR2X3 U5147 ( .A(n8465), .B(\u_DataPath/pc_4_to_ex_i [2]), .Z(n5712) );
  HS65_LH_CNIVX3 U5149 ( .A(\u_DataPath/pc_4_to_ex_i [8]), .Z(n7436) );
  HS65_LH_IVX7 U5150 ( .A(\u_DataPath/data_read_ex_1_i [8]), .Z(n3025) );
  HS65_LH_IVX9 U5151 ( .A(n7673), .Z(n7216) );
  HS65_LH_IVX18 U5152 ( .A(n7672), .Z(n7013) );
  HS65_LH_CNIVX3 U5153 ( .A(\u_DataPath/pc_4_to_ex_i [12]), .Z(n7630) );
  HS65_LH_NAND2X7 U5155 ( .A(\u_DataPath/rs_ex_i [0]), .B(
        \u_DataPath/pc_4_to_ex_i [21]), .Z(n5818) );
  HS65_LH_IVX9 U5157 ( .A(\u_DataPath/data_read_ex_2_i [12]), .Z(n8409) );
  HS65_LH_NAND2X7 U5158 ( .A(\u_DataPath/pc_4_to_ex_i [11]), .B(
        \u_DataPath/pc_4_to_ex_i [10]), .Z(n7431) );
  HS65_LH_NAND2X7 U5159 ( .A(\u_DataPath/pc_4_to_ex_i [15]), .B(
        \u_DataPath/pc_4_to_ex_i [14]), .Z(n7421) );
  HS65_LH_NAND2X7 U5161 ( .A(\u_DataPath/pc_4_to_ex_i [19]), .B(
        \u_DataPath/pc_4_to_ex_i [18]), .Z(n7440) );
  HS65_LH_IVX9 U5163 ( .A(\u_DataPath/u_decode_unit/hdu_0/current_state [0]), 
        .Z(n7196) );
  HS65_LH_IVX7 U5164 ( .A(\u_DataPath/data_read_ex_1_i [19]), .Z(n3145) );
  HS65_LH_NAND2X7 U5165 ( .A(n8596), .B(n9124), .Z(
        \u_DataPath/dataOut_exe_i [29]) );
  HS65_LH_IVX9 U5167 ( .A(n8214), .Z(\u_DataPath/dataOut_exe_i [11]) );
  HS65_LL_NAND2AX4 U5169 ( .A(n4550), .B(n4549), .Z(n8326) );
  HS65_LH_AOI22X6 U5170 ( .A(\u_DataPath/u_execute/link_value_i [11]), .B(
        n7695), .C(n8315), .D(n8353), .Z(n8214) );
  HS65_LL_OAI21X3 U5171 ( .A(n4591), .B(n9539), .C(n4589), .Z(n8327) );
  HS65_LL_NOR2AX3 U5173 ( .A(n4588), .B(n4587), .Z(n4589) );
  HS65_LL_NAND4ABX3 U5174 ( .A(n5176), .B(n5175), .C(n5061), .D(n5174), .Z(
        n8325) );
  HS65_LL_AOI21X2 U5182 ( .A(n5492), .B(n3709), .C(n3708), .Z(n3710) );
  HS65_LL_NOR2AX3 U5185 ( .A(n5058), .B(n5057), .Z(n5059) );
  HS65_LL_NAND2X2 U5187 ( .A(n4089), .B(n4088), .Z(n4099) );
  HS65_LH_IVX9 U5189 ( .A(n4856), .Z(n4857) );
  HS65_LLS_XNOR2X3 U5191 ( .A(n4697), .B(n4696), .Z(n7320) );
  HS65_LLS_XNOR2X3 U5193 ( .A(n3544), .B(n3543), .Z(n3552) );
  HS65_LLS_XNOR2X3 U5194 ( .A(n4547), .B(n4546), .Z(n4548) );
  HS65_LL_AOI21X2 U5196 ( .A(n5173), .B(n2850), .C(n5172), .Z(n5174) );
  HS65_LL_NOR3X1 U5200 ( .A(n4201), .B(n4200), .C(n4199), .Z(n4233) );
  HS65_LL_NOR2X2 U5201 ( .A(n4516), .B(n4515), .Z(n4517) );
  HS65_LL_NOR2X2 U5202 ( .A(n4072), .B(n4071), .Z(n4073) );
  HS65_LL_OAI12X2 U5206 ( .A(n4744), .B(n4468), .C(n4029), .Z(n4037) );
  HS65_LL_OAI22X1 U5207 ( .A(n4747), .B(n4746), .C(n4745), .D(n4744), .Z(n4755) );
  HS65_LH_NOR2X5 U5211 ( .A(n4502), .B(n3321), .Z(n3333) );
  HS65_LL_NOR2X2 U5214 ( .A(n3632), .B(n3631), .Z(n4813) );
  HS65_LH_NAND3X5 U5223 ( .A(n3382), .B(n3381), .C(n3380), .Z(n3395) );
  HS65_LL_AOI22X1 U5226 ( .A(n4294), .B(n4832), .C(n5484), .D(n4828), .Z(n3602) );
  HS65_LH_OAI21X3 U5231 ( .A(n4846), .B(n2791), .C(n4405), .Z(n4406) );
  HS65_LH_NOR3X4 U5234 ( .A(n3931), .B(n3930), .C(n3929), .Z(n3932) );
  HS65_LL_AOI12X2 U5237 ( .A(n5325), .B(n5289), .C(n5365), .Z(n5331) );
  HS65_LL_CBI4I6X2 U5240 ( .A(n2829), .B(n4189), .C(n4188), .D(n5499), .Z(
        n4201) );
  HS65_LH_AOI21X2 U5248 ( .A(n5217), .B(n5216), .C(n5215), .Z(n5225) );
  HS65_LH_NAND2X4 U5249 ( .A(n4618), .B(n4063), .Z(n3380) );
  HS65_LL_AO12X4 U5252 ( .A(n4730), .B(n4729), .C(n4728), .Z(n4731) );
  HS65_LL_AOI12X2 U5253 ( .A(n3883), .B(n4092), .C(n3885), .Z(n3618) );
  HS65_LL_NOR3X1 U5254 ( .A(n4982), .B(n4981), .C(n4980), .Z(n5165) );
  HS65_LL_NAND2X2 U5257 ( .A(n4692), .B(n4691), .Z(n4693) );
  HS65_LH_OAI12X3 U5260 ( .A(n4564), .B(n3337), .C(n3336), .Z(n3352) );
  HS65_LL_OAI12X3 U5261 ( .A(n3003), .B(n3002), .C(n3001), .Z(n3666) );
  HS65_LL_NOR3X1 U5262 ( .A(n4914), .B(n4906), .C(n4923), .Z(n4907) );
  HS65_LL_OAI22X1 U5264 ( .A(n4753), .B(n4332), .C(n4665), .D(n4745), .Z(n3351) );
  HS65_LH_IVX9 U5266 ( .A(n4564), .Z(n4740) );
  HS65_LL_NOR2X2 U5268 ( .A(n4747), .B(n4295), .Z(n4296) );
  HS65_LH_AOI22X3 U5270 ( .A(n5517), .B(n4961), .C(n4743), .D(n4742), .Z(n4756) );
  HS65_LL_OAI12X3 U5271 ( .A(n4176), .B(n3083), .C(n3082), .Z(n3084) );
  HS65_LH_OAI12X3 U5277 ( .A(n3903), .B(n3902), .C(n3901), .Z(n3904) );
  HS65_LH_AOI12X2 U5278 ( .A(n3874), .B(n4822), .C(n3761), .Z(n3762) );
  HS65_LL_CBI4I1X3 U5279 ( .A(n5308), .B(n5307), .C(n5306), .D(n5305), .Z(
        n5326) );
  HS65_LH_NAND2X4 U5281 ( .A(n4168), .B(n4080), .Z(n4084) );
  HS65_LH_NOR2X6 U5292 ( .A(n5198), .B(n5272), .Z(n5275) );
  HS65_LL_NOR2X2 U5304 ( .A(n4177), .B(n3083), .Z(n3071) );
  HS65_LH_OAI12X3 U5306 ( .A(n4523), .B(n4689), .C(n4522), .Z(n4524) );
  HS65_LH_NAND2X7 U5308 ( .A(n1885), .B(\u_DataPath/toPC2_i [31]), .Z(n8130)
         );
  HS65_LH_CNIVX3 U5313 ( .A(n4932), .Z(n4933) );
  HS65_LH_NAND2X7 U5318 ( .A(n3798), .B(n3797), .Z(n4062) );
  HS65_LH_NAND2X4 U5320 ( .A(n4610), .B(n3390), .Z(n3391) );
  HS65_LH_IVX9 U5323 ( .A(n4332), .Z(n4739) );
  HS65_LL_NAND2X2 U5324 ( .A(n3077), .B(n4238), .Z(n4177) );
  HS65_LH_NAND2X4 U5332 ( .A(n5237), .B(n5205), .Z(n5240) );
  HS65_LHS_XOR2X6 U5334 ( .A(n4769), .B(n4186), .Z(n4236) );
  HS65_LH_NOR2X5 U5335 ( .A(n4812), .B(n4321), .Z(n4829) );
  HS65_LH_NAND2X7 U5339 ( .A(n4169), .B(n4168), .Z(n4173) );
  HS65_LL_NOR2X3 U5344 ( .A(n4674), .B(n4613), .Z(n4610) );
  HS65_LL_AOI12X3 U5352 ( .A(n4603), .B(n3273), .C(n3272), .Z(n4689) );
  HS65_LH_IVX7 U5353 ( .A(n4333), .Z(n4334) );
  HS65_LH_IVX7 U5357 ( .A(n4308), .Z(n4780) );
  HS65_LH_NAND2X7 U5359 ( .A(n3787), .B(n3788), .Z(n4477) );
  HS65_LH_NAND2X7 U5361 ( .A(n4258), .B(n4257), .Z(n4264) );
  HS65_LH_IVX9 U5363 ( .A(n4222), .Z(n4851) );
  HS65_LH_AOI21X2 U5364 ( .A(n5301), .B(n5300), .C(n5299), .Z(n5302) );
  HS65_LL_NAND2X2 U5365 ( .A(n3255), .B(n4823), .Z(n3257) );
  HS65_LH_IVX9 U5369 ( .A(n5184), .Z(n4461) );
  HS65_LH_NOR2X6 U5373 ( .A(n3344), .B(n3343), .Z(n4745) );
  HS65_LL_OAI12X2 U5374 ( .A(n5426), .B(n3664), .C(n5228), .Z(n3076) );
  HS65_LH_AOI12X2 U5376 ( .A(n5449), .B(n5448), .C(n5447), .Z(n5473) );
  HS65_LL_OAI12X2 U5378 ( .A(n4374), .B(n3536), .C(n3538), .Z(n3266) );
  HS65_LH_NAND2X7 U5380 ( .A(n1885), .B(\u_DataPath/toPC2_i [29]), .Z(n8133)
         );
  HS65_LL_OAI12X2 U5381 ( .A(n4602), .B(n3353), .C(n3355), .Z(n3272) );
  HS65_LH_NAND2X7 U5382 ( .A(n5269), .B(n5197), .Z(n5272) );
  HS65_LL_NAND3X3 U5383 ( .A(n3488), .B(n3487), .C(n3486), .Z(n4572) );
  HS65_LH_NAND3X3 U5384 ( .A(n3823), .B(n3822), .C(n3821), .Z(n3824) );
  HS65_LH_NOR2X5 U5385 ( .A(n3924), .B(n3923), .Z(n3692) );
  HS65_LL_OAI12X3 U5386 ( .A(n4488), .B(n4486), .C(n4487), .Z(n4724) );
  HS65_LH_NAND2X2 U5389 ( .A(n5412), .B(n5349), .Z(n3947) );
  HS65_LH_AOI21X2 U5393 ( .A(n5295), .B(n4911), .C(n5002), .Z(n4917) );
  HS65_LH_NAND3X3 U5395 ( .A(n5454), .B(n5445), .C(n4011), .Z(n4008) );
  HS65_LH_NAND2X7 U5396 ( .A(n5192), .B(n3200), .Z(n4552) );
  HS65_LH_NOR2X6 U5397 ( .A(n3685), .B(n3684), .Z(n4791) );
  HS65_LH_NOR2X6 U5398 ( .A(n3189), .B(\add_x_50/A[19] ), .Z(n3636) );
  HS65_LH_IVX9 U5400 ( .A(n4079), .Z(n4168) );
  HS65_LH_NAND2X7 U5401 ( .A(\lte_x_57/B[10] ), .B(n3074), .Z(n5426) );
  HS65_LH_NAND2X7 U5404 ( .A(n5263), .B(n4540), .Z(n4547) );
  HS65_LH_NOR2X6 U5413 ( .A(n3586), .B(n3585), .Z(n4222) );
  HS65_LL_OAI12X3 U5414 ( .A(n3875), .B(n3756), .C(n3758), .Z(n4821) );
  HS65_LH_NAND2X4 U5416 ( .A(n5517), .B(n4957), .Z(n4058) );
  HS65_LH_IVX9 U5417 ( .A(n5064), .Z(n3192) );
  HS65_LL_NOR2X2 U5419 ( .A(n4701), .B(n4709), .Z(n3197) );
  HS65_LL_NOR2X2 U5423 ( .A(n5085), .B(n3888), .Z(n3081) );
  HS65_LH_IVX9 U5425 ( .A(n5246), .Z(n3189) );
  HS65_LH_IVX9 U5427 ( .A(n5066), .Z(n3193) );
  HS65_LH_NAND2X7 U5428 ( .A(\lte_x_57/B[11] ), .B(n5077), .Z(n3675) );
  HS65_LL_AOI12X2 U5430 ( .A(n9132), .B(n5868), .C(n9460), .Z(n5758) );
  HS65_LH_NOR2X6 U5431 ( .A(\lte_x_57/B[11] ), .B(n5077), .Z(n3673) );
  HS65_LH_NAND2X7 U5432 ( .A(\lte_x_57/B[10] ), .B(n5386), .Z(n4258) );
  HS65_LH_NOR2X6 U5434 ( .A(n2793), .B(n5203), .Z(n4079) );
  HS65_LH_NAND2X7 U5435 ( .A(\sub_x_51/A[8] ), .B(n5201), .Z(n4277) );
  HS65_LL_NAND2X4 U5436 ( .A(\lte_x_57/B[2] ), .B(n2994), .Z(n4768) );
  HS65_LL_NOR2X2 U5439 ( .A(n4541), .B(n5070), .Z(n4637) );
  HS65_LL_NOR2X5 U5440 ( .A(\lte_x_57/B[6] ), .B(n2998), .Z(n4859) );
  HS65_LH_NAND2X4 U5445 ( .A(n5036), .B(n5350), .Z(n3954) );
  HS65_LH_NOR2X6 U5446 ( .A(n3765), .B(n5209), .Z(n4864) );
  HS65_LL_NAND2X4 U5449 ( .A(n4128), .B(n4127), .Z(n4827) );
  HS65_LL_NAND2X4 U5450 ( .A(n3576), .B(n3575), .Z(n4828) );
  HS65_LL_NAND2X4 U5451 ( .A(n4203), .B(n5077), .Z(n5354) );
  HS65_LH_NAND2X7 U5455 ( .A(n5385), .B(n5386), .Z(n5376) );
  HS65_LH_OAI21X2 U5457 ( .A(n3842), .B(n5218), .C(n3767), .Z(n5222) );
  HS65_LH_OAI12X3 U5458 ( .A(n5265), .B(n5264), .C(n5263), .Z(n5268) );
  HS65_LH_NOR2X6 U5459 ( .A(n5266), .B(n5195), .Z(n5269) );
  HS65_LH_OAI21X2 U5460 ( .A(n5220), .B(n5088), .C(n5219), .Z(n5221) );
  HS65_LH_IVX9 U5465 ( .A(n3633), .Z(n4366) );
  HS65_LH_NOR2X6 U5466 ( .A(\sub_x_51/A[20] ), .B(n5064), .Z(n3453) );
  HS65_LH_NOR2X6 U5467 ( .A(\sub_x_51/A[16] ), .B(n5186), .Z(n4447) );
  HS65_LH_NAND2X5 U5469 ( .A(\lte_x_57/B[11] ), .B(n5496), .Z(n3735) );
  HS65_LL_NAND2X4 U5472 ( .A(n4918), .B(n5066), .Z(n5286) );
  HS65_LH_NAND3X5 U5477 ( .A(n5449), .B(n5437), .C(n5436), .Z(n5456) );
  HS65_LH_NOR2X5 U5481 ( .A(\lte_x_57/B[29] ), .B(n3204), .Z(n5264) );
  HS65_LHS_XOR2X3 U5483 ( .A(n8931), .B(n5560), .Z(\u_DataPath/toPC2_i [28])
         );
  HS65_LH_NOR2X3 U5484 ( .A(\lte_x_57/B[30] ), .B(n2790), .Z(n5195) );
  HS65_LH_NAND2X7 U5485 ( .A(n1885), .B(\u_DataPath/toPC2_i [27]), .Z(n8135)
         );
  HS65_LH_NAND2X7 U5486 ( .A(n4315), .B(n3807), .Z(n3340) );
  HS65_LL_NOR2X3 U5487 ( .A(\sub_x_51/A[22] ), .B(n3194), .Z(n4709) );
  HS65_LL_NOR2X2 U5488 ( .A(n4523), .B(n4519), .Z(n4681) );
  HS65_LH_IVX9 U5489 ( .A(n5079), .Z(n3073) );
  HS65_LH_NAND2X7 U5492 ( .A(n3239), .B(n7317), .Z(n5449) );
  HS65_LH_NAND2X7 U5495 ( .A(\sub_x_51/A[27] ), .B(n4005), .Z(n5009) );
  HS65_LH_AOI21X2 U5497 ( .A(\lte_x_57/B[4] ), .B(n4796), .C(n3844), .Z(n3847)
         );
  HS65_LL_NOR2X3 U5498 ( .A(\add_x_50/A[23] ), .B(n3195), .Z(n4701) );
  HS65_LL_NOR2X2 U5499 ( .A(n5495), .B(n4187), .Z(n4128) );
  HS65_LH_AOI22X1 U5500 ( .A(\sub_x_51/A[20] ), .B(n3826), .C(n2796), .D(
        \sub_x_51/A[18] ), .Z(n3458) );
  HS65_LH_NAND2X4 U5502 ( .A(\u_DataPath/u_execute/A_inALU_i[26] ), .B(n3742), 
        .Z(n3398) );
  HS65_LL_NOR2X3 U5504 ( .A(\u_DataPath/u_execute/A_inALU_i[26] ), .B(n4622), 
        .Z(n4592) );
  HS65_LH_NAND2X7 U5506 ( .A(\u_DataPath/u_execute/A_inALU_i[26] ), .B(n4622), 
        .Z(n4594) );
  HS65_LH_IVX9 U5507 ( .A(n8134), .Z(\u_DataPath/jump_address_i [27]) );
  HS65_LH_NAND2X7 U5509 ( .A(\lte_x_57/B[14] ), .B(n3079), .Z(n3886) );
  HS65_LH_NAND2X7 U5511 ( .A(\lte_x_57/B[30] ), .B(n2790), .Z(n5436) );
  HS65_LH_OR2X9 U5513 ( .A(\lte_x_57/B[30] ), .B(n2790), .Z(n4641) );
  HS65_LL_NOR2X2 U5514 ( .A(n3896), .B(n3903), .Z(n3263) );
  HS65_LH_OAI22X4 U5519 ( .A(n7719), .B(n7854), .C(n7717), .D(n8248), .Z(
        \u_DataPath/data_read_ex_2_i [26]) );
  HS65_LH_OAI22X4 U5520 ( .A(n7719), .B(n7812), .C(n7718), .D(n8271), .Z(
        \u_DataPath/data_read_ex_2_i [30]) );
  HS65_LH_OAI22X4 U5521 ( .A(n7719), .B(n7791), .C(n7717), .D(n8227), .Z(
        \u_DataPath/data_read_ex_2_i [8]) );
  HS65_LH_OAI22X4 U5522 ( .A(n7719), .B(n7826), .C(n7717), .D(n8268), .Z(
        \u_DataPath/data_read_ex_2_i [28]) );
  HS65_LH_NOR2X5 U5526 ( .A(n5084), .B(n3962), .Z(n5366) );
  HS65_LH_OA12X4 U5527 ( .A(n5529), .B(n2830), .C(n3485), .Z(n3487) );
  HS65_LHS_XNOR2X3 U5529 ( .A(n9411), .B(n7307), .Z(
        \u_DataPath/u_execute/link_value_i [28]) );
  HS65_LH_NAND2X4 U5530 ( .A(n3962), .B(n5084), .Z(n3963) );
  HS65_LH_NOR2X5 U5532 ( .A(n3861), .B(n3580), .Z(n3223) );
  HS65_LL_NAND2X4 U5533 ( .A(\sub_x_51/A[22] ), .B(n5251), .Z(n4725) );
  HS65_LL_NOR3X1 U5534 ( .A(n8816), .B(n9051), .C(n7981), .Z(n7953) );
  HS65_LL_NOR2X3 U5535 ( .A(\add_x_50/A[23] ), .B(n5252), .Z(n4718) );
  HS65_LH_IVX7 U5536 ( .A(n3775), .Z(n3776) );
  HS65_LH_AOI22X6 U5540 ( .A(\sub_x_51/A[27] ), .B(n7680), .C(n7682), .D(
        \u_DataPath/u_execute/resAdd1_i [27]), .Z(n8134) );
  HS65_LH_NAND2X5 U5541 ( .A(n4330), .B(n4346), .Z(n5036) );
  HS65_LH_NOR2X3 U5543 ( .A(n3160), .B(n2829), .Z(n3825) );
  HS65_LL_NAND2X2 U5545 ( .A(n8434), .B(n3175), .Z(n3176) );
  HS65_LL_NOR2X3 U5546 ( .A(\lte_x_57/B[28] ), .B(n4902), .Z(n4523) );
  HS65_LH_IVX9 U5552 ( .A(n8078), .Z(\u_DataPath/pc4_to_idexreg_i [30]) );
  HS65_LH_IVX9 U5553 ( .A(n3106), .Z(n4005) );
  HS65_LL_NOR2X3 U5558 ( .A(n2825), .B(n5251), .Z(n5004) );
  HS65_LH_NAND2X4 U5564 ( .A(n3128), .B(n2792), .Z(n3583) );
  HS65_LL_NOR2X2 U5565 ( .A(\lte_x_57/B[14] ), .B(n5392), .Z(n3903) );
  HS65_LH_IVX9 U5566 ( .A(n8150), .Z(\u_DataPath/jump_address_i [15]) );
  HS65_LH_IVX9 U5567 ( .A(n8137), .Z(\u_DataPath/branch_target_i [25]) );
  HS65_LH_OAI22X4 U5568 ( .A(n7719), .B(n7847), .C(n7717), .D(n8208), .Z(
        \u_DataPath/data_read_ex_2_i [23]) );
  HS65_LH_OAI22X4 U5569 ( .A(n7719), .B(n7784), .C(n7717), .D(n8212), .Z(
        \u_DataPath/data_read_ex_2_i [11]) );
  HS65_LH_OAI22X4 U5570 ( .A(n7719), .B(n7739), .C(n7717), .D(n8204), .Z(
        \u_DataPath/data_read_ex_2_i [27]) );
  HS65_LH_OAI22X4 U5571 ( .A(n7719), .B(n7833), .C(n7718), .D(n8269), .Z(
        \u_DataPath/data_read_ex_2_i [29]) );
  HS65_LH_OAI22X4 U5572 ( .A(n7719), .B(n7770), .C(n7717), .D(n8257), .Z(
        \u_DataPath/data_read_ex_2_i [9]) );
  HS65_LH_OAI22X4 U5573 ( .A(n7719), .B(n7910), .C(n7717), .D(n8262), .Z(
        \u_DataPath/data_read_ex_2_i [5]) );
  HS65_LH_OAI22X4 U5574 ( .A(n7719), .B(n7798), .C(n7717), .D(n8244), .Z(
        \u_DataPath/data_read_ex_2_i [6]) );
  HS65_LH_AOI22X4 U5575 ( .A(n2793), .B(n7679), .C(n7681), .D(
        \u_DataPath/u_execute/resAdd1_i [12]), .Z(n8170) );
  HS65_LH_NAND2AX7 U5576 ( .A(n8660), .B(n2797), .Z(n3099) );
  HS65_LH_AOI22X6 U5581 ( .A(\lte_x_57/B[15] ), .B(n7679), .C(n7681), .D(
        \u_DataPath/u_execute/resAdd1_i [15]), .Z(n8150) );
  HS65_LL_NAND2X4 U5582 ( .A(n9284), .B(n2797), .Z(n8379) );
  HS65_LL_OAI12X3 U5583 ( .A(n2951), .B(n8381), .C(n2950), .Z(n3588) );
  HS65_LH_NAND2X7 U5584 ( .A(n1885), .B(\u_DataPath/toPC2_i [25]), .Z(n8137)
         );
  HS65_LL_OAI12X5 U5585 ( .A(n8439), .B(n3170), .C(n3169), .Z(n5251) );
  HS65_LH_NAND2X7 U5587 ( .A(n1885), .B(n8968), .Z(n8078) );
  HS65_LL_MUX21I1X6 U5588 ( .D0(n8449), .D1(n8730), .S0(n3174), .Z(n4902) );
  HS65_LH_NAND2AX7 U5589 ( .A(n8633), .B(n2797), .Z(n8434) );
  HS65_LH_IVX9 U5591 ( .A(n8821), .Z(n7981) );
  HS65_LH_AOI22X4 U5592 ( .A(\add_x_50/A[23] ), .B(n7679), .C(n7682), .D(
        \u_DataPath/u_execute/resAdd1_i [23]), .Z(n8139) );
  HS65_LH_NOR2X6 U5593 ( .A(n4330), .B(n3338), .Z(n3848) );
  HS65_LH_NOR2X3 U5594 ( .A(n3950), .B(n3338), .Z(n4190) );
  HS65_LH_AND2X4 U5595 ( .A(addr_to_iram_28), .B(n7456), .Z(n7457) );
  HS65_LH_NOR2X6 U5596 ( .A(n8673), .B(n2772), .Z(n8381) );
  HS65_LL_OAI21X2 U5597 ( .A(n8653), .B(n2772), .C(n3114), .Z(n8447) );
  HS65_LHS_XNOR2X3 U5600 ( .A(n8880), .B(n5920), .Z(
        \u_DataPath/u_execute/resAdd1_i [26]) );
  HS65_LH_IVX9 U5601 ( .A(n8152), .Z(\u_DataPath/branch_target_i [14]) );
  HS65_LH_IVX9 U5603 ( .A(n8140), .Z(\u_DataPath/branch_target_i [23]) );
  HS65_LH_AOI22X3 U5605 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][3] ), .B(n9226), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][3] ), .D(n9193), .Z(n6450) );
  HS65_LH_AO22X9 U5607 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][8] ), .B(n9254), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][8] ), .D(
        n9244), .Z(n6855) );
  HS65_LH_AOI22X3 U5610 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][0] ), .B(n9246), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][0] ), .D(n9262), .Z(n6205) );
  HS65_LH_AOI22X3 U5612 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][28] ), .B(n9255), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][28] ), .D(
        n9195), .Z(n6522) );
  HS65_LH_AOI22X3 U5613 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][28] ), .B(n9206), 
        .C(n9205), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][28] ), .Z(n7576)
         );
  HS65_LH_AOI22X3 U5614 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][28] ), .B(n9248), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][28] ), .D(
        n9163), .Z(n6535) );
  HS65_LH_AO22X9 U5615 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][28] ), .B(n9469), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][28] ), .D(
        n9475), .Z(n6525) );
  HS65_LH_AOI22X3 U5620 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][26] ), .B(n9188), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][26] ), .D(
        n9190), .Z(n6937) );
  HS65_LH_AOI22X3 U5622 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][26] ), .B(n9255), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][26] ), .D(
        n9195), .Z(n6933) );
  HS65_LH_AO22X9 U5625 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][3] ), .B(n9187), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][3] ), .D(
        n9194), .Z(n6441) );
  HS65_LH_AOI22X3 U5626 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][3] ), .B(n8851), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][3] ), .D(n9264), .Z(n6446) );
  HS65_LH_AOI22X3 U5628 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][30] ), .B(n9206), 
        .C(n9205), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][30] ), .Z(n7530)
         );
  HS65_LH_AOI22X3 U5629 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][30] ), .B(n9204), 
        .C(n9203), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][30] ), .Z(n7529)
         );
  HS65_LH_AOI22X3 U5630 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][8] ), .B(n8938), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][8] ), .D(n9264), .Z(n6653) );
  HS65_LH_NAND2X7 U5631 ( .A(n1885), .B(\u_DataPath/toPC2_i [23]), .Z(n8140)
         );
  HS65_LHS_XOR2X3 U5632 ( .A(n9001), .B(n5584), .Z(\u_DataPath/toPC2_i [24])
         );
  HS65_LH_BFX18 U5633 ( .A(n8316), .Z(n7697) );
  HS65_LL_AO112X9 U5634 ( .A(n8696), .B(n2712), .C(n3102), .D(n3101), .Z(n3103) );
  HS65_LH_NOR2X6 U5635 ( .A(n8954), .B(n7956), .Z(\u_DataPath/u_idexreg/N15 )
         );
  HS65_LH_NOR2X6 U5636 ( .A(n8750), .B(n7956), .Z(\u_DataPath/u_idexreg/N16 )
         );
  HS65_LH_NAND2X7 U5639 ( .A(n1885), .B(n8966), .Z(n8098) );
  HS65_LL_NOR3X1 U5640 ( .A(n3174), .B(n8429), .C(n8430), .Z(n3143) );
  HS65_LH_NAND2X7 U5641 ( .A(n1885), .B(\u_DataPath/toPC2_i [14]), .Z(n8152)
         );
  HS65_LL_NOR3X1 U5644 ( .A(n3184), .B(n8420), .C(n8421), .Z(n3140) );
  HS65_LL_NOR3X1 U5645 ( .A(n3174), .B(n8432), .C(n8433), .Z(n3175) );
  HS65_LH_NAND2X7 U5646 ( .A(n1885), .B(n9020), .Z(n8081) );
  HS65_LH_AOI22X3 U5650 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][19] ), .B(n9247), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][19] ), .D(
        n9227), .Z(n6769) );
  HS65_LH_AOI22X3 U5653 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][14] ), .B(n9247), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][14] ), .D(
        n9227), .Z(n6088) );
  HS65_LH_AOI22X3 U5655 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][9] ), .B(n9191), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][9] ), .D(
        n9471), .Z(n6990) );
  HS65_LH_AOI22X3 U5656 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][29] ), .B(n9247), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][29] ), .D(
        n9227), .Z(n7554) );
  HS65_LH_AOI22X3 U5658 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][29] ), .B(n9250), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][29] ), .D(
        n9265), .Z(n7553) );
  HS65_LH_AO22X9 U5661 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][20] ), .B(n9206), 
        .C(n9205), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][20] ), .Z(n7097)
         );
  HS65_LH_AOI22X3 U5662 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][19] ), .B(n9250), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][19] ), .D(
        n9265), .Z(n6774) );
  HS65_LH_AOI22X3 U5663 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][20] ), .B(n9246), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][20] ), .D(
        n9067), .Z(n6591) );
  HS65_LH_AOI22X3 U5664 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][19] ), .B(n9248), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][19] ), .D(
        n9240), .Z(n6300) );
  HS65_LH_AO22X4 U5665 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][20] ), .B(n9469), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][20] ), .D(
        n9475), .Z(n6588) );
  HS65_LH_AOI22X3 U5669 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][11] ), .B(n9255), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][11] ), .D(
        n9116), .Z(n6502) );
  HS65_LH_AO22X9 U5670 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][23] ), .B(n9254), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][23] ), .D(
        n9244), .Z(n7130) );
  HS65_LH_AOI22X3 U5674 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][19] ), .B(n9255), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][19] ), .D(
        n9116), .Z(n6289) );
  HS65_LH_AOI22X3 U5675 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][15] ), .B(n9255), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][15] ), .D(
        n9195), .Z(n6884) );
  HS65_LH_AO22X9 U5678 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][21] ), .B(n9254), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][21] ), .D(
        n9244), .Z(n6008) );
  HS65_LH_AOI22X3 U5682 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][10] ), .B(n9247), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][10] ), .D(
        n9227), .Z(n7044) );
  HS65_LH_AO22X9 U5683 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][27] ), .B(n9469), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][27] ), .D(
        n8853), .Z(n6314) );
  HS65_LH_AOI22X3 U5685 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][10] ), .B(n8938), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][10] ), .D(
        n9264), .Z(n6713) );
  HS65_LH_AOI22X3 U5688 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][10] ), .B(n9191), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][10] ), .D(
        n9471), .Z(n6711) );
  HS65_LH_AOI22X3 U5689 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][10] ), .B(n9250), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][10] ), .D(
        n9265), .Z(n7049) );
  HS65_LH_AOI22X3 U5691 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][27] ), .B(n9248), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][27] ), .D(
        n9240), .Z(n6321) );
  HS65_LH_AO22X9 U5695 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][6] ), .B(n9254), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][6] ), .D(
        n9244), .Z(n6835) );
  HS65_LH_AOI22X3 U5697 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][17] ), .B(n9159), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][17] ), .D(
        n9265), .Z(n5965) );
  HS65_LH_AO22X9 U5700 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][17] ), .B(n9254), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][17] ), .D(
        n9244), .Z(n5966) );
  HS65_LH_AO22X9 U5703 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][12] ), .B(n9254), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][12] ), .D(
        n9244), .Z(n7150) );
  HS65_LH_AOI22X3 U5706 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][18] ), .B(n9259), 
        .C(n9256), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][18] ), .Z(n7227)
         );
  HS65_LH_AO22X4 U5707 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][18] ), .B(n9258), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][18] ), .D(
        n9245), .Z(n7222) );
  HS65_LH_AOI22X3 U5712 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][18] ), .B(n9188), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][18] ), .D(
        n9190), .Z(n6670) );
  HS65_LH_AOI22X3 U5713 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][18] ), .B(n9191), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][18] ), .D(
        n9471), .Z(n6671) );
  HS65_LH_AOI22X3 U5714 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][24] ), .B(n9248), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][24] ), .D(
        n9240), .Z(n6279) );
  HS65_LH_AOI22X3 U5715 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][18] ), .B(n9247), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][18] ), .D(
        n9227), .Z(n7226) );
  HS65_LH_AOI22X3 U5717 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][25] ), .B(n9191), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][25] ), .D(
        n9471), .Z(n6959) );
  HS65_LH_AO22X4 U5718 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][31] ), .B(n9258), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][31] ), .D(
        n9245), .Z(n7521) );
  HS65_LH_AOI22X3 U5719 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][25] ), .B(n9255), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][25] ), .D(
        n9195), .Z(n6954) );
  HS65_LH_AOI22X3 U5720 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][24] ), .B(n9255), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][24] ), .D(
        n9116), .Z(n6262) );
  HS65_LH_AOI22X3 U5721 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][6] ), .B(n9191), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][6] ), .D(
        n9471), .Z(n6735) );
  HS65_LH_AOI22X3 U5725 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][6] ), .B(n8938), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][6] ), .D(n9264), .Z(n6737) );
  HS65_LH_AO22X4 U5726 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][24] ), .B(n9258), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][24] ), .D(
        n9245), .Z(n5976) );
  HS65_LH_AOI22X3 U5728 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][9] ), .B(n8938), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][9] ), .D(n9264), .Z(n6995) );
  HS65_LH_AOI22X3 U5729 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][16] ), .B(n9247), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][16] ), .D(
        n9227), .Z(n6068) );
  HS65_LH_AOI22X3 U5732 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][16] ), .B(n9259), 
        .C(n9256), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][16] ), .Z(n6069)
         );
  HS65_LH_AO22X4 U5736 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][16] ), .B(n9258), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][16] ), .D(
        n9245), .Z(n6064) );
  HS65_LH_AO22X9 U5739 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][29] ), .B(n9469), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][29] ), .D(
        n9475), .Z(n6913) );
  HS65_LH_AOI22X3 U5740 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][12] ), .B(n8938), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][12] ), .D(
        n9264), .Z(n6693) );
  HS65_LH_AOI22X3 U5741 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][14] ), .B(n9255), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][14] ), .D(
        n9195), .Z(n6864) );
  HS65_LH_AOI22X3 U5742 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][29] ), .B(n9255), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][29] ), .D(
        n9195), .Z(n6906) );
  HS65_LH_AOI22X3 U5744 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][12] ), .B(n9191), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][12] ), .D(
        n9471), .Z(n6691) );
  HS65_LH_AO22X4 U5745 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][25] ), .B(n9258), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][25] ), .D(
        n9245), .Z(n7480) );
  HS65_LH_AO22X9 U5749 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][13] ), .B(n9258), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][13] ), .D(
        n9245), .Z(n7020) );
  HS65_LH_AOI22X3 U5750 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][29] ), .B(n9204), 
        .C(n9203), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][29] ), .Z(n7549)
         );
  HS65_LH_AOI22X3 U5751 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][9] ), .B(n9188), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][9] ), .D(
        n9190), .Z(n6989) );
  HS65_LH_AOI22X3 U5754 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][29] ), .B(n9206), 
        .C(n9205), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][29] ), .Z(n7550)
         );
  HS65_LH_AO22X9 U5756 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][1] ), .B(n9206), 
        .C(n9205), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][1] ), .Z(n7239)
         );
  HS65_LH_AO22X9 U5758 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][1] ), .B(n9258), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][1] ), .D(
        n9245), .Z(n7242) );
  HS65_LH_AO22X9 U5759 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][1] ), .B(n9204), 
        .C(n9203), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][1] ), .Z(n7238)
         );
  HS65_LH_IVX18 U5760 ( .A(n3239), .Z(n5148) );
  HS65_LHS_XNOR2X3 U5761 ( .A(n8881), .B(n5932), .Z(
        \u_DataPath/u_execute/resAdd1_i [24]) );
  HS65_LH_IVX9 U5762 ( .A(n8173), .Z(\u_DataPath/branch_target_i [9]) );
  HS65_LH_NAND2X7 U5763 ( .A(n4620), .B(n3239), .Z(n4431) );
  HS65_LH_IVX9 U5764 ( .A(n8175), .Z(\u_DataPath/branch_target_i [7]) );
  HS65_LH_BFX18 U5765 ( .A(n8368), .Z(n7717) );
  HS65_LH_IVX9 U5767 ( .A(n8142), .Z(\u_DataPath/branch_target_i [21]) );
  HS65_LH_IVX9 U5768 ( .A(n8149), .Z(\u_DataPath/branch_target_i [16]) );
  HS65_LH_NOR2X6 U5769 ( .A(n2813), .B(n8222), .Z(n8305) );
  HS65_LH_NOR2X6 U5770 ( .A(n8641), .B(n3181), .Z(n2890) );
  HS65_LH_IVX9 U5771 ( .A(n8223), .Z(n8300) );
  HS65_LH_NOR2AX6 U5772 ( .A(n8690), .B(n2794), .Z(n8436) );
  HS65_LH_NOR2X6 U5774 ( .A(n8640), .B(n3181), .Z(n3117) );
  HS65_LH_NAND2X7 U5777 ( .A(n8996), .B(n8023), .Z(n7956) );
  HS65_LH_AO22X4 U5779 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][4] ), .B(n9258), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][4] ), .D(
        n9245), .Z(n6022) );
  HS65_LH_AOI22X3 U5781 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][4] ), .B(n9247), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][4] ), .D(n9227), .Z(n6028) );
  HS65_LH_AOI22X3 U5782 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][7] ), .B(n9250), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][7] ), .D(n9265), .Z(n6053) );
  HS65_LH_AOI22X3 U5783 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][7] ), .B(n9247), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][7] ), .D(n9227), .Z(n6048) );
  HS65_LH_AO22X4 U5784 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][7] ), .B(n9258), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][7] ), .D(
        n9245), .Z(n6044) );
  HS65_LH_AOI22X3 U5785 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][7] ), .B(n9188), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][7] ), .D(
        n9190), .Z(n6464) );
  HS65_LH_AOI22X3 U5786 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][7] ), .B(n9191), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][7] ), .D(
        n9471), .Z(n6465) );
  HS65_LH_NAND2X7 U5791 ( .A(n1885), .B(\u_DataPath/toPC2_i [16]), .Z(n8149)
         );
  HS65_LH_NAND2X7 U5792 ( .A(n1885), .B(n9016), .Z(n8087) );
  HS65_LH_NAND2X7 U5793 ( .A(n1885), .B(\u_DataPath/toPC2_i [7]), .Z(n8175) );
  HS65_LH_NAND2X7 U5794 ( .A(n1885), .B(\u_DataPath/toPC2_i [9]), .Z(n8173) );
  HS65_LH_NAND2X7 U5795 ( .A(n1885), .B(\u_DataPath/toPC2_i [10]), .Z(n8172)
         );
  HS65_LH_NOR2X6 U5796 ( .A(n9111), .B(n8071), .Z(n7950) );
  HS65_LH_IVX9 U5797 ( .A(n7705), .Z(n7703) );
  HS65_LH_NOR2X6 U5798 ( .A(n7455), .B(n7454), .Z(n7387) );
  HS65_LH_NAND2X7 U5800 ( .A(n9438), .B(n8186), .Z(n8222) );
  HS65_LL_NOR3X1 U5801 ( .A(n9045), .B(n9069), .C(n8071), .Z(
        \u_DataPath/cw_to_ex_i [17]) );
  HS65_LL_OAI21X2 U5802 ( .A(\u_DataPath/dataOut_exe_i [4]), .B(n3178), .C(
        n2944), .Z(n2945) );
  HS65_LH_IVX9 U5803 ( .A(n7705), .Z(n7702) );
  HS65_LL_OAI12X3 U5804 ( .A(n9131), .B(n5842), .C(n9033), .Z(n5932) );
  HS65_LH_NAND2X7 U5805 ( .A(n1885), .B(n6861), .Z(n8368) );
  HS65_LH_NOR2X6 U5806 ( .A(n7474), .B(n7473), .Z(n7406) );
  HS65_LH_NAND2X7 U5807 ( .A(n1885), .B(\u_DataPath/toPC2_i [21]), .Z(n8142)
         );
  HS65_LH_NOR2X6 U5811 ( .A(n8739), .B(n8071), .Z(n8513) );
  HS65_LH_IVX9 U5813 ( .A(n7808), .Z(n7812) );
  HS65_LH_IVX9 U5814 ( .A(n5605), .Z(n5587) );
  HS65_LH_IVX9 U5816 ( .A(n7721), .Z(n7725) );
  HS65_LH_NAND2X7 U5817 ( .A(n7386), .B(n7385), .Z(n7454) );
  HS65_LHS_XNOR2X3 U5818 ( .A(n8987), .B(n5924), .Z(
        \u_DataPath/u_execute/resAdd1_i [22]) );
  HS65_LH_NAND2X7 U5819 ( .A(addr_to_iram_18), .B(n7470), .Z(n7471) );
  HS65_LH_IVX9 U5821 ( .A(n7850), .Z(n7854) );
  HS65_LH_NAND2X7 U5822 ( .A(addr_to_iram_20), .B(n7467), .Z(n7468) );
  HS65_LL_NAND2X2 U5823 ( .A(n8157), .B(n2710), .Z(n2964) );
  HS65_LHS_XNOR2X3 U5824 ( .A(n9234), .B(n7305), .Z(
        \u_DataPath/u_execute/link_value_i [22]) );
  HS65_LH_IVX9 U5826 ( .A(n7401), .Z(n8038) );
  HS65_LH_IVX9 U5827 ( .A(n7787), .Z(n7791) );
  HS65_LH_IVX9 U5831 ( .A(n7822), .Z(n7826) );
  HS65_LH_IVX9 U5834 ( .A(n8361), .Z(n7708) );
  HS65_LH_NAND2X5 U5836 ( .A(n3090), .B(n8380), .Z(n2991) );
  HS65_LH_IVX9 U5838 ( .A(n7843), .Z(n7847) );
  HS65_LH_IVX7 U5839 ( .A(n7405), .Z(n7979) );
  HS65_LH_IVX9 U5841 ( .A(n7892), .Z(n7896) );
  HS65_LH_NOR2X6 U5842 ( .A(n7380), .B(n7452), .Z(n7467) );
  HS65_LH_NOR2X6 U5843 ( .A(n7382), .B(n7452), .Z(n7470) );
  HS65_LHS_XOR2X3 U5844 ( .A(n7453), .B(n7452), .Z(\u_DataPath/pc_4_i [18]) );
  HS65_LH_NOR2X6 U5845 ( .A(n7449), .B(n7448), .Z(n7362) );
  HS65_LH_IVX9 U5846 ( .A(n7749), .Z(n7753) );
  HS65_LH_IVX9 U5847 ( .A(n7829), .Z(n7833) );
  HS65_LH_IVX9 U5848 ( .A(n7864), .Z(n7868) );
  HS65_LH_IVX9 U5849 ( .A(n7801), .Z(n7805) );
  HS65_LH_IVX9 U5850 ( .A(n7356), .Z(n7385) );
  HS65_LH_IVX9 U5851 ( .A(n7836), .Z(n7840) );
  HS65_LH_NOR2X6 U5853 ( .A(n7451), .B(n7450), .Z(n7389) );
  HS65_LH_IVX9 U5854 ( .A(n7794), .Z(n7798) );
  HS65_LH_IVX9 U5855 ( .A(n7857), .Z(n7861) );
  HS65_LH_IVX9 U5856 ( .A(n7885), .Z(n7889) );
  HS65_LH_IVX9 U5857 ( .A(n7906), .Z(n7910) );
  HS65_LH_IVX9 U5858 ( .A(n7899), .Z(n7903) );
  HS65_LH_IVX9 U5859 ( .A(n7759), .Z(n7763) );
  HS65_LH_IVX9 U5860 ( .A(n7735), .Z(n7739) );
  HS65_LH_IVX9 U5862 ( .A(n7913), .Z(n7917) );
  HS65_LH_IVX9 U5863 ( .A(n7766), .Z(n7770) );
  HS65_LH_NOR2X6 U5864 ( .A(n7335), .B(n7334), .Z(n7401) );
  HS65_LH_IVX9 U5865 ( .A(n7871), .Z(n7875) );
  HS65_LH_OAI12X3 U5866 ( .A(n8972), .B(n2799), .C(n9130), .Z(n5693) );
  HS65_LH_OAI12X3 U5868 ( .A(n9056), .B(n2799), .C(n5573), .Z(n5605) );
  HS65_LH_IVX9 U5869 ( .A(n7728), .Z(n7732) );
  HS65_LH_OAI12X3 U5870 ( .A(n9392), .B(n2799), .C(n9239), .Z(n5686) );
  HS65_LH_NAND2X7 U5871 ( .A(n1885), .B(\u_DataPath/toPC2_i [4]), .Z(n8178) );
  HS65_LH_OR2X9 U5872 ( .A(n9125), .B(n3980), .Z(n2843) );
  HS65_LH_IVX9 U5873 ( .A(n7742), .Z(n7746) );
  HS65_LH_NAND2X5 U5874 ( .A(n7693), .B(n9138), .Z(n8304) );
  HS65_LH_NAND2X7 U5875 ( .A(addr_to_iram_6), .B(n7464), .Z(n7465) );
  HS65_LL_AND2X9 U5876 ( .A(n4846), .B(n3293), .Z(n3379) );
  HS65_LH_NAND2X7 U5877 ( .A(n7361), .B(n7461), .Z(n7448) );
  HS65_LH_NOR2X6 U5880 ( .A(n6481), .B(n6480), .Z(n6485) );
  HS65_LH_NAND2X7 U5881 ( .A(n7398), .B(n7397), .Z(n8021) );
  HS65_LH_NAND2X7 U5883 ( .A(n7368), .B(n7461), .Z(n7356) );
  HS65_LH_NAND2X7 U5884 ( .A(n8441), .B(n2814), .Z(n8361) );
  HS65_LH_NAND2X7 U5885 ( .A(n7410), .B(n7614), .Z(n7405) );
  HS65_LH_NAND2X7 U5886 ( .A(n1885), .B(\u_DataPath/toPC2_i [3]), .Z(n8179) );
  HS65_LH_NAND2X7 U5888 ( .A(n6757), .B(n7439), .Z(n7631) );
  HS65_LL_OR2X4 U5889 ( .A(n3174), .B(n8384), .Z(n2940) );
  HS65_LH_IVX7 U5890 ( .A(n9144), .Z(n8043) );
  HS65_LL_NAND2X4 U5892 ( .A(n8156), .B(n2800), .Z(n8371) );
  HS65_LH_NAND2X7 U5893 ( .A(n7377), .B(n7376), .Z(n7450) );
  HS65_LHS_XNOR2X6 U5894 ( .A(n7343), .B(n7461), .Z(\u_DataPath/pc_4_i [10])
         );
  HS65_LH_NAND2X7 U5895 ( .A(n8020), .B(n7615), .Z(n7335) );
  HS65_LH_BFX18 U5896 ( .A(n7692), .Z(n7693) );
  HS65_LHS_XOR2X6 U5897 ( .A(n7620), .B(n7619), .Z(
        \u_DataPath/u_execute/link_value_i [5]) );
  HS65_LH_IVX9 U5898 ( .A(n3465), .Z(n4630) );
  HS65_LH_IVX4 U5900 ( .A(n7955), .Z(n7393) );
  HS65_LL_NAND2X4 U5901 ( .A(n2896), .B(n2895), .Z(n2916) );
  HS65_LH_NOR2X6 U5903 ( .A(n7375), .B(n7374), .Z(n7376) );
  HS65_LL_NAND2X4 U5904 ( .A(n2915), .B(n2914), .Z(n2917) );
  HS65_LH_IVX9 U5905 ( .A(n7370), .Z(n7461) );
  HS65_LH_NOR2X6 U5906 ( .A(n7370), .B(n7369), .Z(n7377) );
  HS65_LH_NOR2X6 U5907 ( .A(n7354), .B(n7353), .Z(n8047) );
  HS65_LL_NOR2X5 U5908 ( .A(n5959), .B(n5957), .Z(n6129) );
  HS65_LH_NAND3X3 U5909 ( .A(opcode_i[2]), .B(n7400), .C(n7403), .Z(n7614) );
  HS65_LH_NAND2X7 U5910 ( .A(n6490), .B(n6489), .Z(n6494) );
  HS65_LH_NAND2X7 U5911 ( .A(opcode_i[1]), .B(n7332), .Z(n7615) );
  HS65_LH_NAND2X4 U5913 ( .A(opcode_i[1]), .B(n7403), .Z(n7967) );
  HS65_LH_AOI21X6 U5914 ( .A(n3148), .B(\u_DataPath/from_mem_data_out_i [28]), 
        .C(n3115), .Z(n7653) );
  HS65_LL_NOR2X5 U5915 ( .A(n5959), .B(n5951), .Z(n6112) );
  HS65_LL_NOR2X5 U5917 ( .A(n6182), .B(n6185), .Z(n6272) );
  HS65_LH_BFX18 U5918 ( .A(n8180), .Z(n7680) );
  HS65_LH_NAND2X7 U5922 ( .A(n2812), .B(n6163), .Z(n6164) );
  HS65_LL_NAND2X5 U5927 ( .A(\u_DataPath/reg_write_i ), .B(n2892), .Z(n8041)
         );
  HS65_LL_NOR2X5 U5928 ( .A(n5959), .B(n5950), .Z(n6114) );
  HS65_LL_NOR2X5 U5929 ( .A(n5958), .B(n5960), .Z(n6130) );
  HS65_LL_IVX7 U5930 ( .A(n3529), .Z(n7309) );
  HS65_LH_NOR2AX3 U5931 ( .A(\u_DataPath/from_alu_data_out_i [26]), .B(n3148), 
        .Z(n3108) );
  HS65_LH_NAND2X7 U5932 ( .A(n7411), .B(n7392), .Z(n7955) );
  HS65_LH_NAND2X7 U5933 ( .A(n7368), .B(n7367), .Z(n7369) );
  HS65_LH_NOR2X6 U5934 ( .A(n3302), .B(n5161), .Z(n3465) );
  HS65_LL_NOR2X5 U5935 ( .A(n5959), .B(n5960), .Z(n6121) );
  HS65_LH_NAND2X7 U5936 ( .A(n8017), .B(n5938), .Z(n5937) );
  HS65_LH_NAND2X7 U5937 ( .A(n8801), .B(n9346), .Z(n7973) );
  HS65_LH_NAND2X7 U5938 ( .A(\u_DataPath/jaddr_i [20]), .B(n5938), .Z(n5939)
         );
  HS65_LH_NAND2X7 U5939 ( .A(n7408), .B(n7404), .Z(n7613) );
  HS65_LH_NAND2X7 U5940 ( .A(n7342), .B(n7341), .Z(n7370) );
  HS65_LH_IVX9 U5942 ( .A(n7936), .Z(n7944) );
  HS65_LH_CNIVX3 U5943 ( .A(n8122), .Z(\u_DataPath/pc_4_to_ex_i [2]) );
  HS65_LH_CNIVX3 U5944 ( .A(n8119), .Z(\u_DataPath/pc_4_to_ex_i [4]) );
  HS65_LH_CNIVX3 U5945 ( .A(n8126), .Z(\u_DataPath/u_execute/link_value_i [0])
         );
  HS65_LH_CNIVX3 U5946 ( .A(n8365), .Z(\u_DataPath/cw_memwb_i [2]) );
  HS65_LH_CNIVX3 U5947 ( .A(n8034), .Z(\u_DataPath/cw_tomem_i [7]) );
  HS65_LH_IVX9 U5948 ( .A(n8127), .Z(n8180) );
  HS65_LL_NAND2X7 U5951 ( .A(n2871), .B(n7649), .Z(n8029) );
  HS65_LH_NOR2X5 U5952 ( .A(n5707), .B(n5712), .Z(n5534) );
  HS65_LL_NAND2X7 U5954 ( .A(n2871), .B(n7673), .Z(n6488) );
  HS65_LL_IVX7 U5955 ( .A(n3528), .Z(n3529) );
  HS65_LL_NAND2X7 U5956 ( .A(n2871), .B(n7648), .Z(n8028) );
  HS65_LH_NAND2X4 U5957 ( .A(n5698), .B(n5645), .Z(n5649) );
  HS65_LH_NAND2X7 U5958 ( .A(n5540), .B(n5593), .Z(n5574) );
  HS65_LH_NAND2X5 U5959 ( .A(n5536), .B(n5648), .Z(n5538) );
  HS65_LH_IVX9 U5960 ( .A(n7400), .Z(n7392) );
  HS65_LH_NOR2X6 U5961 ( .A(n9422), .B(rst), .Z(n8465) );
  HS65_LH_NAND2X7 U5962 ( .A(n6755), .B(n7423), .Z(n6756) );
  HS65_LH_NOR2X6 U5963 ( .A(n7415), .B(n6750), .Z(n7417) );
  HS65_LH_NOR2X6 U5964 ( .A(\u_DataPath/immediate_ext_dec_i [0]), .B(n8031), 
        .Z(n7954) );
  HS65_LH_NAND2X7 U5965 ( .A(n5749), .B(n5795), .Z(n5826) );
  HS65_LH_NAND2X7 U5966 ( .A(n5741), .B(n5801), .Z(n5777) );
  HS65_LH_NAND3X3 U5967 ( .A(opcode_i[3]), .B(n7408), .C(n8019), .Z(n7957) );
  HS65_LH_NOR2X5 U5969 ( .A(n5910), .B(n5915), .Z(n5735) );
  HS65_LH_IVX4 U5970 ( .A(n5801), .Z(n5804) );
  HS65_LH_NAND2X4 U5971 ( .A(n5772), .B(n5771), .Z(n5783) );
  HS65_LH_NOR2X3 U5972 ( .A(n9465), .B(rst), .Z(\u_DataPath/idex_rt_i [2]) );
  HS65_LL_NAND2X7 U5973 ( .A(n6479), .B(n2815), .Z(n6184) );
  HS65_LH_NOR2X6 U5974 ( .A(\u_DataPath/jaddr_i [20]), .B(n2804), .Z(n5949) );
  HS65_LH_NOR2X6 U5976 ( .A(n7364), .B(n7382), .Z(n7379) );
  HS65_LH_NOR2X3 U5977 ( .A(opcode_i[5]), .B(n7391), .Z(n7404) );
  HS65_LH_NAND2AX4 U5978 ( .A(n7714), .B(n9349), .Z(n7650) );
  HS65_LH_NAND2AX4 U5979 ( .A(n7715), .B(n9176), .Z(n7932) );
  HS65_LH_IVX9 U5980 ( .A(\u_DataPath/immediate_ext_dec_i [3]), .Z(n8031) );
  HS65_LH_IVX9 U5981 ( .A(addr_to_iram_16), .Z(n7453) );
  HS65_LH_NOR2X6 U5982 ( .A(n5890), .B(n5895), .Z(n5801) );
  HS65_LH_IVX9 U5983 ( .A(n5720), .Z(n5554) );
  HS65_LH_NOR2X6 U5985 ( .A(n5874), .B(n5879), .Z(n5749) );
  HS65_LH_CNIVX3 U5986 ( .A(n5562), .Z(n5563) );
  HS65_LH_NAND2X7 U5987 ( .A(opcode_i[0]), .B(opcode_i[2]), .Z(n7964) );
  HS65_LH_IVX9 U5988 ( .A(n5728), .Z(n5553) );
  HS65_LH_BFX18 U5989 ( .A(n8181), .Z(n7682) );
  HS65_LL_NAND2X7 U5990 ( .A(n8441), .B(n8758), .Z(n8310) );
  HS65_LH_NAND2X7 U5991 ( .A(addr_to_iram_6), .B(addr_to_iram_7), .Z(n7340) );
  HS65_LH_IVX9 U5992 ( .A(n5818), .Z(n5750) );
  HS65_LH_NOR2X6 U5993 ( .A(n7196), .B(
        \u_DataPath/u_decode_unit/hdu_0/current_state [1]), .Z(n7215) );
  HS65_LH_IVX9 U5994 ( .A(n5923), .Z(n5753) );
  HS65_LH_IVX9 U5995 ( .A(n5724), .Z(n5552) );
  HS65_LH_NOR2X6 U5996 ( .A(n7442), .B(n7440), .Z(n6757) );
  HS65_LH_NAND2X7 U5997 ( .A(addr_to_iram_0), .B(addr_to_iram_1), .Z(n7337) );
  HS65_LL_AND2X4 U5998 ( .A(n2876), .B(n2875), .Z(n2877) );
  HS65_LH_NAND2X7 U5999 ( .A(\u_DataPath/pc_4_to_ex_i [2]), .B(
        \u_DataPath/pc_4_to_ex_i [3]), .Z(n7415) );
  HS65_LH_NOR2X6 U6000 ( .A(n5808), .B(n5789), .Z(n5774) );
  HS65_LH_NOR2X6 U6001 ( .A(n6753), .B(n7421), .Z(n6755) );
  HS65_LH_NOR2X6 U6002 ( .A(n5797), .B(n5800), .Z(n5741) );
  HS65_LH_NOR2X6 U6003 ( .A(n6754), .B(n7431), .Z(n7423) );
  HS65_LL_NOR2X3 U6004 ( .A(n7013), .B(n7216), .Z(n7310) );
  HS65_LH_NAND2X7 U6005 ( .A(addr_to_iram_2), .B(addr_to_iram_3), .Z(n7336) );
  HS65_LL_IVX9 U6006 ( .A(n2865), .Z(n2871) );
  HS65_LH_NOR2X6 U6007 ( .A(n5770), .B(n5773), .Z(n5743) );
  HS65_LH_NAND2X7 U6008 ( .A(n5666), .B(n5665), .Z(n5671) );
  HS65_LH_IVX9 U6009 ( .A(addr_to_iram_14), .Z(n7455) );
  HS65_LH_NOR2X2 U6010 ( .A(n9230), .B(rst), .Z(\u_DataPath/u_memwbreg/N73 )
         );
  HS65_LH_NAND2X7 U6011 ( .A(addr_to_iram_4), .B(addr_to_iram_5), .Z(n7344) );
  HS65_LH_IVX9 U6012 ( .A(n5673), .Z(n5555) );
  HS65_LH_IVX4 U6013 ( .A(opcode_i[1]), .Z(n7408) );
  HS65_LH_NOR2X6 U6014 ( .A(opcode_i[0]), .B(opcode_i[2]), .Z(n8019) );
  HS65_LH_IVX9 U6015 ( .A(opcode_i[5]), .Z(n7965) );
  HS65_LH_NOR2X6 U6016 ( .A(n5567), .B(n5570), .Z(n5542) );
  HS65_LH_NOR2X6 U6017 ( .A(n5688), .B(n5692), .Z(n5593) );
  HS65_LH_IVX4 U6018 ( .A(n5653), .Z(n5703) );
  HS65_LH_CNIVX3 U6019 ( .A(n5567), .Z(n5568) );
  HS65_LH_NAND2X7 U6020 ( .A(addr_to_iram_12), .B(addr_to_iram_13), .Z(n7384)
         );
  HS65_LH_IVX9 U6021 ( .A(opcode_i[2]), .Z(n7411) );
  HS65_LH_NAND2X7 U6022 ( .A(addr_to_iram_14), .B(addr_to_iram_15), .Z(n7366)
         );
  HS65_LH_NAND2X7 U6023 ( .A(opcode_i[1]), .B(opcode_i[0]), .Z(n7400) );
  HS65_LH_NAND2X7 U6024 ( .A(addr_to_iram_17), .B(addr_to_iram_16), .Z(n7382)
         );
  HS65_LH_NOR2X6 U6025 ( .A(n5600), .B(n5586), .Z(n5571) );
  HS65_LH_NAND2X4 U6026 ( .A(n5818), .B(n5817), .Z(n5822) );
  HS65_LH_NOR2X6 U6027 ( .A(n5589), .B(n5592), .Z(n5540) );
  HS65_LH_CNIVX3 U6028 ( .A(n5874), .Z(n5875) );
  HS65_LH_NAND2X7 U6029 ( .A(addr_to_iram_8), .B(addr_to_iram_9), .Z(n7360) );
  HS65_LH_IVX9 U6030 ( .A(n5927), .Z(n5756) );
  HS65_LH_IVX9 U6031 ( .A(addr_to_iram_25), .Z(n7474) );
  HS65_LH_IVX9 U6032 ( .A(n5610), .Z(n5548) );
  HS65_LH_IVX9 U6033 ( .A(addr_to_iram_27), .Z(n7606) );
  HS65_LH_IVX9 U6034 ( .A(addr_to_iram_23), .Z(n7451) );
  HS65_LH_IVX9 U6035 ( .A(addr_to_iram_10), .Z(n7449) );
  HS65_LH_IVX9 U6036 ( .A(n5919), .Z(n5755) );
  HS65_LH_NAND2X7 U6037 ( .A(addr_to_iram_19), .B(addr_to_iram_18), .Z(n7364)
         );
  HS65_LH_IVX9 U6038 ( .A(n5716), .Z(n5551) );
  HS65_LH_NAND2X7 U6039 ( .A(n2803), .B(n8035), .Z(n7210) );
  HS65_LH_IVX9 U6040 ( .A(addr_to_iram_22), .Z(n7375) );
  HS65_LH_NOR2X6 U6041 ( .A(n5695), .B(n5700), .Z(n5536) );
  HS65_LH_IVX9 U6042 ( .A(n5931), .Z(n5754) );
  HS65_LH_IVX9 U6043 ( .A(n5624), .Z(n5547) );
  HS65_LH_NAND2X7 U6044 ( .A(addr_to_iram_10), .B(addr_to_iram_11), .Z(n7355)
         );
  HS65_LH_CNIVX3 U6045 ( .A(n5638), .Z(n5639) );
  HS65_LH_IVX9 U6046 ( .A(addr_to_iram_20), .Z(n7381) );
  HS65_LH_NOR2X6 U6047 ( .A(\u_DataPath/jaddr_i [24]), .B(n2811), .Z(n6169) );
  HS65_LH_IVX9 U6048 ( .A(addr_to_iram_12), .Z(n7357) );
  HS65_LH_NAND2X7 U6050 ( .A(n8526), .B(\u_DataPath/pc_4_to_ex_i [28]), .Z(
        n5559) );
  HS65_LH_IVX9 U6051 ( .A(\u_DataPath/pc_4_to_ex_i [21]), .Z(n7632) );
  HS65_LH_NAND2X7 U6052 ( .A(\u_DataPath/pc_4_to_ex_i [5]), .B(
        \u_DataPath/pc_4_to_ex_i [4]), .Z(n6750) );
  HS65_LH_IVX7 U6053 ( .A(\u_DataPath/data_read_ex_2_i [6]), .Z(n2926) );
  HS65_LH_IVX9 U6054 ( .A(\u_DataPath/pc_4_to_ex_i [27]), .Z(n7634) );
  HS65_LH_IVX9 U6055 ( .A(\u_DataPath/pc_4_to_ex_i [23]), .Z(n7628) );
  HS65_LH_NAND2X7 U6056 ( .A(n8526), .B(\u_DataPath/pc_4_to_ex_i [29]), .Z(
        n5673) );
  HS65_LH_IVX7 U6057 ( .A(\u_DataPath/data_read_ex_2_i [8]), .Z(n3026) );
  HS65_LH_NAND2X7 U6058 ( .A(n8512), .B(\u_DataPath/pc_4_to_ex_i [15]), .Z(
        n5772) );
  HS65_LH_IVX9 U6059 ( .A(\u_DataPath/pc_4_to_ex_i [20]), .Z(n7442) );
  HS65_LH_IVX7 U6060 ( .A(\u_DataPath/from_alu_data_out_i [4]), .Z(n2942) );
  HS65_LH_NOR2X3 U6061 ( .A(n8467), .B(\u_DataPath/pc_4_to_ex_i [4]), .Z(n5653) );
  HS65_LH_IVX9 U6062 ( .A(n7932), .Z(n2865) );
  HS65_LH_IVX9 U6063 ( .A(n7652), .Z(n6748) );
  HS65_LH_CNIVX3 U6064 ( .A(\u_DataPath/data_read_ex_1_i [26]), .Z(n3112) );
  HS65_LH_IVX9 U6065 ( .A(\u_DataPath/cw_to_ex_i [3]), .Z(n3283) );
  HS65_LH_OR2X9 U6067 ( .A(\u_DataPath/rs_ex_i [1]), .B(
        \u_DataPath/pc_4_to_ex_i [22]), .Z(n5922) );
  HS65_LH_NAND2X7 U6068 ( .A(n8525), .B(\u_DataPath/pc_4_to_ex_i [9]), .Z(
        n5892) );
  HS65_LH_OR2X9 U6069 ( .A(\u_DataPath/rs_ex_i [3]), .B(
        \u_DataPath/pc_4_to_ex_i [24]), .Z(n5930) );
  HS65_LH_NAND2X7 U6070 ( .A(n8526), .B(\u_DataPath/pc_4_to_ex_i [30]), .Z(
        n5667) );
  HS65_LH_IVX7 U6071 ( .A(\u_DataPath/data_read_ex_2_i [11]), .Z(n3010) );
  HS65_LH_NAND2X7 U6072 ( .A(\u_DataPath/rs_ex_i [2]), .B(
        \u_DataPath/pc_4_to_ex_i [23]), .Z(n5841) );
  HS65_LH_IVX9 U6073 ( .A(\u_DataPath/cw_tomem_i [7]), .Z(n3435) );
  HS65_LH_IVX9 U6074 ( .A(\u_DataPath/cw_tomem_i [3]), .Z(n8162) );
  HS65_LH_NAND2X7 U6075 ( .A(n8526), .B(\u_DataPath/pc_4_to_ex_i [22]), .Z(
        n5640) );
  HS65_LH_IVX9 U6076 ( .A(\u_DataPath/rs_ex_i [2]), .Z(n2868) );
  HS65_LH_NAND2X7 U6077 ( .A(n8510), .B(\u_DataPath/pc_4_to_ex_i [13]), .Z(
        n5602) );
  HS65_LH_NAND2X7 U6078 ( .A(\u_DataPath/rs_ex_i [3]), .B(
        \u_DataPath/pc_4_to_ex_i [24]), .Z(n5931) );
  HS65_LH_NAND2X7 U6079 ( .A(n8515), .B(\u_DataPath/pc_4_to_ex_i [25]), .Z(
        n5786) );
  HS65_LH_NAND2X7 U6080 ( .A(n8515), .B(\u_DataPath/pc_4_to_ex_i [26]), .Z(
        n5919) );
  HS65_LH_NAND2X7 U6081 ( .A(n8526), .B(\u_DataPath/pc_4_to_ex_i [21]), .Z(
        n5716) );
  HS65_LH_IVX9 U6082 ( .A(\u_DataPath/u_idexreg/N13 ), .Z(n8035) );
  HS65_LH_OR2X9 U6083 ( .A(n8526), .B(\u_DataPath/pc_4_to_ex_i [21]), .Z(n5715) );
  HS65_LH_IVX4 U6084 ( .A(n8515), .Z(n2867) );
  HS65_LH_IVX9 U6085 ( .A(\u_DataPath/data_read_ex_2_i [3]), .Z(n2986) );
  HS65_LH_NAND2X7 U6086 ( .A(n8515), .B(\u_DataPath/pc_4_to_ex_i [27]), .Z(
        n5767) );
  HS65_LH_IVX9 U6087 ( .A(\u_DataPath/rs_ex_i [1]), .Z(n2864) );
  HS65_LH_NAND2X7 U6088 ( .A(n8515), .B(\u_DataPath/pc_4_to_ex_i [28]), .Z(
        n5927) );
  HS65_LH_NAND2X7 U6089 ( .A(n8515), .B(\u_DataPath/pc_4_to_ex_i [29]), .Z(
        n5762) );
  HS65_LH_NAND2X7 U6090 ( .A(n8526), .B(\u_DataPath/pc_4_to_ex_i [20]), .Z(
        n5610) );
  HS65_LH_NAND2X7 U6091 ( .A(n8474), .B(\u_DataPath/pc_4_to_ex_i [7]), .Z(
        n5900) );
  HS65_LH_NAND2X7 U6092 ( .A(n8504), .B(\u_DataPath/pc_4_to_ex_i [14]), .Z(
        n5677) );
  HS65_LH_NAND2X7 U6093 ( .A(n8515), .B(\u_DataPath/pc_4_to_ex_i [30]), .Z(
        n5867) );
  HS65_LH_IVX7 U6094 ( .A(\u_DataPath/data_read_ex_2_i [13]), .Z(n3066) );
  HS65_LH_NAND2X7 U6095 ( .A(n8526), .B(\u_DataPath/pc_4_to_ex_i [19]), .Z(
        n5631) );
  HS65_LH_IVX7 U6096 ( .A(\u_DataPath/from_mem_data_out_i [7]), .Z(n2927) );
  HS65_LH_NAND2X7 U6097 ( .A(n8512), .B(\u_DataPath/pc_4_to_ex_i [15]), .Z(
        n5569) );
  HS65_LH_IVX9 U6098 ( .A(\u_DataPath/cw_to_ex_i [0]), .Z(n5062) );
  HS65_LH_NAND2X7 U6099 ( .A(n8526), .B(\u_DataPath/pc_4_to_ex_i [18]), .Z(
        n5624) );
  HS65_LH_NOR2X3 U6100 ( .A(\u_DataPath/cw_to_ex_i [2]), .B(
        \u_DataPath/cw_to_ex_i [1]), .Z(n3284) );
  HS65_LH_NAND2X7 U6101 ( .A(n8526), .B(\u_DataPath/pc_4_to_ex_i [16]), .Z(
        n5681) );
  HS65_LH_NAND2X7 U6102 ( .A(n8526), .B(\u_DataPath/pc_4_to_ex_i [17]), .Z(
        n5618) );
  HS65_LL_NOR2X2 U6103 ( .A(n8526), .B(\u_DataPath/pc_4_to_ex_i [17]), .Z(
        n5616) );
  HS65_LH_NAND2X7 U6104 ( .A(n8469), .B(\u_DataPath/pc_4_to_ex_i [10]), .Z(
        n5685) );
  HS65_LH_NOR2X6 U6105 ( .A(n9446), .B(rst), .Z(n8181) );
  HS65_LH_NAND2X7 U6106 ( .A(n8526), .B(\u_DataPath/pc_4_to_ex_i [25]), .Z(
        n5728) );
  HS65_LH_NAND2X7 U6107 ( .A(n8526), .B(\u_DataPath/pc_4_to_ex_i [26]), .Z(
        n5564) );
  HS65_LH_NAND2X7 U6108 ( .A(\u_DataPath/pc_4_to_ex_i [7]), .B(
        \u_DataPath/pc_4_to_ex_i [6]), .Z(n7435) );
  HS65_LH_NAND2X7 U6109 ( .A(n8506), .B(\u_DataPath/pc_4_to_ex_i [11]), .Z(
        n5591) );
  HS65_LH_IVX7 U6110 ( .A(\u_DataPath/data_read_ex_1_i [7]), .Z(n2930) );
  HS65_LH_NAND2X7 U6111 ( .A(n8526), .B(\u_DataPath/pc_4_to_ex_i [24]), .Z(
        n5583) );
  HS65_LH_NAND2X7 U6112 ( .A(\u_DataPath/idex_rt_i [4]), .B(
        \u_DataPath/pc_4_to_ex_i [20]), .Z(n5825) );
  HS65_LH_NAND2X7 U6113 ( .A(n8526), .B(\u_DataPath/pc_4_to_ex_i [27]), .Z(
        n5720) );
  HS65_LH_NAND2X7 U6115 ( .A(\u_DataPath/rs_ex_i [1]), .B(
        \u_DataPath/pc_4_to_ex_i [22]), .Z(n5923) );
  HS65_LH_NAND2X7 U6116 ( .A(n8508), .B(\u_DataPath/pc_4_to_ex_i [12]), .Z(
        n5603) );
  HS65_LH_NAND2X7 U6117 ( .A(n8526), .B(\u_DataPath/pc_4_to_ex_i [23]), .Z(
        n5724) );
  HS65_LH_IVX9 U6118 ( .A(Data_out_fromRAM[7]), .Z(n8224) );
  HS65_LH_IVX9 U6119 ( .A(Data_out_fromRAM[23]), .Z(n8220) );
  HS65_LL_NOR4X4 U6121 ( .A(n5179), .B(n5178), .C(n8326), .D(n8327), .Z(n5180)
         );
  HS65_LL_NAND3X2 U6122 ( .A(n8328), .B(n8329), .C(n8330), .Z(n5178) );
  HS65_LL_NOR2X2 U6124 ( .A(n8323), .B(n8322), .Z(n5177) );
  HS65_LL_NAND3X2 U6126 ( .A(n8336), .B(n8335), .C(n8334), .Z(n5182) );
  HS65_LL_CBI4I1X3 U6127 ( .A(n8780), .B(n9329), .C(n9044), .D(n8598), .Z(
        \u_DataPath/dataOut_exe_i [19]) );
  HS65_LL_NOR3X2 U6129 ( .A(n3755), .B(n3754), .C(n3753), .Z(n3774) );
  HS65_LH_OAI12X3 U6130 ( .A(n8310), .B(n8350), .C(n8233), .Z(
        \u_DataPath/dataOut_exe_i [10]) );
  HS65_LH_OAI12X3 U6131 ( .A(n8310), .B(n8342), .C(n8286), .Z(
        \u_DataPath/dataOut_exe_i [2]) );
  HS65_LL_NAND3X2 U6132 ( .A(n4422), .B(n4421), .C(n4420), .Z(n4423) );
  HS65_LL_NAND3AX3 U6135 ( .A(n2851), .B(n3307), .C(n3306), .Z(n3308) );
  HS65_LL_AOI21X3 U6136 ( .A(n7327), .B(n4764), .C(n4763), .Z(n8336) );
  HS65_LL_NAND4ABX3 U6138 ( .A(n3369), .B(n3368), .C(n3367), .D(n3366), .Z(
        n3370) );
  HS65_LL_NAND2AX4 U6141 ( .A(n4099), .B(n4098), .Z(n8348) );
  HS65_LL_NAND2AX4 U6142 ( .A(n3819), .B(n3818), .Z(n8338) );
  HS65_LL_NAND2X2 U6143 ( .A(n5492), .B(n4140), .Z(n4141) );
  HS65_LL_NAND4ABX3 U6144 ( .A(n4455), .B(n4454), .C(n4453), .D(n4452), .Z(
        n4456) );
  HS65_LL_NAND2AX4 U6147 ( .A(n3657), .B(n3656), .Z(n3658) );
  HS65_LL_NAND2AX4 U6149 ( .A(n5476), .B(n5475), .Z(n5477) );
  HS65_LL_NOR2AX3 U6153 ( .A(n4076), .B(n4075), .Z(n4089) );
  HS65_LL_NAND4ABX3 U6156 ( .A(n4855), .B(n4854), .C(n4853), .D(n4852), .Z(
        n4856) );
  HS65_LLS_XNOR2X3 U6157 ( .A(n3638), .B(n3637), .Z(n3639) );
  HS65_LHS_XNOR2X6 U6158 ( .A(n3457), .B(n3456), .Z(n3505) );
  HS65_LLS_XNOR2X3 U6159 ( .A(n4373), .B(n4372), .Z(n4397) );
  HS65_LL_NOR2AX3 U6160 ( .A(n3602), .B(n3601), .Z(n3603) );
  HS65_LLS_XNOR2X3 U6161 ( .A(n2858), .B(n3619), .Z(n3620) );
  HS65_LL_NAND2X2 U6166 ( .A(n4074), .B(n4073), .Z(n4075) );
  HS65_LL_AND2X4 U6168 ( .A(n4774), .B(n3652), .Z(n2861) );
  HS65_LLS_XNOR2X3 U6171 ( .A(n4600), .B(n4599), .Z(n4635) );
  HS65_LL_NOR2AX3 U6172 ( .A(n4233), .B(n4232), .Z(n4234) );
  HS65_LL_NAND3X2 U6173 ( .A(n3412), .B(n3411), .C(n3410), .Z(n3413) );
  HS65_LL_NOR3X1 U6174 ( .A(n4037), .B(n4036), .C(n4035), .Z(n4054) );
  HS65_LHS_XNOR2X6 U6175 ( .A(n3909), .B(n3908), .Z(n3936) );
  HS65_LL_NOR2AX3 U6177 ( .A(n3701), .B(n3700), .Z(n3702) );
  HS65_LLS_XNOR2X3 U6180 ( .A(n4026), .B(n4025), .Z(n4056) );
  HS65_LL_OAI12X3 U6182 ( .A(n4427), .B(n4714), .C(n4426), .Z(n4428) );
  HS65_LL_NAND4ABX3 U6187 ( .A(n4359), .B(n4358), .C(n4357), .D(n4356), .Z(
        n8344) );
  HS65_LL_OR2X4 U6188 ( .A(n4485), .B(n4484), .Z(n4497) );
  HS65_LL_NOR2AX3 U6189 ( .A(n3618), .B(n3617), .Z(n3619) );
  HS65_LLS_XNOR2X3 U6191 ( .A(n4179), .B(n4178), .Z(n4180) );
  HS65_LH_OAI21X3 U6192 ( .A(n4942), .B(n4630), .C(n3810), .Z(n3811) );
  HS65_LL_NAND3AX3 U6193 ( .A(n3474), .B(n3473), .C(n3472), .Z(n3480) );
  HS65_LL_NAND3X2 U6194 ( .A(n4835), .B(n4834), .C(n4833), .Z(n4855) );
  HS65_LH_NAND3X5 U6195 ( .A(n4134), .B(n4133), .C(n4132), .Z(n4135) );
  HS65_LH_NAND2X4 U6196 ( .A(n5486), .B(n4391), .Z(n4228) );
  HS65_LL_NOR4ABX2 U6197 ( .A(n4628), .B(n4627), .C(n4626), .D(n4625), .Z(
        n4629) );
  HS65_LH_OAI21X3 U6198 ( .A(n4954), .B(n4630), .C(n3722), .Z(n3754) );
  HS65_LH_NOR3X4 U6199 ( .A(n3395), .B(n3394), .C(n3393), .Z(n3415) );
  HS65_LL_OAI112X1 U6205 ( .A(n3988), .B(n2848), .C(n3989), .D(n3987), .Z(
        n4022) );
  HS65_LL_OAI211X1 U6206 ( .A(n4951), .B(n4630), .C(n3550), .D(n3549), .Z(
        n3551) );
  HS65_LH_OAI21X3 U6208 ( .A(n5499), .B(n4289), .C(n4157), .Z(n4158) );
  HS65_LL_NAND3X2 U6209 ( .A(n4390), .B(n4389), .C(n4388), .Z(n4394) );
  HS65_LL_NAND3X2 U6210 ( .A(n3934), .B(n3933), .C(n3932), .Z(n3935) );
  HS65_LL_OAI21X2 U6211 ( .A(n4476), .B(n4440), .C(n4439), .Z(n4454) );
  HS65_LL_NOR2AX3 U6213 ( .A(n4941), .B(n4940), .Z(n5176) );
  HS65_LH_OAI211X3 U6215 ( .A(n4753), .B(n3320), .C(n4752), .D(n4751), .Z(
        n4754) );
  HS65_LL_OAI12X2 U6222 ( .A(n5432), .B(n5431), .C(n5430), .Z(n5442) );
  HS65_LH_AOI21X2 U6225 ( .A(n4712), .B(n4711), .C(n4710), .Z(n4713) );
  HS65_LL_NOR3X1 U6229 ( .A(n3352), .B(n3351), .C(n3350), .Z(n3367) );
  HS65_LL_AOI22X1 U6230 ( .A(n4667), .B(n3331), .C(n4836), .D(n3696), .Z(n3332) );
  HS65_LH_NAND2X5 U6231 ( .A(n5492), .B(n4345), .Z(n4357) );
  HS65_LH_NAND2X4 U6233 ( .A(n4038), .B(n5484), .Z(n3745) );
  HS65_LL_IVX2 U6234 ( .A(n4405), .Z(n4502) );
  HS65_LL_AOI22X1 U6235 ( .A(n5510), .B(n4567), .C(n4667), .D(n3835), .Z(n3654) );
  HS65_LH_NAND2AX4 U6236 ( .A(n3615), .B(n3666), .Z(n3616) );
  HS65_LL_NAND3X2 U6237 ( .A(n4002), .B(n4001), .C(n4000), .Z(n4016) );
  HS65_LH_AOI21X2 U6238 ( .A(n5517), .B(n5163), .C(n4656), .Z(n4670) );
  HS65_LL_NAND4ABX3 U6239 ( .A(n5166), .B(n4995), .C(n5165), .D(n5169), .Z(
        n4996) );
  HS65_LL_NAND2X2 U6242 ( .A(n4667), .B(n4480), .Z(n3411) );
  HS65_LH_AOI12X2 U6244 ( .A(n4536), .B(n4535), .C(n4534), .Z(n4537) );
  HS65_LH_AOI21X2 U6245 ( .A(n4461), .B(n4711), .C(n5290), .Z(n4462) );
  HS65_LL_NOR2AX3 U6250 ( .A(n5322), .B(n5321), .Z(n5323) );
  HS65_LH_OAI22X3 U6251 ( .A(n4630), .B(n4983), .C(n4738), .D(n4574), .Z(n4575) );
  HS65_LH_IVX9 U6252 ( .A(n8130), .Z(\u_DataPath/branch_target_i [31]) );
  HS65_LL_AOI21X2 U6255 ( .A(n5275), .B(n5274), .C(n5273), .Z(n5276) );
  HS65_LH_OAI211X3 U6256 ( .A(n4846), .B(n4622), .C(n4621), .D(n4748), .Z(
        n4626) );
  HS65_LHS_XNOR2X6 U6261 ( .A(n4264), .B(n4263), .Z(n4265) );
  HS65_LLS_XOR2X3 U6262 ( .A(n3770), .B(n3769), .Z(n3771) );
  HS65_LH_NOR2AX3 U6265 ( .A(n4400), .B(n3206), .Z(n3208) );
  HS65_LH_OAI21X3 U6267 ( .A(n2787), .B(n4846), .C(n4844), .Z(n3721) );
  HS65_LL_AOI21X2 U6268 ( .A(n4294), .B(n5483), .C(n3866), .Z(n3867) );
  HS65_LH_OAI211X3 U6269 ( .A(n2998), .B(n4846), .C(n4845), .D(n4844), .Z(
        n4847) );
  HS65_LL_OAI22X1 U6270 ( .A(n3320), .B(n4564), .C(n4659), .D(n4746), .Z(n3547) );
  HS65_LL_OAI12X2 U6273 ( .A(n4305), .B(n9540), .C(n4220), .Z(n4230) );
  HS65_LL_AOI21X2 U6274 ( .A(n4673), .B(n4828), .C(n4226), .Z(n4227) );
  HS65_LH_OAI21X3 U6275 ( .A(n3718), .B(n4070), .C(n3717), .Z(n3755) );
  HS65_LH_OAI21X3 U6279 ( .A(n4662), .B(n4440), .C(n3626), .Z(n3632) );
  HS65_LH_OAI21X3 U6280 ( .A(n4613), .B(n3692), .C(n3630), .Z(n3631) );
  HS65_LHS_XNOR2X6 U6281 ( .A(n4173), .B(n4172), .Z(n4174) );
  HS65_LL_NOR2X2 U6283 ( .A(n4665), .B(n4746), .Z(n4666) );
  HS65_LH_OAI21X3 U6284 ( .A(n4330), .B(n4311), .C(n4310), .Z(n4312) );
  HS65_LL_NAND3X2 U6285 ( .A(n3833), .B(n3832), .C(n3831), .Z(n4410) );
  HS65_LH_OAI12X3 U6291 ( .A(n5340), .B(n5339), .C(n5338), .Z(n5359) );
  HS65_LH_IVX9 U6292 ( .A(n3835), .Z(n4563) );
  HS65_LH_AOI21X2 U6295 ( .A(n4352), .B(n4863), .C(n4351), .Z(n4353) );
  HS65_LH_NAND3X5 U6298 ( .A(n5461), .B(n5440), .C(n5470), .Z(n5441) );
  HS65_LH_AO12X4 U6300 ( .A(n5379), .B(n5378), .C(n5377), .Z(n2838) );
  HS65_LH_OAI12X3 U6309 ( .A(n3888), .B(n3887), .C(n3886), .Z(n3889) );
  HS65_LH_OAI21X2 U6311 ( .A(n5214), .B(n5091), .C(n4767), .Z(n5215) );
  HS65_LH_NOR2X3 U6314 ( .A(n4292), .B(n4281), .Z(n3866) );
  HS65_LHS_XNOR2X6 U6315 ( .A(n3876), .B(n4822), .Z(n3877) );
  HS65_LL_OAI12X2 U6319 ( .A(n4747), .B(n4511), .C(n3385), .Z(n3394) );
  HS65_LH_IVX9 U6322 ( .A(n8133), .Z(\u_DataPath/branch_target_i [29]) );
  HS65_LH_AOI21X2 U6323 ( .A(n5237), .B(n5236), .C(n5235), .Z(n5238) );
  HS65_LL_OAI12X2 U6324 ( .A(n5154), .B(n5153), .C(n5152), .Z(n5155) );
  HS65_LH_NOR2AX3 U6325 ( .A(n3246), .B(n3357), .Z(n3358) );
  HS65_LH_AND2X4 U6327 ( .A(n1885), .B(\u_DataPath/toPC2_i [30]), .Z(
        \u_DataPath/branch_target_i [30]) );
  HS65_LH_NOR2AX3 U6328 ( .A(n4904), .B(n4932), .Z(n4905) );
  HS65_LL_NAND2X4 U6329 ( .A(n3197), .B(n4704), .Z(n3199) );
  HS65_LL_NOR2AX3 U6330 ( .A(n3157), .B(n3633), .Z(n3191) );
  HS65_LL_AO12X9 U6332 ( .A(n4184), .B(n2997), .C(n2996), .Z(n4863) );
  HS65_LH_AOI21X2 U6333 ( .A(n5250), .B(n5249), .C(n5248), .Z(n5257) );
  HS65_LH_NAND2X4 U6334 ( .A(n5086), .B(n5117), .Z(n5121) );
  HS65_LH_AOI21X2 U6336 ( .A(n4237), .B(n4239), .C(n3667), .Z(n3668) );
  HS65_LL_AOI12X3 U6338 ( .A(n4239), .B(n3077), .C(n3076), .Z(n4176) );
  HS65_LH_NOR2X6 U6340 ( .A(n5007), .B(n5006), .Z(n5461) );
  HS65_LL_NAND2X4 U6341 ( .A(n4596), .B(n3201), .Z(n4638) );
  HS65_LH_NAND2X2 U6342 ( .A(n5065), .B(n5129), .Z(n5069) );
  HS65_LH_NAND2X4 U6346 ( .A(n5068), .B(n5134), .Z(n5138) );
  HS65_LL_NOR2AX3 U6350 ( .A(n3258), .B(n4079), .Z(n3899) );
  HS65_LH_OAI12X3 U6352 ( .A(n5399), .B(n5398), .C(n5397), .Z(n5400) );
  HS65_LL_IVX7 U6353 ( .A(n4321), .Z(n3326) );
  HS65_LL_NAND3X2 U6354 ( .A(n5355), .B(n5361), .C(n5363), .Z(n5377) );
  HS65_LH_NAND3X3 U6356 ( .A(n4673), .B(n5486), .C(n4573), .Z(n4282) );
  HS65_LL_NAND2AX4 U6357 ( .A(n3249), .B(n4375), .Z(n3454) );
  HS65_LH_NOR4ABX2 U6358 ( .A(n5171), .B(n5164), .C(n5163), .D(n5162), .Z(
        n5168) );
  HS65_LH_CBI4I6X2 U6359 ( .A(n5362), .B(n5388), .C(n5355), .D(n4885), .Z(
        n4886) );
  HS65_LH_AOI21X2 U6363 ( .A(n5412), .B(n5342), .C(n5341), .Z(n5353) );
  HS65_LH_IVX9 U6367 ( .A(n4077), .Z(n3258) );
  HS65_LH_IVX9 U6368 ( .A(n5391), .Z(n5355) );
  HS65_LH_IVX9 U6370 ( .A(n5110), .Z(n4175) );
  HS65_LL_OAI12X3 U6371 ( .A(n4077), .B(n4169), .C(n4078), .Z(n3900) );
  HS65_LL_NAND2X4 U6373 ( .A(n3261), .B(n4259), .Z(n4171) );
  HS65_LL_NAND3X3 U6375 ( .A(n3573), .B(n3572), .C(n3571), .Z(n4832) );
  HS65_LH_NAND3X5 U6378 ( .A(n5459), .B(n5012), .C(n5017), .Z(n5054) );
  HS65_LL_NOR2X2 U6380 ( .A(n4770), .B(n4765), .Z(n2997) );
  HS65_LHS_XOR2X6 U6382 ( .A(n9355), .B(n7637), .Z(
        \u_DataPath/u_execute/link_value_i [31]) );
  HS65_LL_NOR2X3 U6387 ( .A(n3372), .B(n5193), .Z(n4596) );
  HS65_LL_OAI12X2 U6388 ( .A(n4859), .B(n4350), .C(n4861), .Z(n4351) );
  HS65_LH_AOI21X2 U6390 ( .A(n5223), .B(n5222), .C(n5221), .Z(n5224) );
  HS65_LH_NOR3X4 U6391 ( .A(n5439), .B(n5438), .C(n5456), .Z(n5470) );
  HS65_LH_NOR2X3 U6393 ( .A(n4812), .B(n4613), .Z(n4850) );
  HS65_LH_OAI21X2 U6394 ( .A(n5125), .B(n5247), .C(n5434), .Z(n5248) );
  HS65_LH_IVX9 U6397 ( .A(n5107), .Z(n4237) );
  HS65_LH_NAND3X5 U6398 ( .A(n5446), .B(n5445), .C(n5309), .Z(n5318) );
  HS65_LL_OAI12X3 U6400 ( .A(n4578), .B(n3416), .C(n3418), .Z(n4603) );
  HS65_LH_AND2X4 U6403 ( .A(n3886), .B(n3614), .Z(n2858) );
  HS65_LL_NOR2X3 U6405 ( .A(n3756), .B(n3759), .Z(n4823) );
  HS65_LH_NOR2X6 U6407 ( .A(\sub_x_51/A[8] ), .B(n3072), .Z(n4270) );
  HS65_LH_CNIVX3 U6408 ( .A(n4444), .Z(n4445) );
  HS65_LL_OAI12X2 U6409 ( .A(n4861), .B(n4347), .C(n5219), .Z(n2999) );
  HS65_LH_NAND2X4 U6411 ( .A(n5492), .B(n5491), .Z(n5493) );
  HS65_LL_NOR2AX3 U6413 ( .A(n5092), .B(n2995), .Z(n3593) );
  HS65_LH_NOR2X6 U6414 ( .A(n3854), .B(n3853), .Z(n4289) );
  HS65_LH_AOI21X2 U6416 ( .A(n5406), .B(n5405), .C(n5404), .Z(n5410) );
  HS65_LH_OAI21X3 U6417 ( .A(n3379), .B(n5529), .C(n4621), .Z(n4559) );
  HS65_LL_NOR2X2 U6420 ( .A(n4859), .B(n4347), .Z(n3000) );
  HS65_LH_IVX9 U6421 ( .A(n4674), .Z(n4536) );
  HS65_LL_NOR2X2 U6422 ( .A(n4113), .B(n4112), .Z(n4381) );
  HS65_LH_AOI21X2 U6424 ( .A(n5388), .B(n5372), .C(n5371), .Z(n5379) );
  HS65_LH_NAND2X7 U6425 ( .A(n3224), .B(n3223), .Z(n4382) );
  HS65_LL_NOR2X3 U6426 ( .A(n4444), .B(n4447), .Z(n4375) );
  HS65_LL_NAND2X4 U6431 ( .A(\sub_x_51/A[21] ), .B(n3193), .Z(n4460) );
  HS65_LL_NOR2X3 U6433 ( .A(\sub_x_51/A[21] ), .B(n3193), .Z(n4458) );
  HS65_LL_NAND3X3 U6434 ( .A(n5445), .B(n5453), .C(n4011), .Z(n4014) );
  HS65_LL_NAND3X2 U6437 ( .A(n5286), .B(n5292), .C(n5255), .Z(n3992) );
  HS65_LL_NOR2X3 U6439 ( .A(n3128), .B(n3187), .Z(n5245) );
  HS65_LH_NAND2X7 U6441 ( .A(\sub_x_51/A[8] ), .B(n3072), .Z(n4272) );
  HS65_LH_OAI12X3 U6442 ( .A(n5265), .B(n5264), .C(n5147), .Z(n4640) );
  HS65_LL_NAND2X2 U6443 ( .A(n3726), .B(n3725), .Z(n4066) );
  HS65_LH_NAND2X4 U6445 ( .A(n3898), .B(n3897), .Z(n3909) );
  HS65_LH_NOR2X6 U6446 ( .A(n5246), .B(\add_x_50/A[19] ), .Z(n3536) );
  HS65_LH_NAND2X7 U6449 ( .A(\sub_x_51/A[16] ), .B(n5186), .Z(n4448) );
  HS65_LH_NOR2X5 U6453 ( .A(n4630), .B(n4963), .Z(n4534) );
  HS65_LH_IVX9 U6454 ( .A(n4367), .Z(n5294) );
  HS65_LL_HA1X4 U6455 ( .A0(n2849), .B0(n9357), .CO(n7638), .S0(
        \u_DataPath/u_execute/link_value_i [29]) );
  HS65_LH_OAI12X3 U6457 ( .A(n4522), .B(n4519), .C(n4521), .Z(n4686) );
  HS65_LH_NAND3X5 U6461 ( .A(n3346), .B(n3625), .C(n3345), .Z(n4741) );
  HS65_LH_AOI21X2 U6463 ( .A(n5509), .B(n7321), .C(n4654), .Z(n4655) );
  HS65_LL_OAI12X2 U6466 ( .A(n4594), .B(n5191), .C(n5009), .Z(n3202) );
  HS65_LH_AOI21X2 U6467 ( .A(n3941), .B(n5040), .C(n5343), .Z(n3943) );
  HS65_LH_NAND2X4 U6468 ( .A(n5220), .B(n4894), .Z(n4892) );
  HS65_LL_NAND2X4 U6471 ( .A(\lte_x_57/B[4] ), .B(n5208), .Z(n3875) );
  HS65_LH_AOI21X2 U6472 ( .A(n5350), .B(n5334), .C(n5333), .Z(n5339) );
  HS65_LL_NAND2X2 U6473 ( .A(n5009), .B(n4594), .Z(n4931) );
  HS65_LL_NOR2X2 U6480 ( .A(n4818), .B(n4336), .Z(n3255) );
  HS65_LH_NAND2AX7 U6481 ( .A(n5014), .B(n2856), .Z(n5010) );
  HS65_LL_NOR2X3 U6482 ( .A(n3073), .B(n3039), .Z(n4023) );
  HS65_LL_OAI12X2 U6485 ( .A(n5131), .B(n4701), .C(n4703), .Z(n3196) );
  HS65_LH_NAND2X7 U6489 ( .A(n5009), .B(n5008), .Z(n5438) );
  HS65_LH_OAI22X4 U6490 ( .A(n7701), .B(n7791), .C(n7699), .D(n8232), .Z(
        \u_DataPath/data_read_ex_1_i [8]) );
  HS65_LL_NAND2X4 U6493 ( .A(\sub_x_51/A[18] ), .B(n3188), .Z(n4367) );
  HS65_LL_NAND2X5 U6497 ( .A(n3062), .B(n3061), .Z(n5203) );
  HS65_LL_NAND2AX7 U6500 ( .A(n2841), .B(n3141), .Z(n5186) );
  HS65_LL_AO22X4 U6501 ( .A(\lte_x_57/B[28] ), .B(n2796), .C(
        \u_DataPath/u_execute/A_inALU_i[26] ), .D(n4796), .Z(n2854) );
  HS65_LH_AOI211X2 U6502 ( .A(n2798), .B(n8702), .C(n8398), .D(n8397), .Z(
        \u_DataPath/mem_writedata_out_i [9]) );
  HS65_LL_NAND2X5 U6503 ( .A(n3177), .B(n3176), .Z(n5064) );
  HS65_LL_NAND2AX7 U6504 ( .A(n2845), .B(n3144), .Z(n5246) );
  HS65_LH_NAND2X5 U6508 ( .A(\lte_x_57/B[6] ), .B(n3742), .Z(n3730) );
  HS65_LH_NAND2X4 U6510 ( .A(n4882), .B(n4881), .Z(n5220) );
  HS65_LH_OAI22X4 U6514 ( .A(n7701), .B(n7746), .C(n7700), .D(n8312), .Z(
        \u_DataPath/data_read_ex_1_i [31]) );
  HS65_LH_OAI22X4 U6515 ( .A(n7719), .B(n8298), .C(n7718), .D(n8297), .Z(
        \u_DataPath/data_read_ex_2_i [3]) );
  HS65_LH_OAI22X4 U6516 ( .A(n7701), .B(n7812), .C(n7700), .D(n8289), .Z(
        \u_DataPath/data_read_ex_1_i [30]) );
  HS65_LH_OAI22X4 U6517 ( .A(n7701), .B(n7826), .C(n7700), .D(n8295), .Z(
        \u_DataPath/data_read_ex_1_i [28]) );
  HS65_LH_OAI22X4 U6518 ( .A(n7719), .B(n7725), .C(n7718), .D(n8367), .Z(
        \u_DataPath/data_read_ex_2_i [0]) );
  HS65_LH_OAI22X4 U6519 ( .A(n7701), .B(n7854), .C(n7699), .D(n8251), .Z(
        \u_DataPath/data_read_ex_1_i [26]) );
  HS65_LH_OR2X4 U6522 ( .A(n3239), .B(n7321), .Z(n4679) );
  HS65_LL_NAND2X4 U6524 ( .A(\sub_x_51/A[5] ), .B(n3949), .Z(n3758) );
  HS65_LHS_XOR2X3 U6525 ( .A(n8995), .B(n5565), .Z(\u_DataPath/toPC2_i [26])
         );
  HS65_LL_AO12X9 U6528 ( .A(n4880), .B(n8388), .C(n4878), .Z(n5089) );
  HS65_LH_NAND2X7 U6529 ( .A(n8422), .B(n3140), .Z(n3141) );
  HS65_LL_NOR2X2 U6531 ( .A(n4330), .B(n4346), .Z(n5336) );
  HS65_LL_OR2X4 U6533 ( .A(\lte_x_57/B[30] ), .B(n5312), .Z(n4687) );
  HS65_LH_NOR2AX6 U6536 ( .A(n3975), .B(n5190), .Z(n4601) );
  HS65_LH_NAND2X7 U6537 ( .A(n8424), .B(n3133), .Z(n3134) );
  HS65_LH_NAND2X4 U6538 ( .A(n3039), .B(n4796), .Z(n3736) );
  HS65_LL_NAND2X4 U6540 ( .A(n3239), .B(n4208), .Z(n4662) );
  HS65_LL_NOR2X3 U6542 ( .A(\sub_x_51/A[5] ), .B(n3949), .Z(n3756) );
  HS65_LL_AO12X4 U6546 ( .A(n2957), .B(n8370), .C(n3219), .Z(n5508) );
  HS65_LH_OAI22X4 U6547 ( .A(n7719), .B(n7868), .C(n7718), .D(n8276), .Z(
        \u_DataPath/data_read_ex_2_i [15]) );
  HS65_LH_OAI22X4 U6548 ( .A(n7719), .B(n7753), .C(n7717), .D(n8190), .Z(
        \u_DataPath/data_read_ex_2_i [17]) );
  HS65_LH_OAI22X4 U6549 ( .A(n7701), .B(n7889), .C(n7700), .D(n8285), .Z(
        \u_DataPath/data_read_ex_1_i [22]) );
  HS65_LH_OAI22X4 U6550 ( .A(n7701), .B(n7798), .C(n7699), .D(n8247), .Z(
        \u_DataPath/data_read_ex_1_i [6]) );
  HS65_LH_OAI22X4 U6551 ( .A(n7701), .B(n7732), .C(n7699), .D(n8235), .Z(
        \u_DataPath/data_read_ex_1_i [10]) );
  HS65_LH_OAI22X4 U6552 ( .A(n7701), .B(n7910), .C(n7700), .D(n8265), .Z(
        \u_DataPath/data_read_ex_1_i [5]) );
  HS65_LH_OAI22X4 U6553 ( .A(n7719), .B(n7819), .C(n7718), .D(n8274), .Z(
        \u_DataPath/data_read_ex_2_i [20]) );
  HS65_LH_OAI22X4 U6554 ( .A(n7701), .B(n7819), .C(n7700), .D(n8292), .Z(
        \u_DataPath/data_read_ex_1_i [20]) );
  HS65_LH_OAI22X4 U6555 ( .A(n7701), .B(n7770), .C(n7699), .D(n8261), .Z(
        \u_DataPath/data_read_ex_1_i [9]) );
  HS65_LH_OAI22X4 U6556 ( .A(n7719), .B(n7903), .C(n7717), .D(n8199), .Z(
        \u_DataPath/data_read_ex_2_i [21]) );
  HS65_LH_OAI22X4 U6557 ( .A(n7701), .B(n7868), .C(n7700), .D(n8303), .Z(
        \u_DataPath/data_read_ex_1_i [15]) );
  HS65_LH_OAI22X4 U6558 ( .A(n7719), .B(n7763), .C(n7717), .D(n8236), .Z(
        \u_DataPath/data_read_ex_2_i [12]) );
  HS65_LH_OAI22X4 U6559 ( .A(n7701), .B(n7763), .C(n7699), .D(n8240), .Z(
        \u_DataPath/data_read_ex_1_i [12]) );
  HS65_LH_OAI22X4 U6560 ( .A(n7701), .B(n7840), .C(n7699), .D(n8256), .Z(
        \u_DataPath/data_read_ex_1_i [25]) );
  HS65_LH_OAI22X4 U6561 ( .A(n7701), .B(n7861), .C(n7699), .D(n8254), .Z(
        \u_DataPath/data_read_ex_1_i [14]) );
  HS65_LH_OAI22X4 U6562 ( .A(n7701), .B(n7833), .C(n7700), .D(n8319), .Z(
        \u_DataPath/data_read_ex_1_i [29]) );
  HS65_LH_NOR2X3 U6564 ( .A(n4918), .B(n3338), .Z(n3827) );
  HS65_LL_NAND2X4 U6567 ( .A(n2978), .B(n2831), .Z(n2979) );
  HS65_LH_NAND2AX7 U6569 ( .A(n8610), .B(n2797), .Z(n8431) );
  HS65_LH_NAND2AX7 U6570 ( .A(n8647), .B(n2797), .Z(n7329) );
  HS65_LH_NOR2X3 U6571 ( .A(n5529), .B(n3338), .Z(n3716) );
  HS65_LL_OR2X18 U6572 ( .A(n9538), .B(n3222), .Z(n2829) );
  HS65_LH_NOR2X5 U6573 ( .A(n4189), .B(n3338), .Z(n5495) );
  HS65_LH_NAND2AX7 U6574 ( .A(n8630), .B(n2797), .Z(n8437) );
  HS65_LH_NAND2AX7 U6577 ( .A(n8661), .B(n2797), .Z(n8422) );
  HS65_LH_NOR2X2 U6580 ( .A(n5497), .B(n2968), .Z(n5213) );
  HS65_LL_OAI12X5 U6581 ( .A(n8391), .B(n2934), .C(n2933), .Z(n4346) );
  HS65_LL_OAI22X1 U6583 ( .A(n6861), .B(n8226), .C(n7716), .D(n8064), .Z(
        \u_DataPath/data_read_ex_2_i [7]) );
  HS65_LH_AOI22X3 U6585 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][8] ), .B(n9188), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][8] ), .D(
        n9190), .Z(n6650) );
  HS65_LH_OAI22X4 U6586 ( .A(n7701), .B(n8226), .C(n7699), .D(n8225), .Z(
        \u_DataPath/data_read_ex_1_i [7]) );
  HS65_LH_OAI22X4 U6587 ( .A(n7719), .B(n8282), .C(n7718), .D(n8281), .Z(
        \u_DataPath/data_read_ex_2_i [2]) );
  HS65_LL_OAI12X3 U6588 ( .A(n9127), .B(n5584), .C(n9025), .Z(n5729) );
  HS65_LH_IVX18 U6595 ( .A(n3338), .Z(n2792) );
  HS65_LH_AOI22X3 U6598 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][31] ), .B(n9206), 
        .C(n9205), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][31] ), .Z(n7499)
         );
  HS65_LH_AOI22X3 U6601 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][0] ), .B(n9248), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][0] ), .D(
        n9240), .Z(n6209) );
  HS65_LH_AO22X4 U6602 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][31] ), .B(n9469), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][31] ), .D(
        n9475), .Z(n6608) );
  HS65_LH_AOI22X3 U6603 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][31] ), .B(n9255), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][31] ), .D(
        n9195), .Z(n6605) );
  HS65_LH_AOI22X3 U6605 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][30] ), .B(n9255), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][30] ), .D(
        n9195), .Z(n6565) );
  HS65_LH_AO22X4 U6606 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][30] ), .B(n9469), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][30] ), .D(
        n9475), .Z(n6568) );
  HS65_LH_AO22X4 U6607 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][31] ), .B(n9364), 
        .C(n9253), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][31] ), .Z(n7522)
         );
  HS65_LH_AOI22X3 U6608 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][31] ), .B(n9250), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][31] ), .D(
        n9265), .Z(n7506) );
  HS65_LL_IVX7 U6611 ( .A(n3940), .Z(n4871) );
  HS65_LH_OAI31X5 U6616 ( .A(\u_DataPath/dataOut_exe_i [1]), .B(n8222), .C(
        n8164), .D(n8302), .Z(n8307) );
  HS65_LH_OAI21X2 U6617 ( .A(n8071), .B(n8586), .C(n8359), .Z(n7952) );
  HS65_LH_CBI4I6X2 U6618 ( .A(n9419), .B(n7973), .C(n7968), .D(n7974), .Z(
        n7969) );
  HS65_LL_NOR2AX6 U6619 ( .A(n3118), .B(n3117), .Z(\lte_x_57/B[28] ) );
  HS65_LH_OAI22X3 U6620 ( .A(n9317), .B(n8071), .C(n7978), .D(n8363), .Z(n7980) );
  HS65_LL_IVX4 U6621 ( .A(\lte_x_57/B[7] ), .Z(n4330) );
  HS65_LH_AOI22X1 U6624 ( .A(n9243), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][17] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][17] ), .D(n9009), 
        .Z(n5947) );
  HS65_LH_AO22X9 U6626 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][20] ), .B(n9363), 
        .C(n9097), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][20] ), .Z(n7111)
         );
  HS65_LH_AOI22X1 U6627 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][20] ), .B(n9188), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][20] ), .D(
        n8854), .Z(n6589) );
  HS65_LH_AO22X9 U6628 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][16] ), .B(n9469), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][16] ), .D(
        n9475), .Z(n6171) );
  HS65_LH_AOI22X1 U6629 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][18] ), .B(n9096), 
        .C(n9158), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][18] ), .Z(n7220)
         );
  HS65_LH_AO22X9 U6631 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][21] ), .B(n9363), 
        .C(n9257), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][21] ), .Z(n6009)
         );
  HS65_LH_AOI22X3 U6632 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][5] ), .B(n9255), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][5] ), .D(
        n9195), .Z(n6625) );
  HS65_LH_AOI22X3 U6634 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][24] ), .B(n9191), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][24] ), .D(
        n9471), .Z(n6271) );
  HS65_LH_AO22X9 U6636 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][17] ), .B(n9363), 
        .C(n9257), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][17] ), .Z(n5967)
         );
  HS65_LH_AO22X9 U6637 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][16] ), .B(n9363), 
        .C(n9097), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][16] ), .Z(n6075)
         );
  HS65_LH_AOI22X1 U6643 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][1] ), .B(n9096), 
        .C(n9158), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][1] ), .Z(n7240)
         );
  HS65_LH_AOI22X3 U6645 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][16] ), .B(n9226), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][16] ), .D(
        n9193), .Z(n6190) );
  HS65_LH_AOI22X3 U6646 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][16] ), .B(n9248), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][16] ), .D(
        n9240), .Z(n6189) );
  HS65_LH_AOI22X3 U6650 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][22] ), .B(n9255), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][22] ), .D(
        n9195), .Z(n6545) );
  HS65_LH_AO22X4 U6652 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][5] ), .B(n9469), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][5] ), .D(
        n9475), .Z(n6628) );
  HS65_LH_AOI22X1 U6653 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][5] ), .B(n9188), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][5] ), .D(
        n8854), .Z(n6629) );
  HS65_LH_AO22X9 U6654 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][14] ), .B(n9363), 
        .C(n9097), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][14] ), .Z(n6095)
         );
  HS65_LH_AOI22X3 U6660 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][23] ), .B(n9191), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][23] ), .D(
        n9471), .Z(n6337) );
  HS65_LH_AOI22X3 U6662 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][23] ), .B(n8938), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][23] ), .D(
        n9264), .Z(n6342) );
  HS65_LH_AOI22X3 U6663 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][15] ), .B(n8950), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][15] ), .D(
        n9471), .Z(n6889) );
  HS65_LH_AOI22X3 U6665 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][11] ), .B(n8938), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][11] ), .D(
        n9264), .Z(n6509) );
  HS65_LH_AOI22X3 U6667 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][11] ), .B(n9191), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][11] ), .D(
        n9471), .Z(n6507) );
  HS65_LH_AOI22X3 U6669 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][27] ), .B(n9246), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][27] ), .D(
        n9262), .Z(n6317) );
  HS65_LH_AOI22X3 U6674 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][14] ), .B(n9191), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][14] ), .D(
        n9471), .Z(n6869) );
  HS65_LL_NAND3AX3 U6676 ( .A(n3218), .B(n3217), .C(n3216), .Z(n3221) );
  HS65_LL_NAND2X4 U6678 ( .A(addr_to_iram_26), .B(n7406), .Z(n7605) );
  HS65_LH_IVX7 U6679 ( .A(n8103), .Z(\u_DataPath/pc4_to_idexreg_i [14]) );
  HS65_LL_NAND2X2 U6680 ( .A(n8419), .B(n3042), .Z(n3044) );
  HS65_LL_NOR2X3 U6681 ( .A(n2967), .B(n2966), .Z(n3940) );
  HS65_LH_NAND2X4 U6682 ( .A(n8798), .B(n8513), .Z(n7974) );
  HS65_LH_NOR2X6 U6683 ( .A(n8676), .B(n3181), .Z(n2985) );
  HS65_LL_NAND3X5 U6688 ( .A(n8727), .B(n2813), .C(n8186), .Z(n8302) );
  HS65_LHS_XNOR2X6 U6689 ( .A(n7390), .B(n7406), .Z(\u_DataPath/pc_4_i [28])
         );
  HS65_LH_NOR2X6 U6690 ( .A(n8631), .B(n3181), .Z(n3037) );
  HS65_LL_AO12X4 U6691 ( .A(n8698), .B(n2710), .C(n3064), .Z(n3065) );
  HS65_LHS_XOR2X3 U6693 ( .A(n8999), .B(n5842), .Z(
        \u_DataPath/u_execute/resAdd1_i [23]) );
  HS65_LHS_XOR2X3 U6694 ( .A(n8922), .B(n5641), .Z(\u_DataPath/toPC2_i [22])
         );
  HS65_LH_AOI22X1 U6695 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][2] ), .B(n9098), 
        .C(n9200), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][2] ), .Z(n6145)
         );
  HS65_LH_AOI22X3 U6697 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][4] ), .B(n9250), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][4] ), .D(n9265), .Z(n6033) );
  HS65_LH_AOI22X3 U6700 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][4] ), .B(n9206), 
        .C(n9205), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][4] ), .Z(n6021)
         );
  HS65_LH_AOI22X3 U6701 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][4] ), .B(n9204), 
        .C(n9203), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][4] ), .Z(n6020)
         );
  HS65_LHS_XOR2X6 U6705 ( .A(n7455), .B(n7454), .Z(\u_DataPath/pc_4_i [16]) );
  HS65_LH_AOI21X2 U6707 ( .A(n8725), .B(n9076), .C(n8071), .Z(n7975) );
  HS65_LL_NAND2AX4 U6708 ( .A(n2959), .B(n9018), .Z(n8374) );
  HS65_LH_NAND2X5 U6709 ( .A(n1885), .B(n8961), .Z(n8084) );
  HS65_LH_AOI12X2 U6710 ( .A(n9388), .B(n5884), .C(n9461), .Z(n5837) );
  HS65_LH_AOI12X2 U6712 ( .A(n9396), .B(n5884), .C(n9437), .Z(n5830) );
  HS65_LH_NOR2X5 U6719 ( .A(n8669), .B(n3149), .Z(n2966) );
  HS65_LH_NOR2X5 U6723 ( .A(n8667), .B(n3149), .Z(n3158) );
  HS65_LL_NAND2X2 U6724 ( .A(n3215), .B(n9018), .Z(n3217) );
  HS65_LL_NAND2X4 U6725 ( .A(addr_to_iram_24), .B(n7389), .Z(n7473) );
  HS65_LH_NOR2X5 U6727 ( .A(n9463), .B(n3018), .Z(n8400) );
  HS65_LH_NOR2X6 U6728 ( .A(n9268), .B(n3178), .Z(n2928) );
  HS65_LL_NAND2X2 U6729 ( .A(n8724), .B(n2710), .Z(n3004) );
  HS65_LH_NOR2X5 U6731 ( .A(n9401), .B(n3028), .Z(n8393) );
  HS65_LH_NOR2X5 U6732 ( .A(\u_DataPath/dataOut_exe_i [27]), .B(n3178), .Z(
        n3102) );
  HS65_LL_NAND2AX4 U6733 ( .A(n2949), .B(n2948), .Z(n8382) );
  HS65_LH_NAND2X7 U6735 ( .A(n8774), .B(n2712), .Z(n3237) );
  HS65_LL_NAND2X2 U6736 ( .A(n2710), .B(n8263), .Z(n2936) );
  HS65_LL_NAND2AX7 U6737 ( .A(n2899), .B(n2898), .Z(n3214) );
  HS65_LL_OAI12X3 U6738 ( .A(n8045), .B(n8043), .C(n1885), .Z(n8044) );
  HS65_LH_OAI12X3 U6739 ( .A(n9129), .B(n5902), .C(n8974), .Z(n5904) );
  HS65_LH_OAI12X3 U6740 ( .A(n8888), .B(n5894), .C(n8977), .Z(n5896) );
  HS65_LH_OAI12X3 U6741 ( .A(n9312), .B(n5894), .C(n9237), .Z(n5888) );
  HS65_LHS_XNOR2X6 U6742 ( .A(n7381), .B(n7467), .Z(\u_DataPath/pc_4_i [22])
         );
  HS65_LH_BFX18 U6744 ( .A(n7708), .Z(n7706) );
  HS65_LHS_XNOR2X6 U6745 ( .A(n7375), .B(n7371), .Z(\u_DataPath/pc_4_i [24])
         );
  HS65_LH_NOR2X5 U6746 ( .A(n7453), .B(n7452), .Z(n7372) );
  HS65_LH_NOR2X5 U6747 ( .A(n7357), .B(n7356), .Z(n7358) );
  HS65_LHS_XNOR2X6 U6748 ( .A(n9216), .B(n9181), .Z(
        \u_DataPath/u_execute/link_value_i [10]) );
  HS65_LH_NOR2X5 U6749 ( .A(\u_DataPath/dataOut_exe_i [20]), .B(n3980), .Z(
        n8432) );
  HS65_LH_NAND2X4 U6750 ( .A(n3090), .B(n8396), .Z(n3035) );
  HS65_LL_OAI12X12 U6751 ( .A(n8010), .B(n8004), .C(n1885), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N151 ) );
  HS65_LH_NAND2X4 U6753 ( .A(n3090), .B(n8395), .Z(n3030) );
  HS65_LL_NOR2AX3 U6754 ( .A(n2897), .B(n2916), .Z(n2898) );
  HS65_LH_NOR2X5 U6755 ( .A(\u_DataPath/dataOut_exe_i [19]), .B(n3980), .Z(
        n8429) );
  HS65_LHS_XOR2X6 U6757 ( .A(n7449), .B(n7448), .Z(\u_DataPath/pc_4_i [12]) );
  HS65_LH_NAND3X5 U6758 ( .A(Data_out_fromRAM[31]), .B(n8164), .C(n2813), .Z(
        n7314) );
  HS65_LH_NOR3X4 U6759 ( .A(\u_DataPath/dataOut_exe_i [1]), .B(n8220), .C(
        n8164), .Z(n7312) );
  HS65_LH_NAND2X4 U6760 ( .A(n3090), .B(n8425), .Z(n3132) );
  HS65_LH_OR2X9 U6761 ( .A(n8727), .B(n9144), .Z(n8454) );
  HS65_LH_NOR2X5 U6763 ( .A(\u_DataPath/dataOut_exe_i [18]), .B(n3980), .Z(
        n8426) );
  HS65_LL_NAND2X4 U6764 ( .A(n3090), .B(n8371), .Z(n3218) );
  HS65_LHS_XNOR2X6 U6768 ( .A(n7345), .B(n7464), .Z(\u_DataPath/pc_4_i [8]) );
  HS65_LL_NOR2AX3 U6770 ( .A(n1885), .B(n7674), .Z(n7660) );
  HS65_LL_NOR2X3 U6772 ( .A(n2910), .B(n2894), .Z(n2897) );
  HS65_LH_NOR2X5 U6773 ( .A(n7617), .B(n7616), .Z(n7418) );
  HS65_LH_NAND3X5 U6776 ( .A(opcode_i[0]), .B(n7411), .C(n7403), .Z(n7409) );
  HS65_LH_AOI21X6 U6777 ( .A(n3148), .B(\u_DataPath/from_mem_data_out_i [26]), 
        .C(n3108), .Z(n7659) );
  HS65_LH_NOR2X3 U6778 ( .A(\u_DataPath/dataOut_exe_i [14]), .B(n2782), .Z(
        n8414) );
  HS65_LL_NAND2AX14 U6779 ( .A(n2884), .B(n2883), .Z(n3234) );
  HS65_LH_NOR2X5 U6780 ( .A(n7447), .B(n7446), .Z(n7338) );
  HS65_LH_NAND2X4 U6781 ( .A(n5912), .B(n5911), .Z(n5917) );
  HS65_LL_NOR2X6 U6782 ( .A(n6188), .B(n6183), .Z(n6345) );
  HS65_LH_IVX7 U6783 ( .A(n7613), .Z(n7397) );
  HS65_LH_NOR2X6 U6784 ( .A(n5959), .B(n5952), .Z(n6110) );
  HS65_LH_AO22X9 U6785 ( .A(n9360), .B(n7944), .C(n8906), .D(n7943), .Z(
        \u_DataPath/RFaddr_out_memwb_i [4]) );
  HS65_LH_AO22X9 U6786 ( .A(n9452), .B(n7944), .C(n8819), .D(n7943), .Z(
        \u_DataPath/RFaddr_out_memwb_i [1]) );
  HS65_LH_AO22X9 U6787 ( .A(n9435), .B(n7944), .C(n9046), .D(n7943), .Z(
        \u_DataPath/RFaddr_out_memwb_i [2]) );
  HS65_LH_AO22X9 U6788 ( .A(n9436), .B(n7944), .C(n8820), .D(n7943), .Z(
        \u_DataPath/RFaddr_out_memwb_i [0]) );
  HS65_LH_AO22X9 U6789 ( .A(n9434), .B(n7944), .C(n9112), .D(n7943), .Z(
        \u_DataPath/RFaddr_out_memwb_i [3]) );
  HS65_LH_OAI12X3 U6791 ( .A(n9085), .B(n9238), .C(n9086), .Z(n5713) );
  HS65_LH_IVX7 U6792 ( .A(n7608), .Z(n7332) );
  HS65_LLS_XNOR2X3 U6793 ( .A(\u_DataPath/idex_rt_i [0]), .B(n3529), .Z(n2915)
         );
  HS65_LH_NAND3X5 U6794 ( .A(n7964), .B(n7399), .C(n7404), .Z(n7410) );
  HS65_LLS_XNOR2X3 U6795 ( .A(n8812), .B(n9059), .Z(n6490) );
  HS65_LLS_XNOR2X3 U6796 ( .A(\u_DataPath/idex_rt_i [2]), .B(n6488), .Z(n2896)
         );
  HS65_LLS_XNOR2X3 U6797 ( .A(\u_DataPath/idex_rt_i [4]), .B(n8029), .Z(n2895)
         );
  HS65_LH_OAI12X3 U6798 ( .A(n8887), .B(n5914), .C(n8985), .Z(n5916) );
  HS65_LLS_XNOR2X3 U6799 ( .A(n2872), .B(n8028), .Z(n2873) );
  HS65_LH_NOR2X5 U6801 ( .A(n3435), .B(n7351), .Z(n3437) );
  HS65_LH_NOR3X4 U6802 ( .A(\u_DataPath/cw_tomem_i [7]), .B(
        \u_DataPath/cw_tomem_i [8]), .C(n7351), .Z(n8163) );
  HS65_LH_NAND2X4 U6803 ( .A(n5786), .B(n5785), .Z(n5788) );
  HS65_LH_IVX18 U6804 ( .A(n8310), .Z(n8315) );
  HS65_LH_NAND2X4 U6805 ( .A(n5892), .B(n5891), .Z(n5897) );
  HS65_LH_NAND2X4 U6806 ( .A(n5907), .B(n5906), .Z(n5909) );
  HS65_LH_NAND2X7 U6807 ( .A(n5623), .B(n5626), .Z(n5632) );
  HS65_LH_NOR2X5 U6808 ( .A(n8466), .B(\u_DataPath/pc_4_to_ex_i [3]), .Z(n5707) );
  HS65_LH_NAND2X4 U6809 ( .A(n5913), .B(n5858), .Z(n5860) );
  HS65_LH_NAND2X4 U6810 ( .A(n5863), .B(n5862), .Z(n5864) );
  HS65_LH_NAND2X7 U6811 ( .A(n5542), .B(n5571), .Z(n5544) );
  HS65_LH_IVX7 U6813 ( .A(n5774), .Z(n5780) );
  HS65_LH_NAND2X4 U6814 ( .A(n5767), .B(n5766), .Z(n5769) );
  HS65_LH_NAND2X4 U6815 ( .A(n5583), .B(n5582), .Z(n5585) );
  HS65_LH_NAND2X4 U6816 ( .A(n5883), .B(n5882), .Z(n5885) );
  HS65_LH_NAND2X4 U6817 ( .A(n5841), .B(n5840), .Z(n5843) );
  HS65_LL_AND2X4 U6818 ( .A(n3435), .B(n3436), .Z(n7352) );
  HS65_LH_NOR2X6 U6819 ( .A(n7340), .B(n7344), .Z(n7341) );
  HS65_LH_NAND2X7 U6820 ( .A(n5743), .B(n5774), .Z(n5745) );
  HS65_LH_NAND2X7 U6821 ( .A(n8466), .B(\u_DataPath/pc_4_to_ex_i [3]), .Z(
        n5912) );
  HS65_LH_NOR2X6 U6822 ( .A(n2804), .B(n8017), .Z(n5944) );
  HS65_LLS_XNOR2X3 U6823 ( .A(\u_DataPath/rs_ex_i [0]), .B(n3528), .Z(n2874)
         );
  HS65_LH_NOR2X6 U6825 ( .A(n7366), .B(n7384), .Z(n7367) );
  HS65_LHS_XNOR2X6 U6826 ( .A(addr_to_iram_0), .B(n7330), .Z(
        \u_DataPath/pc_4_i [3]) );
  HS65_LH_NOR2X3 U6827 ( .A(n7965), .B(opcode_i[4]), .Z(n7929) );
  HS65_LL_NAND3X2 U6828 ( .A(n8019), .B(n7965), .C(n7933), .Z(n7934) );
  HS65_LH_NAND2X4 U6829 ( .A(n5564), .B(n5563), .Z(n5566) );
  HS65_LH_NAND3X5 U6831 ( .A(opcode_i[2]), .B(opcode_i[4]), .C(n8070), .Z(
        n7608) );
  HS65_LL_NAND4ABX3 U6833 ( .A(\u_DataPath/regfile_addr_out_towb_i [3]), .B(
        \u_DataPath/regfile_addr_out_towb_i [4]), .C(n3528), .D(n7310), .Z(
        n2892) );
  HS65_LH_NOR2X3 U6834 ( .A(n9221), .B(rst), .Z(\u_DataPath/rs_ex_i [3]) );
  HS65_LH_NOR2X5 U6835 ( .A(opcode_i[5]), .B(opcode_i[3]), .Z(n8070) );
  HS65_LH_OAI12X3 U6836 ( .A(n5877), .B(n5874), .C(n5876), .Z(n5748) );
  HS65_LH_OAI12X3 U6838 ( .A(n5685), .B(n5589), .C(n5591), .Z(n5539) );
  HS65_LL_NOR3X1 U6839 ( .A(opcode_i[3]), .B(opcode_i[1]), .C(opcode_i[4]), 
        .Z(n7933) );
  HS65_LH_IVX7 U6840 ( .A(n5871), .Z(n5781) );
  HS65_LH_NAND2X4 U6841 ( .A(n5728), .B(n5727), .Z(n5730) );
  HS65_LH_NAND2X4 U6842 ( .A(n5720), .B(n5719), .Z(n5722) );
  HS65_LL_AND2X4 U6843 ( .A(n8162), .B(n3433), .Z(n3436) );
  HS65_LH_NOR2X6 U6844 ( .A(n5898), .B(n5903), .Z(n5737) );
  HS65_LH_NAND2X7 U6845 ( .A(n5733), .B(n5732), .Z(n5759) );
  HS65_LH_IVX7 U6846 ( .A(n5887), .Z(n5805) );
  HS65_LL_NAND4ABX3 U6847 ( .A(\u_DataPath/RFaddr_out_memwb_i [0]), .B(
        \u_DataPath/RFaddr_out_memwb_i [1]), .C(n2880), .D(n8027), .Z(n2881)
         );
  HS65_LH_IVX7 U6848 ( .A(n5681), .Z(n5620) );
  HS65_LH_IVX4 U6849 ( .A(n5907), .Z(n5855) );
  HS65_LH_NAND2X4 U6850 ( .A(\u_DataPath/immediate_ext_dec_i [0]), .B(
        \u_DataPath/immediate_ext_dec_i [1]), .Z(n7982) );
  HS65_LH_IVX7 U6851 ( .A(n5677), .Z(n5578) );
  HS65_LH_NOR2X6 U6852 ( .A(n5851), .B(n5854), .Z(n5849) );
  HS65_LH_IVX7 U6853 ( .A(n5811), .Z(n5812) );
  HS65_LH_OAI12X3 U6854 ( .A(n5811), .B(n5808), .C(n5810), .Z(n5778) );
  HS65_LH_NAND2X4 U6855 ( .A(n5923), .B(n5922), .Z(n5925) );
  HS65_LH_NAND2X4 U6857 ( .A(n5927), .B(n5926), .Z(n5929) );
  HS65_LH_OAI12X3 U6858 ( .A(n5664), .B(n5660), .C(n5662), .Z(n5658) );
  HS65_LH_OAI12X3 U6859 ( .A(n5893), .B(n5890), .C(n5892), .Z(n5802) );
  HS65_LH_NAND3X5 U6860 ( .A(\u_DataPath/cw_tomem_i [8]), .B(n3435), .C(n3429), 
        .Z(n3430) );
  HS65_LH_NAND2X7 U6861 ( .A(n8465), .B(\u_DataPath/pc_4_to_ex_i [2]), .Z(
        n5913) );
  HS65_LH_NOR2X5 U6862 ( .A(\u_DataPath/idex_rt_i [3]), .B(
        \u_DataPath/pc_4_to_ex_i [19]), .Z(n5874) );
  HS65_LLS_XOR2X3 U6863 ( .A(n8515), .B(\u_DataPath/RFaddr_out_memwb_i [4]), 
        .Z(n2884) );
  HS65_LH_NAND2X7 U6864 ( .A(n8510), .B(\u_DataPath/pc_4_to_ex_i [13]), .Z(
        n5810) );
  HS65_LH_IVX9 U6865 ( .A(n7648), .Z(\u_DataPath/regfile_addr_out_towb_i [3])
         );
  HS65_LH_NOR2X5 U6866 ( .A(n8469), .B(\u_DataPath/pc_4_to_ex_i [10]), .Z(
        n5592) );
  HS65_LH_NAND2X4 U6867 ( .A(n8515), .B(\u_DataPath/pc_4_to_ex_i [31]), .Z(
        n5733) );
  HS65_LH_NOR2X5 U6868 ( .A(n8515), .B(\u_DataPath/pc_4_to_ex_i [29]), .Z(
        n5760) );
  HS65_LH_OR2X9 U6869 ( .A(n8515), .B(\u_DataPath/pc_4_to_ex_i [28]), .Z(n5926) );
  HS65_LH_NOR2X5 U6870 ( .A(n8515), .B(\u_DataPath/pc_4_to_ex_i [27]), .Z(
        n5765) );
  HS65_LH_OR2X9 U6871 ( .A(n8515), .B(\u_DataPath/pc_4_to_ex_i [26]), .Z(n5918) );
  HS65_LH_NOR2X5 U6872 ( .A(n8525), .B(\u_DataPath/pc_4_to_ex_i [9]), .Z(n5688) );
  HS65_LH_NOR2X5 U6873 ( .A(n8526), .B(\u_DataPath/pc_4_to_ex_i [19]), .Z(
        n5629) );
  HS65_LH_NOR2X5 U6874 ( .A(n8526), .B(\u_DataPath/pc_4_to_ex_i [28]), .Z(
        n5557) );
  HS65_LH_NAND2X7 U6875 ( .A(n8506), .B(\u_DataPath/pc_4_to_ex_i [11]), .Z(
        n5799) );
  HS65_LH_NOR2X5 U6876 ( .A(n8526), .B(\u_DataPath/pc_4_to_ex_i [30]), .Z(
        n5669) );
  HS65_LH_NAND2X4 U6877 ( .A(n8526), .B(\u_DataPath/pc_4_to_ex_i [31]), .Z(
        n5666) );
  HS65_LH_NAND2X7 U6878 ( .A(n8524), .B(\u_DataPath/pc_4_to_ex_i [8]), .Z(
        n5893) );
  HS65_LH_OR2X9 U6879 ( .A(\u_DataPath/rs_ex_i [0]), .B(
        \u_DataPath/pc_4_to_ex_i [21]), .Z(n5817) );
  HS65_LLS_XNOR2X6 U6880 ( .A(\u_DataPath/idex_rt_i [0]), .B(
        \u_DataPath/RFaddr_out_memwb_i [0]), .Z(n2907) );
  HS65_LLS_XNOR2X3 U6881 ( .A(\u_DataPath/idex_rt_i [2]), .B(
        \u_DataPath/RFaddr_out_memwb_i [2]), .Z(n2905) );
  HS65_LH_NOR2X5 U6882 ( .A(\u_DataPath/idex_rt_i [4]), .B(
        \u_DataPath/pc_4_to_ex_i [20]), .Z(n5823) );
  HS65_LH_NAND2X7 U6883 ( .A(n8523), .B(\u_DataPath/pc_4_to_ex_i [6]), .Z(
        n5901) );
  HS65_LH_NAND2X7 U6884 ( .A(n8467), .B(\u_DataPath/pc_4_to_ex_i [4]), .Z(
        n5907) );
  HS65_LH_OR2X9 U6885 ( .A(n8526), .B(\u_DataPath/pc_4_to_ex_i [25]), .Z(n5727) );
  HS65_LH_NOR2X5 U6886 ( .A(\u_DataPath/cw_tomem_i [8]), .B(
        \u_DataPath/cw_tomem_i [6]), .Z(n3433) );
  HS65_LH_IVX9 U6887 ( .A(\u_DataPath/cw_to_ex_i [19]), .Z(n8358) );
  HS65_LH_IVX9 U6888 ( .A(\u_DataPath/dataOut_exe_i [7]), .Z(n8455) );
  HS65_LH_NOR2X5 U6891 ( .A(n8524), .B(\u_DataPath/pc_4_to_ex_i [8]), .Z(n5692) );
  HS65_LH_NOR2X5 U6892 ( .A(n8523), .B(\u_DataPath/pc_4_to_ex_i [6]), .Z(n5700) );
  HS65_LH_NOR2X5 U6893 ( .A(\u_DataPath/pc_4_to_ex_i [5]), .B(n8522), .Z(n5650) );
  HS65_LH_NOR2X5 U6894 ( .A(n8474), .B(\u_DataPath/pc_4_to_ex_i [7]), .Z(n5695) );
  HS65_LL_OAI12X3 U6895 ( .A(n7664), .B(n7665), .C(n7663), .Z(n7652) );
  HS65_LL_NAND3X3 U6896 ( .A(n9142), .B(n8357), .C(n5530), .Z(n7665) );
  HS65_LL_CBI4I1X3 U6904 ( .A(n8970), .B(n8757), .C(n9044), .D(n8594), .Z(
        \u_DataPath/dataOut_exe_i [28]) );
  HS65_LL_NOR2AX3 U6907 ( .A(n8351), .B(n8348), .Z(n4100) );
  HS65_LL_NAND3AX3 U6908 ( .A(n8338), .B(n8340), .C(n8341), .Z(n3882) );
  HS65_LH_AOI12X6 U6909 ( .A(n9269), .B(n8356), .C(n7712), .Z(n7658) );
  HS65_LL_NAND2AX4 U6910 ( .A(n4497), .B(n4496), .Z(n4498) );
  HS65_LL_NAND2AX4 U6912 ( .A(n5060), .B(n5059), .Z(n5061) );
  HS65_LL_OAI21X2 U6914 ( .A(n8310), .B(n8351), .C(n8258), .Z(
        \u_DataPath/dataOut_exe_i [9]) );
  HS65_LL_AO112X4 U6915 ( .A(n7325), .B(n4395), .C(n4394), .D(n4393), .Z(n4396) );
  HS65_LHS_XNOR2X6 U6917 ( .A(n4139), .B(n4138), .Z(n4140) );
  HS65_LL_AO12X4 U6919 ( .A(n4671), .B(n4062), .C(n3816), .Z(n2852) );
  HS65_LLS_XNOR2X3 U6921 ( .A(n3281), .B(n3280), .Z(n3282) );
  HS65_LLS_XNOR2X3 U6922 ( .A(n4418), .B(n4417), .Z(n4419) );
  HS65_LL_NOR4ABX4 U6923 ( .A(n3655), .B(n3654), .C(n3653), .D(n2861), .Z(
        n3656) );
  HS65_LL_NOR2AX3 U6924 ( .A(n3498), .B(n3497), .Z(n3503) );
  HS65_LLS_XNOR2X3 U6926 ( .A(n3364), .B(n3363), .Z(n3365) );
  HS65_LL_NAND3AX3 U6927 ( .A(n3873), .B(n3872), .C(n3871), .Z(n3879) );
  HS65_LL_OAI12X2 U6928 ( .A(n4492), .B(n4695), .C(n4491), .Z(n4493) );
  HS65_LL_NOR2AX3 U6930 ( .A(n3748), .B(n3747), .Z(n3749) );
  HS65_LLS_XNOR2X3 U6931 ( .A(n2847), .B(n4450), .Z(n4451) );
  HS65_LL_AOI21X2 U6933 ( .A(n5517), .B(n4993), .C(n4409), .Z(n4422) );
  HS65_LLS_XNOR2X3 U6935 ( .A(n3500), .B(n3499), .Z(n3501) );
  HS65_LLS_XNOR2X3 U6937 ( .A(n4735), .B(n4734), .Z(n4736) );
  HS65_LL_OAI12X2 U6938 ( .A(n4463), .B(n4714), .C(n4462), .Z(n4464) );
  HS65_LH_OAI21X3 U6941 ( .A(n4846), .B(n3200), .C(n4561), .Z(n4566) );
  HS65_LL_OAI12X2 U6943 ( .A(n3635), .B(n4714), .C(n3634), .Z(n3638) );
  HS65_LL_AOI21X2 U6944 ( .A(n5510), .B(n4570), .C(n3461), .Z(n3481) );
  HS65_LL_AOI21X2 U6945 ( .A(n3326), .B(n4062), .C(n4061), .Z(n4076) );
  HS65_LL_NAND2AX4 U6948 ( .A(n5474), .B(n2853), .Z(n5475) );
  HS65_LL_NAND4ABX3 U6949 ( .A(n4811), .B(n4810), .C(n4809), .D(n4808), .Z(
        n4815) );
  HS65_LL_NAND4ABX3 U6950 ( .A(n4231), .B(n4230), .C(n4229), .D(n4228), .Z(
        n4232) );
  HS65_LL_NAND3AX3 U6951 ( .A(n5381), .B(n2838), .C(n5380), .Z(n5382) );
  HS65_LL_NOR2AX3 U6952 ( .A(n3870), .B(n3869), .Z(n3871) );
  HS65_LL_NAND3AX3 U6954 ( .A(n4939), .B(n4938), .C(n4937), .Z(n4940) );
  HS65_LL_OAI12X3 U6956 ( .A(n2823), .B(n3907), .C(n3906), .Z(n3908) );
  HS65_LL_NOR2X2 U6959 ( .A(n4738), .B(n4430), .Z(n4455) );
  HS65_LL_AND3X4 U6960 ( .A(n5473), .B(n5472), .C(n5471), .Z(n2853) );
  HS65_LHS_XNOR2X6 U6964 ( .A(n3612), .B(n3611), .Z(n3613) );
  HS65_LH_NAND2AX4 U6966 ( .A(n5421), .B(n2859), .Z(n5047) );
  HS65_LL_NOR4ABX2 U6967 ( .A(n5169), .B(n5168), .C(n5167), .D(n5166), .Z(
        n5170) );
  HS65_LL_OAI21X2 U6969 ( .A(n3868), .B(n4812), .C(n3867), .Z(n3869) );
  HS65_LL_NAND4ABX3 U6970 ( .A(n4057), .B(n3699), .C(n3698), .D(n3697), .Z(
        n3700) );
  HS65_LL_NOR2AX3 U6971 ( .A(n3496), .B(n3495), .Z(n3868) );
  HS65_LH_NAND2X4 U6972 ( .A(n4461), .B(n4706), .Z(n4463) );
  HS65_LL_NAND3AX3 U6974 ( .A(n3900), .B(n3610), .C(n3609), .Z(n3611) );
  HS65_LH_CBI4I1X3 U6975 ( .A(n4796), .B(n4836), .C(n4795), .D(\lte_x_57/B[3] ), .Z(n4797) );
  HS65_LL_AOI21X2 U6977 ( .A(n4647), .B(n4646), .C(n4645), .Z(n4648) );
  HS65_LL_OR2X4 U6979 ( .A(n4171), .B(n3265), .Z(n2828) );
  HS65_LL_NOR2AX3 U6980 ( .A(n4576), .B(n4575), .Z(n4585) );
  HS65_LH_NAND2AX7 U6981 ( .A(n4559), .B(n4558), .Z(n4560) );
  HS65_LL_AOI22X1 U6982 ( .A(n5484), .B(n4851), .C(n4850), .D(n4849), .Z(n4852) );
  HS65_LH_AOI21X2 U6983 ( .A(n5484), .B(n4780), .C(n4312), .Z(n4319) );
  HS65_LH_AOI21X2 U6985 ( .A(n5517), .B(n4962), .C(n3914), .Z(n3934) );
  HS65_LL_NAND2X2 U6986 ( .A(n3208), .B(n4639), .Z(n3210) );
  HS65_LH_AOI21X2 U6990 ( .A(n4836), .B(n5479), .C(n3855), .Z(n3872) );
  HS65_LL_AO12X4 U6992 ( .A(n4536), .B(n3605), .C(n3244), .Z(n2851) );
  HS65_LH_AOI21X2 U6993 ( .A(n5505), .B(n4851), .C(n4223), .Z(n4229) );
  HS65_LH_OAI12X3 U6998 ( .A(n5359), .B(n5358), .C(n5357), .Z(n5383) );
  HS65_LL_NAND2AX4 U7000 ( .A(n3259), .B(n3263), .Z(n3265) );
  HS65_LHS_XOR2X3 U7002 ( .A(n4354), .B(n4353), .Z(n4355) );
  HS65_LH_AOI21X2 U7003 ( .A(n4121), .B(n4120), .C(n4738), .Z(n4122) );
  HS65_LLS_XOR2X3 U7005 ( .A(n3763), .B(n3762), .Z(n3764) );
  HS65_LLS_XNOR2X3 U7008 ( .A(n4772), .B(n4771), .Z(n4773) );
  HS65_LH_CBI4I1X3 U7011 ( .A(n5424), .B(n5376), .C(n5375), .D(n5374), .Z(
        n5378) );
  HS65_LH_OAI21X2 U7012 ( .A(n3944), .B(n3943), .C(n3942), .Z(n3945) );
  HS65_LH_NOR4ABX2 U7013 ( .A(n5295), .B(n5288), .C(n5287), .D(n5306), .Z(
        n5289) );
  HS65_LH_AND2X4 U7015 ( .A(n3974), .B(n3973), .Z(n2848) );
  HS65_LH_AOI21X2 U7020 ( .A(n4323), .B(n4322), .C(n4321), .Z(n4329) );
  HS65_LH_AOI31X2 U7023 ( .A(n4116), .B(n4115), .C(n4114), .D(n4440), .Z(n3229) );
  HS65_LL_OA12X9 U7024 ( .A(n3760), .B(n3257), .C(n3256), .Z(n2823) );
  HS65_LH_OAI21X2 U7029 ( .A(n5360), .B(n5355), .C(n5361), .Z(n5032) );
  HS65_LH_NAND2AX4 U7030 ( .A(n4969), .B(n4968), .Z(n4981) );
  HS65_LH_NAND3AX3 U7032 ( .A(n5407), .B(n5337), .C(n5037), .Z(n5038) );
  HS65_LL_AOI12X2 U7033 ( .A(n5130), .B(n5129), .C(n5128), .Z(n5137) );
  HS65_LL_NOR2AX6 U7034 ( .A(n2994), .B(n2789), .Z(n4842) );
  HS65_LL_AOI22X1 U7035 ( .A(n3239), .B(n7679), .C(n7681), .D(
        \u_DataPath/u_execute/resAdd1_i [31]), .Z(n8128) );
  HS65_LH_AOI21X2 U7036 ( .A(n5151), .B(n5150), .C(n5149), .Z(n5152) );
  HS65_LL_NAND2AX4 U7038 ( .A(n3464), .B(n3463), .Z(n3835) );
  HS65_LHS_XNOR2X6 U7041 ( .A(n9041), .B(n5670), .Z(\u_DataPath/toPC2_i [31])
         );
  HS65_LH_NAND2X2 U7042 ( .A(n5114), .B(n5081), .Z(n5087) );
  HS65_LL_IVX2 U7043 ( .A(n4170), .Z(n4082) );
  HS65_LL_MUX21I1X3 U7045 ( .D0(n4571), .D1(n5502), .S0(n5092), .Z(n4146) );
  HS65_LH_NAND2AX7 U7046 ( .A(n4903), .B(n4930), .Z(n4932) );
  HS65_LL_AOI12X2 U7047 ( .A(n5262), .B(n5261), .C(n5260), .Z(n5271) );
  HS65_LL_NAND2AX4 U7048 ( .A(n3647), .B(n3646), .Z(n3865) );
  HS65_LL_NAND2X2 U7050 ( .A(n3000), .B(n4864), .Z(n3003) );
  HS65_LL_AOI22X1 U7052 ( .A(n8313), .B(n9434), .C(n7694), .D(
        \u_DataPath/u_execute/link_value_i [30]), .Z(n8287) );
  HS65_LL_AO22X4 U7053 ( .A(\lte_x_57/B[30] ), .B(n7680), .C(n7682), .D(
        \u_DataPath/u_execute/resAdd1_i [30]), .Z(
        \u_DataPath/jump_address_i [30]) );
  HS65_LL_OAI12X3 U7054 ( .A(n5245), .B(n4426), .C(n5244), .Z(n4369) );
  HS65_LH_NAND3X5 U7055 ( .A(n3734), .B(n3733), .C(n3732), .Z(n3801) );
  HS65_LH_NOR2X2 U7056 ( .A(n3888), .B(n5083), .Z(n5086) );
  HS65_LH_NOR2X2 U7057 ( .A(n3954), .B(n3972), .Z(n3946) );
  HS65_LH_NOR2X2 U7058 ( .A(n5107), .B(n5080), .Z(n5081) );
  HS65_LH_NAND2AX7 U7060 ( .A(n4190), .B(n3462), .Z(n3464) );
  HS65_LL_OAI12X2 U7061 ( .A(n4272), .B(n5080), .C(n5227), .Z(n5230) );
  HS65_LL_NOR2X2 U7062 ( .A(n3633), .B(n5245), .Z(n5065) );
  HS65_LH_AOI21X2 U7063 ( .A(n3961), .B(n5371), .C(n5362), .Z(n3965) );
  HS65_LH_OAI21X2 U7064 ( .A(n5232), .B(n3888), .C(n3886), .Z(n5118) );
  HS65_LH_IVX9 U7065 ( .A(n3593), .Z(n4440) );
  HS65_LH_NAND2X5 U7066 ( .A(n4189), .B(n5211), .Z(n5347) );
  HS65_LH_IVX9 U7068 ( .A(n4849), .Z(n4624) );
  HS65_LH_CBI4I6X2 U7069 ( .A(n4922), .B(n4921), .C(n4920), .D(n4919), .Z(
        n4924) );
  HS65_LL_NAND3X2 U7070 ( .A(n4920), .B(n5005), .C(n5433), .Z(n4914) );
  HS65_LH_OAI21X2 U7073 ( .A(n3633), .B(n5126), .C(n5125), .Z(n5130) );
  HS65_LH_OAI12X3 U7074 ( .A(n4768), .B(n4765), .C(n4767), .Z(n2996) );
  HS65_LH_AOI21X2 U7078 ( .A(n4796), .B(\sub_x_51/A[8] ), .C(n3859), .Z(n3864)
         );
  HS65_LH_CNIVX3 U7081 ( .A(n5237), .Z(n3966) );
  HS65_LH_AOI21X2 U7082 ( .A(n3994), .B(n5003), .C(n5002), .Z(n3995) );
  HS65_LH_NAND2AX7 U7083 ( .A(n2854), .B(n4118), .Z(n4849) );
  HS65_LL_NOR2AX3 U7087 ( .A(n3248), .B(n3536), .Z(n3267) );
  HS65_LL_NAND2AX4 U7088 ( .A(n3389), .B(n3388), .Z(n3390) );
  HS65_LL_AOI22X1 U7090 ( .A(\lte_x_57/B[29] ), .B(n7680), .C(n7682), .D(
        \u_DataPath/u_execute/resAdd1_i [29]), .Z(n8132) );
  HS65_LL_NOR2X3 U7092 ( .A(n3713), .B(n3712), .Z(n4070) );
  HS65_LH_NAND2AX7 U7093 ( .A(n3329), .B(n3328), .Z(n3330) );
  HS65_LH_NAND2X4 U7096 ( .A(n4374), .B(n3248), .Z(n4380) );
  HS65_LL_OAI12X3 U7097 ( .A(n4277), .B(n4046), .C(n4048), .Z(n4260) );
  HS65_LL_AOI21X2 U7098 ( .A(\lte_x_57/B[3] ), .B(n3742), .C(n3476), .Z(n3477)
         );
  HS65_LH_AOI21X2 U7100 ( .A(n5362), .B(n5361), .C(n5360), .Z(n5370) );
  HS65_LL_NOR2AX3 U7101 ( .A(n3246), .B(n3353), .Z(n3273) );
  HS65_LH_NOR2X5 U7103 ( .A(n5208), .B(n3948), .Z(n5341) );
  HS65_LL_NAND2AX4 U7105 ( .A(n5186), .B(\sub_x_51/A[16] ), .Z(n5027) );
  HS65_LH_NAND2X5 U7106 ( .A(n5208), .B(n3948), .Z(n5412) );
  HS65_LH_NOR2X5 U7108 ( .A(n3993), .B(n5246), .Z(n5002) );
  HS65_LH_NAND2X5 U7109 ( .A(n4283), .B(n5201), .Z(n5337) );
  HS65_LHS_XOR2X3 U7111 ( .A(n5529), .B(n5067), .Z(n4983) );
  HS65_LH_CNIVX3 U7112 ( .A(n3765), .Z(n3766) );
  HS65_LL_NOR2AX3 U7115 ( .A(n4778), .B(n3729), .Z(n3388) );
  HS65_LL_NAND3X2 U7116 ( .A(n3569), .B(n3458), .C(n3583), .Z(n4570) );
  HS65_LL_AOI22X1 U7118 ( .A(\sub_x_51/A[13] ), .B(n3826), .C(n2793), .D(n5498), .Z(n3401) );
  HS65_LH_AO22X9 U7121 ( .A(\lte_x_57/B[28] ), .B(n7680), .C(n7682), .D(
        \u_DataPath/u_execute/resAdd1_i [28]), .Z(
        \u_DataPath/jump_address_i [28]) );
  HS65_LH_OAI12X3 U7122 ( .A(n3886), .B(n5396), .C(n5115), .Z(n3080) );
  HS65_LHS_XNOR2X6 U7123 ( .A(n2824), .B(n5064), .Z(n4984) );
  HS65_LHS_XNOR2X3 U7124 ( .A(n2780), .B(n5487), .Z(n5488) );
  HS65_LL_NOR2AX3 U7126 ( .A(n3917), .B(n2855), .Z(n3320) );
  HS65_LL_NOR2X2 U7129 ( .A(n5366), .B(n5360), .Z(n4884) );
  HS65_LH_CNIVX3 U7136 ( .A(n3729), .Z(n3734) );
  HS65_LL_NAND2X5 U7138 ( .A(n3012), .B(n3011), .Z(n5077) );
  HS65_LL_NOR2X3 U7139 ( .A(\lte_x_57/B[6] ), .B(n5089), .Z(n4818) );
  HS65_LHS_XNOR2X6 U7140 ( .A(\lte_x_57/B[6] ), .B(n5089), .Z(n4943) );
  HS65_LH_OR2X4 U7141 ( .A(n2780), .B(n5508), .Z(n5489) );
  HS65_LL_CBI4I1X3 U7142 ( .A(n5507), .B(n5508), .C(n5506), .D(n2780), .Z(
        n5514) );
  HS65_LL_NAND2X2 U7143 ( .A(\lte_x_57/B[2] ), .B(n5092), .Z(n4802) );
  HS65_LL_OAI12X2 U7145 ( .A(n5298), .B(n5304), .C(n5284), .Z(n4919) );
  HS65_LL_AOI22X3 U7146 ( .A(n3940), .B(n3826), .C(n2780), .D(n5498), .Z(n4468) );
  HS65_LL_NOR2AX3 U7149 ( .A(n3742), .B(n4871), .Z(n3228) );
  HS65_LL_NOR2X3 U7150 ( .A(\lte_x_57/B[15] ), .B(n2788), .Z(n5396) );
  HS65_LH_IVX9 U7151 ( .A(n2969), .Z(n3777) );
  HS65_LH_IVX9 U7156 ( .A(n5186), .Z(n2795) );
  HS65_LH_OR2X4 U7158 ( .A(n3239), .B(n7317), .Z(n4636) );
  HS65_LL_NAND2AX7 U7160 ( .A(n2846), .B(n3134), .Z(n5187) );
  HS65_LL_MUX21I1X3 U7161 ( .D0(n7676), .D1(n8730), .S0(
        \u_DataPath/cw_to_ex_i [14]), .Z(n5067) );
  HS65_LH_NOR2X5 U7162 ( .A(n4032), .B(n5079), .Z(n5424) );
  HS65_LH_AO22X9 U7163 ( .A(\sub_x_51/A[22] ), .B(n7680), .C(n7682), .D(
        \u_DataPath/u_execute/resAdd1_i [22]), .Z(
        \u_DataPath/jump_address_i [22]) );
  HS65_LH_OAI21X3 U7165 ( .A(n8288), .B(n8317), .C(n7696), .Z(
        \u_DataPath/from_mem_data_out_i [30]) );
  HS65_LH_AO222X4 U7166 ( .A(n7706), .B(n8969), .C(n7685), .D(n9281), .E(n7691), .F(n9406), .Z(addr_to_iram_29) );
  HS65_LH_IVX9 U7168 ( .A(n5392), .Z(n3079) );
  HS65_LH_OAI21X3 U7169 ( .A(n8318), .B(n8317), .C(n7697), .Z(
        \u_DataPath/from_mem_data_out_i [29]) );
  HS65_LH_OAI21X3 U7170 ( .A(n8294), .B(n8317), .C(n7696), .Z(
        \u_DataPath/from_mem_data_out_i [28]) );
  HS65_LH_OAI21X3 U7171 ( .A(n8216), .B(n8317), .C(n7697), .Z(
        \u_DataPath/from_mem_data_out_i [27]) );
  HS65_LH_AO22X9 U7173 ( .A(\lte_x_57/B[3] ), .B(n7680), .C(n7682), .D(
        \u_DataPath/u_execute/resAdd1_i [3]), .Z(
        \u_DataPath/jump_address_i [3]) );
  HS65_LL_CBI4I1X3 U7174 ( .A(n5507), .B(n3949), .C(n5506), .D(\sub_x_51/A[5] ), .Z(n3727) );
  HS65_LH_AO22X9 U7175 ( .A(\lte_x_57/B[10] ), .B(n7680), .C(n7682), .D(
        \u_DataPath/u_execute/resAdd1_i [10]), .Z(
        \u_DataPath/jump_address_i [10]) );
  HS65_LH_AO22X9 U7176 ( .A(n7680), .B(\u_DataPath/u_execute/A_inALU_i[26] ), 
        .C(n7682), .D(\u_DataPath/u_execute/resAdd1_i [26]), .Z(
        \u_DataPath/jump_address_i [26]) );
  HS65_LH_NOR2AX3 U7177 ( .A(\sub_x_51/A[5] ), .B(n2830), .Z(n3729) );
  HS65_LH_AO22X9 U7178 ( .A(\sub_x_51/A[16] ), .B(n7680), .C(n7682), .D(
        \u_DataPath/u_execute/resAdd1_i [16]), .Z(
        \u_DataPath/jump_address_i [16]) );
  HS65_LL_NOR3AX2 U7181 ( .A(n8989), .B(n8800), .C(n7981), .Z(n7983) );
  HS65_LH_OAI21X3 U7184 ( .A(n8311), .B(n8317), .C(n7697), .Z(
        \u_DataPath/from_mem_data_out_i [31]) );
  HS65_LHS_XOR2X3 U7185 ( .A(n3239), .B(n7321), .Z(n5163) );
  HS65_LH_NAND4ABX3 U7187 ( .A(n8752), .B(n8686), .C(n9367), .D(n8362), .Z(
        \u_DataPath/cw_exmem_i [10]) );
  HS65_LH_AO22X9 U7188 ( .A(\lte_x_57/B[14] ), .B(n7680), .C(n7682), .D(
        \u_DataPath/u_execute/resAdd1_i [14]), .Z(
        \u_DataPath/jump_address_i [14]) );
  HS65_LH_OR2X4 U7190 ( .A(n7321), .B(n5148), .Z(n5151) );
  HS65_LH_OAI21X3 U7191 ( .A(n8202), .B(n8317), .C(n7697), .Z(
        \u_DataPath/from_mem_data_out_i [21]) );
  HS65_LH_OAI21X3 U7192 ( .A(n8250), .B(n8317), .C(n7697), .Z(
        \u_DataPath/from_mem_data_out_i [26]) );
  HS65_LH_OAI21X3 U7193 ( .A(n8284), .B(n8317), .C(n7696), .Z(
        \u_DataPath/from_mem_data_out_i [22]) );
  HS65_LH_OAI21X3 U7194 ( .A(n8187), .B(n8317), .C(n7696), .Z(
        \u_DataPath/from_mem_data_out_i [16]) );
  HS65_LH_OAI21X3 U7195 ( .A(n8291), .B(n8317), .C(n7696), .Z(
        \u_DataPath/from_mem_data_out_i [20]) );
  HS65_LH_OAI21X3 U7196 ( .A(n8193), .B(n8317), .C(n7697), .Z(
        \u_DataPath/from_mem_data_out_i [17]) );
  HS65_LL_NAND3AX3 U7197 ( .A(n3060), .B(n3059), .C(n9543), .Z(n3061) );
  HS65_LH_OAI21X3 U7198 ( .A(n8242), .B(n8317), .C(n7697), .Z(
        \u_DataPath/from_mem_data_out_i [18]) );
  HS65_LHS_XOR2X3 U7199 ( .A(n9002), .B(n5768), .Z(
        \u_DataPath/u_execute/resAdd1_i [27]) );
  HS65_LH_NAND2X5 U7200 ( .A(n3950), .B(n3949), .Z(n5349) );
  HS65_LH_OAI21X3 U7201 ( .A(n8220), .B(n8317), .C(n7697), .Z(
        \u_DataPath/from_mem_data_out_i [23]) );
  HS65_LH_OAI21X3 U7202 ( .A(n8197), .B(n8317), .C(n7697), .Z(
        \u_DataPath/from_mem_data_out_i [19]) );
  HS65_LH_OAI21X3 U7203 ( .A(n8260), .B(n8317), .C(n7697), .Z(
        \u_DataPath/from_mem_data_out_i [25]) );
  HS65_LH_AO22X9 U7204 ( .A(n3039), .B(n7680), .C(n7682), .D(
        \u_DataPath/u_execute/resAdd1_i [9]), .Z(
        \u_DataPath/jump_address_i [9]) );
  HS65_LH_OAI21X3 U7205 ( .A(n8231), .B(n8317), .C(n7697), .Z(
        \u_DataPath/from_mem_data_out_i [24]) );
  HS65_LL_OAI22X1 U7206 ( .A(n6861), .B(n7896), .C(n7716), .D(n8067), .Z(
        \u_DataPath/data_read_ex_2_i [19]) );
  HS65_LL_OAI22X1 U7207 ( .A(n6861), .B(n7732), .C(n7716), .D(n8062), .Z(
        \u_DataPath/data_read_ex_2_i [10]) );
  HS65_LH_NAND2X4 U7208 ( .A(Data_out_fromRAM[15]), .B(n8300), .Z(n8301) );
  HS65_LL_OR2X4 U7209 ( .A(n3940), .B(n2968), .Z(n5094) );
  HS65_LH_NAND2X4 U7210 ( .A(Data_out_fromRAM[13]), .B(n8300), .Z(n8167) );
  HS65_LH_NAND2X4 U7211 ( .A(Data_out_fromRAM[14]), .B(n8300), .Z(n8253) );
  HS65_LL_MUX21I1X6 U7212 ( .D0(n8450), .D1(n8730), .S0(
        \u_DataPath/cw_to_ex_i [14]), .Z(n5312) );
  HS65_LH_AO22X9 U7213 ( .A(n5192), .B(n7680), .C(n7682), .D(
        \u_DataPath/u_execute/resAdd1_i [24]), .Z(
        \u_DataPath/jump_address_i [24]) );
  HS65_LH_AO22X9 U7214 ( .A(\add_x_50/A[19] ), .B(n7680), .C(n7682), .D(
        \u_DataPath/u_execute/resAdd1_i [19]), .Z(
        \u_DataPath/jump_address_i [19]) );
  HS65_LH_NAND2X4 U7215 ( .A(Data_out_fromRAM[12]), .B(n8300), .Z(n8239) );
  HS65_LH_AO222X4 U7216 ( .A(n7706), .B(n8968), .C(n7691), .D(n8619), .E(n9022), .F(n7685), .Z(addr_to_iram_28) );
  HS65_LH_NAND2X4 U7217 ( .A(Data_out_fromRAM[11]), .B(n8300), .Z(n8215) );
  HS65_LH_NAND2X4 U7218 ( .A(Data_out_fromRAM[10]), .B(n8300), .Z(n8234) );
  HS65_LH_NAND2X4 U7219 ( .A(Data_out_fromRAM[9]), .B(n8300), .Z(n8259) );
  HS65_LL_AO112X4 U7220 ( .A(n8719), .B(n2712), .C(n3167), .D(n3166), .Z(n2825) );
  HS65_LH_NAND2X4 U7221 ( .A(Data_out_fromRAM[8]), .B(n8300), .Z(n8230) );
  HS65_LLS_XOR2X3 U7222 ( .A(addr_to_iram_29), .B(n7457), .Z(
        \u_DataPath/pc_4_i [31]) );
  HS65_LL_AO112X4 U7224 ( .A(n8691), .B(n2710), .C(n3172), .D(n3171), .Z(n2824) );
  HS65_LH_OR2X9 U7226 ( .A(n3006), .B(n3005), .Z(n4203) );
  HS65_LH_AO22X9 U7229 ( .A(n7680), .B(\lte_x_57/B[7] ), .C(n7682), .D(
        \u_DataPath/u_execute/resAdd1_i [7]), .Z(
        \u_DataPath/jump_address_i [7]) );
  HS65_LH_AOI22X3 U7230 ( .A(\sub_x_51/A[5] ), .B(n7679), .C(n7681), .D(
        \u_DataPath/u_execute/resAdd1_i [5]), .Z(n8177) );
  HS65_LH_AO222X4 U7231 ( .A(n7706), .B(n8967), .C(n7691), .D(n9453), .E(n9280), .F(n7685), .Z(addr_to_iram_27) );
  HS65_LHS_XNOR2X6 U7232 ( .A(n7407), .B(n7456), .Z(\u_DataPath/pc_4_i [30])
         );
  HS65_LH_OR3X9 U7233 ( .A(\u_DataPath/cw_exmem_i [3]), .B(n7948), .C(
        \u_DataPath/u_idexreg/N13 ), .Z(\u_DataPath/u_idexreg/N10 ) );
  HS65_LL_OR2X4 U7234 ( .A(n2977), .B(n2772), .Z(n2831) );
  HS65_LL_OAI12X3 U7236 ( .A(n3181), .B(n9282), .C(n2929), .Z(\lte_x_57/B[7] )
         );
  HS65_LH_AOI211X3 U7237 ( .A(n8023), .B(n8603), .C(\u_DataPath/u_idexreg/N15 ), .D(\u_DataPath/u_idexreg/N16 ), .Z(n7960) );
  HS65_LH_NOR3X4 U7238 ( .A(n7963), .B(n8990), .C(n7962), .Z(n7989) );
  HS65_LL_OA12X4 U7239 ( .A(n9288), .B(n3181), .C(n3111), .Z(n2806) );
  HS65_LL_OAI12X3 U7240 ( .A(n9128), .B(n5787), .C(n9031), .Z(n5920) );
  HS65_LHS_XOR2X3 U7242 ( .A(n9008), .B(n5787), .Z(
        \u_DataPath/u_execute/resAdd1_i [25]) );
  HS65_LH_OR2X9 U7243 ( .A(n8658), .B(n3181), .Z(n2826) );
  HS65_LL_OR2X4 U7244 ( .A(n8629), .B(n3181), .Z(n3041) );
  HS65_LH_IVX9 U7245 ( .A(n9538), .Z(n2968) );
  HS65_LH_AOI22X3 U7248 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][30] ), .B(n8950), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][30] ), .D(
        n8855), .Z(n6570) );
  HS65_LH_AOI22X3 U7249 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][3] ), .B(n9248), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][3] ), .D(
        n9240), .Z(n6449) );
  HS65_LL_NAND3AX3 U7250 ( .A(n2937), .B(n2936), .C(n2935), .Z(n3950) );
  HS65_LHS_XNOR2X6 U7251 ( .A(n8908), .B(n2807), .Z(
        \u_DataPath/u_execute/resAdd1_i [14]) );
  HS65_LH_OA112X18 U7252 ( .A(n8642), .B(n3149), .C(n3238), .D(n3237), .Z(
        n3239) );
  HS65_LH_AO222X4 U7253 ( .A(n7706), .B(n9020), .C(n7691), .D(n8618), .E(n8877), .F(n7685), .Z(addr_to_iram_26) );
  HS65_LH_AO222X4 U7254 ( .A(n7706), .B(n8966), .C(n7690), .D(
        \u_DataPath/jump_address_i [17]), .E(n8837), .F(n7686), .Z(
        addr_to_iram_15) );
  HS65_LH_OA12X9 U7255 ( .A(n8671), .B(n3149), .C(n3135), .Z(n3136) );
  HS65_LL_NOR4ABX2 U7256 ( .A(n8740), .B(n8186), .C(n9350), .D(n9286), .Z(
        n8166) );
  HS65_LL_NOR2X2 U7257 ( .A(n3218), .B(n8369), .Z(n2957) );
  HS65_LHS_XNOR2X3 U7258 ( .A(n9223), .B(n6758), .Z(
        \u_DataPath/u_execute/link_value_i [24]) );
  HS65_LHS_XNOR2X6 U7260 ( .A(n9093), .B(n5880), .Z(
        \u_DataPath/u_execute/resAdd1_i [19]) );
  HS65_LHS_XOR2X6 U7261 ( .A(n7606), .B(n7605), .Z(\u_DataPath/pc_4_i [29]) );
  HS65_LH_AOI12X2 U7262 ( .A(n9390), .B(n5678), .C(n9272), .Z(n5579) );
  HS65_LH_BFX9 U7263 ( .A(n8368), .Z(n7718) );
  HS65_LH_AOI22X3 U7267 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][20] ), .B(n9255), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][20] ), .D(
        n9195), .Z(n6585) );
  HS65_LH_AOI22X3 U7268 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][1] ), .B(n9472), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][1] ), .D(
        n9468), .Z(n6240) );
  HS65_LH_BFX9 U7269 ( .A(n8320), .Z(n7698) );
  HS65_LH_BFX9 U7271 ( .A(n8320), .Z(n7700) );
  HS65_LHS_XOR2X3 U7272 ( .A(n9292), .B(n7627), .Z(
        \u_DataPath/u_execute/link_value_i [23]) );
  HS65_LL_AOI12X6 U7273 ( .A(n9318), .B(n2820), .C(n8036), .Z(n8526) );
  HS65_LH_AND2X4 U7274 ( .A(n8806), .B(n8513), .Z(n7949) );
  HS65_LH_OAI12X3 U7275 ( .A(n9394), .B(n5587), .C(n9393), .Z(n5678) );
  HS65_LL_NAND3X2 U7276 ( .A(n8901), .B(n7994), .C(n8513), .Z(n7998) );
  HS65_LH_AO222X4 U7277 ( .A(n7706), .B(n8964), .C(n7691), .D(n9328), .E(n9450), .F(n7685), .Z(addr_to_iram_25) );
  HS65_LH_AO222X4 U7278 ( .A(n7706), .B(n8883), .C(n7690), .D(
        \u_DataPath/jump_address_i [23]), .E(n9323), .F(n7685), .Z(
        addr_to_iram_21) );
  HS65_LH_AO222X4 U7279 ( .A(n7706), .B(n8965), .C(n7690), .D(n9379), .E(n9320), .F(n7685), .Z(addr_to_iram_19) );
  HS65_LHS_XNOR2X6 U7280 ( .A(n7388), .B(n7387), .Z(\u_DataPath/pc_4_i [17])
         );
  HS65_LH_BFX9 U7281 ( .A(n8320), .Z(n7699) );
  HS65_LL_NAND2AX4 U7282 ( .A(n2965), .B(n2964), .Z(n2967) );
  HS65_LH_OAI12X3 U7283 ( .A(n9277), .B(n5790), .C(n9347), .Z(n2807) );
  HS65_LH_OAI12X3 U7284 ( .A(n9277), .B(n5790), .C(n9347), .Z(n5872) );
  HS65_LH_IVX9 U7285 ( .A(n5813), .Z(n5790) );
  HS65_LH_AOI12X2 U7287 ( .A(n9424), .B(n5682), .C(n9274), .Z(n5621) );
  HS65_LH_AOI12X2 U7288 ( .A(n9397), .B(n5682), .C(n5634), .Z(n5636) );
  HS65_LHS_XOR2X6 U7289 ( .A(n7472), .B(n7471), .Z(\u_DataPath/pc_4_i [21]) );
  HS65_LH_AOI12X2 U7291 ( .A(n9386), .B(n5605), .C(n9417), .Z(n5607) );
  HS65_LH_AOI12X2 U7292 ( .A(n9341), .B(n5686), .C(n9423), .Z(n5598) );
  HS65_LHS_XOR2X3 U7295 ( .A(n7474), .B(n7473), .Z(\u_DataPath/pc_4_i [27]) );
  HS65_LH_NOR2X3 U7299 ( .A(n8703), .B(n8071), .Z(n8468) );
  HS65_LH_NOR2X5 U7301 ( .A(n3030), .B(n8393), .Z(n3031) );
  HS65_LL_MUXI21X2 U7302 ( .D0(n9338), .D1(n8452), .S0(n3090), .Z(n3982) );
  HS65_LHS_XOR2X3 U7303 ( .A(n9295), .B(n9075), .Z(
        \u_DataPath/u_execute/link_value_i [21]) );
  HS65_LH_BFX9 U7304 ( .A(n8472), .Z(n7742) );
  HS65_LH_NAND2X4 U7306 ( .A(n8764), .B(n3107), .Z(n3024) );
  HS65_LHS_XNOR2X6 U7309 ( .A(n7383), .B(n7470), .Z(\u_DataPath/pc_4_i [20])
         );
  HS65_LHS_XNOR2X3 U7310 ( .A(n7378), .B(n7389), .Z(\u_DataPath/pc_4_i [26])
         );
  HS65_LH_BFX9 U7311 ( .A(n8480), .Z(n7787) );
  HS65_LH_OAI12X3 U7312 ( .A(n8971), .B(n5699), .C(n9147), .Z(n5701) );
  HS65_LH_BFX9 U7313 ( .A(n7708), .Z(n7707) );
  HS65_LHS_XNOR2X6 U7314 ( .A(n7373), .B(n7372), .Z(\u_DataPath/pc_4_i [19])
         );
  HS65_LHS_XNOR2X6 U7315 ( .A(n7363), .B(n7362), .Z(\u_DataPath/pc_4_i [13])
         );
  HS65_LHS_XNOR2X6 U7316 ( .A(n7359), .B(n7358), .Z(\u_DataPath/pc_4_i [15])
         );
  HS65_LH_NOR2X5 U7317 ( .A(\u_DataPath/dataOut_exe_i [25]), .B(n3980), .Z(
        n8444) );
  HS65_LL_OAI12X18 U7318 ( .A(n8720), .B(n8012), .C(n1885), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N132 ) );
  HS65_LL_OAI12X12 U7319 ( .A(n8005), .B(n3532), .C(n1885), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N144 ) );
  HS65_LL_OAI12X12 U7321 ( .A(n8004), .B(n8689), .C(n1885), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N153 ) );
  HS65_LH_BFX9 U7322 ( .A(n8489), .Z(n7850) );
  HS65_LHS_XNOR2X6 U7323 ( .A(n9214), .B(n9013), .Z(
        \u_DataPath/u_execute/link_value_i [7]) );
  HS65_LL_OAI12X18 U7324 ( .A(n8009), .B(n8012), .C(n1885), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N137 ) );
  HS65_LL_OAI12X18 U7326 ( .A(n3532), .B(n8012), .C(n1885), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N136 ) );
  HS65_LHS_XOR2X6 U7327 ( .A(n7463), .B(n7462), .Z(\u_DataPath/pc_4_i [11]) );
  HS65_LHS_XOR2X6 U7328 ( .A(n7466), .B(n7465), .Z(\u_DataPath/pc_4_i [9]) );
  HS65_LH_BFX9 U7329 ( .A(n8462), .Z(n7721) );
  HS65_LL_OAI12X18 U7330 ( .A(n8726), .B(n8012), .C(n1885), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N133 ) );
  HS65_LH_AND3X9 U7331 ( .A(n2990), .B(n2989), .C(n9103), .Z(n7670) );
  HS65_LH_BFX9 U7332 ( .A(n8485), .Z(n7822) );
  HS65_LHS_XOR2X3 U7333 ( .A(n7451), .B(n7450), .Z(\u_DataPath/pc_4_i [25]) );
  HS65_LL_OAI12X12 U7334 ( .A(n8005), .B(n7644), .C(n1885), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N145 ) );
  HS65_LL_OAI12X18 U7335 ( .A(n2720), .B(n8012), .C(n1885), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N135 ) );
  HS65_LL_OAI12X12 U7337 ( .A(n8005), .B(n8726), .C(n1885), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N141 ) );
  HS65_LH_BFX9 U7338 ( .A(n8483), .Z(n7808) );
  HS65_LL_OAI12X12 U7339 ( .A(n8005), .B(n8720), .C(n1885), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N140 ) );
  HS65_LH_BFX9 U7341 ( .A(n8495), .Z(n7892) );
  HS65_LH_BFX9 U7342 ( .A(n8499), .Z(n7913) );
  HS65_LH_BFX9 U7343 ( .A(n8491), .Z(n7864) );
  HS65_LH_BFX9 U7344 ( .A(n8493), .Z(n7878) );
  HS65_LH_BFX9 U7345 ( .A(n8481), .Z(n7794) );
  HS65_LH_BFX9 U7346 ( .A(n8476), .Z(n7759) );
  HS65_LH_BFX9 U7347 ( .A(n8497), .Z(n7906) );
  HS65_LH_BFX9 U7348 ( .A(n6278), .Z(n7000) );
  HS65_LH_BFX9 U7349 ( .A(n7588), .Z(n7508) );
  HS65_LH_BFX9 U7350 ( .A(n8490), .Z(n7857) );
  HS65_LH_BFX9 U7351 ( .A(n6132), .Z(n7502) );
  HS65_LH_NAND2X4 U7352 ( .A(opcode_i[3]), .B(n7393), .Z(n7966) );
  HS65_LH_BFX9 U7353 ( .A(n8486), .Z(n7829) );
  HS65_LL_OAI12X3 U7354 ( .A(n3184), .B(n8375), .C(n2976), .Z(n2978) );
  HS65_LH_BFX9 U7355 ( .A(n6245), .Z(n6992) );
  HS65_LL_NOR2AX3 U7356 ( .A(n7674), .B(n9066), .Z(n2990) );
  HS65_LH_OAI21X3 U7357 ( .A(opcode_i[0]), .B(n7608), .C(n7409), .Z(n7334) );
  HS65_LH_BFX9 U7358 ( .A(n8488), .Z(n7843) );
  HS65_LH_BFX9 U7359 ( .A(n8492), .Z(n7871) );
  HS65_LH_IVX9 U7360 ( .A(n5572), .Z(n2799) );
  HS65_LH_BFX9 U7361 ( .A(n8477), .Z(n7766) );
  HS65_LH_BFX9 U7362 ( .A(n6120), .Z(n7577) );
  HS65_LH_BFX9 U7363 ( .A(n6272), .Z(n6993) );
  HS65_LH_BFX9 U7364 ( .A(n8487), .Z(n7836) );
  HS65_LH_BFX9 U7365 ( .A(n6119), .Z(n7578) );
  HS65_LHS_XNOR2X6 U7366 ( .A(n7339), .B(n7338), .Z(\u_DataPath/pc_4_i [7]) );
  HS65_LH_BFX9 U7367 ( .A(n6345), .Z(n6999) );
  HS65_LH_BFX9 U7368 ( .A(n5980), .Z(n7560) );
  HS65_LH_BFX9 U7369 ( .A(n8470), .Z(n7728) );
  HS65_LL_AND2X4 U7370 ( .A(n9362), .B(n2989), .Z(n2918) );
  HS65_LH_BFX9 U7371 ( .A(n6113), .Z(n7518) );
  HS65_LH_BFX9 U7372 ( .A(n6128), .Z(n7585) );
  HS65_LH_BFX9 U7373 ( .A(n5981), .Z(n7595) );
  HS65_LH_BFX9 U7374 ( .A(n8494), .Z(n7885) );
  HS65_LH_BFX9 U7375 ( .A(n8496), .Z(n7899) );
  HS65_LH_BFX9 U7376 ( .A(n6498), .Z(n6973) );
  HS65_LH_BFX9 U7377 ( .A(n8473), .Z(n7749) );
  HS65_LH_BFX9 U7378 ( .A(n6129), .Z(n7580) );
  HS65_LH_BFX9 U7379 ( .A(n8478), .Z(n7773) );
  HS65_LH_BFX9 U7380 ( .A(n8479), .Z(n7780) );
  HS65_LH_BFX9 U7381 ( .A(n8471), .Z(n7735) );
  HS65_LH_BFX9 U7382 ( .A(n6112), .Z(n7515) );
  HS65_LH_BFX9 U7383 ( .A(n8484), .Z(n7815) );
  HS65_LHS_XOR2X3 U7384 ( .A(n7617), .B(n7616), .Z(
        \u_DataPath/u_execute/link_value_i [6]) );
  HS65_LH_BFX9 U7385 ( .A(n8482), .Z(n7801) );
  HS65_LH_BFX9 U7386 ( .A(n7692), .Z(n7694) );
  HS65_LH_BFX9 U7387 ( .A(n7692), .Z(n7695) );
  HS65_LH_BFX9 U7388 ( .A(n6530), .Z(n6918) );
  HS65_LH_BFX9 U7389 ( .A(n6131), .Z(n7503) );
  HS65_LL_NOR2X5 U7390 ( .A(n5961), .B(n5939), .Z(n6017) );
  HS65_LL_NOR2X5 U7391 ( .A(n6175), .B(n6188), .Z(n6264) );
  HS65_LHS_XOR2X6 U7392 ( .A(n9169), .B(n9316), .Z(n6480) );
  HS65_LH_BFX9 U7393 ( .A(n6528), .Z(n6917) );
  HS65_LL_NOR2X5 U7394 ( .A(n6175), .B(n6182), .Z(n6529) );
  HS65_LH_BFX9 U7395 ( .A(n6347), .Z(n6895) );
  HS65_LL_NOR2X5 U7396 ( .A(n5959), .B(n5939), .Z(n6016) );
  HS65_LH_OR2X9 U7397 ( .A(\u_DataPath/cw_to_ex_i [1]), .B(n7315), .Z(n4305)
         );
  HS65_LH_BFX9 U7398 ( .A(n6121), .Z(n7501) );
  HS65_LL_NOR2X5 U7399 ( .A(n5958), .B(n5939), .Z(n6014) );
  HS65_LL_NOR2X5 U7400 ( .A(n5963), .B(n5939), .Z(n6015) );
  HS65_LH_BFX9 U7401 ( .A(n6340), .Z(n6890) );
  HS65_LL_NOR2X5 U7402 ( .A(n2870), .B(n2869), .Z(n2889) );
  HS65_LH_BFX9 U7403 ( .A(n7684), .Z(n7686) );
  HS65_LH_BFX9 U7404 ( .A(n7684), .Z(n7685) );
  HS65_LH_BFX9 U7405 ( .A(n3465), .Z(n5517) );
  HS65_LH_BFX9 U7406 ( .A(n6114), .Z(n7517) );
  HS65_LH_BFX9 U7407 ( .A(n7684), .Z(n7687) );
  HS65_LH_AND3X4 U7408 ( .A(\u_DataPath/cw_tomem_i [5]), .B(n3438), .C(n7352), 
        .Z(n3561) );
  HS65_LH_BFX9 U7409 ( .A(n6130), .Z(n7579) );
  HS65_LH_NOR2X3 U7410 ( .A(\u_DataPath/dataOut_exe_i [15]), .B(n2782), .Z(
        n8417) );
  HS65_LL_AND3X4 U7411 ( .A(\u_DataPath/cw_tomem_i [4]), .B(n3434), .C(n7352), 
        .Z(n3562) );
  HS65_LH_NAND2X4 U7412 ( .A(\u_DataPath/pc_4_to_ex_i [4]), .B(n7618), .Z(
        n7619) );
  HS65_LL_NOR2X2 U7413 ( .A(n8158), .B(n9066), .Z(n2948) );
  HS65_LH_IVX2 U7416 ( .A(n8698), .Z(n6760) );
  HS65_LH_BFX9 U7418 ( .A(n6109), .Z(n7510) );
  HS65_LH_NAND2X4 U7419 ( .A(n5709), .B(n5708), .Z(n5714) );
  HS65_LH_BFX9 U7420 ( .A(n7587), .Z(n7293) );
  HS65_LL_NAND3X2 U7421 ( .A(n7309), .B(n7216), .C(n7013), .Z(n3531) );
  HS65_LH_BFX9 U7422 ( .A(n8314), .Z(n7692) );
  HS65_LH_BFX9 U7423 ( .A(n8180), .Z(n7679) );
  HS65_LH_OAI21X3 U7424 ( .A(opcode_i[1]), .B(n7398), .C(n7611), .Z(n8020) );
  HS65_LL_MUXI21X2 U7426 ( .D0(\u_DataPath/from_alu_data_out_i [11]), .D1(
        \u_DataPath/from_mem_data_out_i [11]), .S0(n3148), .Z(n8213) );
  HS65_LHS_XNOR2X3 U7428 ( .A(\u_DataPath/pc_4_to_ex_i [2]), .B(n7420), .Z(
        \u_DataPath/u_execute/link_value_i [3]) );
  HS65_LH_OAI12X3 U7429 ( .A(n5710), .B(n5707), .C(n5709), .Z(n5533) );
  HS65_LL_MUXI21X2 U7430 ( .D0(\u_DataPath/from_alu_data_out_i [25]), .D1(
        \u_DataPath/from_mem_data_out_i [25]), .S0(n3148), .Z(n8445) );
  HS65_LH_IVX9 U7431 ( .A(write_byte_snps_wire), .Z(n3553) );
  HS65_LLS_XNOR2X3 U7432 ( .A(n7014), .B(n2893), .Z(n2910) );
  HS65_LH_OAI12X3 U7433 ( .A(n8975), .B(n8759), .C(n9024), .Z(n5819) );
  HS65_LL_NAND3X2 U7434 ( .A(n6488), .B(n7014), .C(n3529), .Z(n3530) );
  HS65_LL_MUXI21X2 U7435 ( .D0(\u_DataPath/from_alu_data_out_i [22]), .D1(
        \u_DataPath/from_mem_data_out_i [22]), .S0(n3235), .Z(n8273) );
  HS65_LH_BFX9 U7436 ( .A(n8183), .Z(n7684) );
  HS65_LL_NAND3X2 U7437 ( .A(n5279), .B(n5329), .C(n3292), .Z(n3293) );
  HS65_LL_NOR2X5 U7438 ( .A(n6182), .B(n6174), .Z(n6528) );
  HS65_LL_NOR2X5 U7439 ( .A(n6184), .B(n6176), .Z(n6530) );
  HS65_LH_MUXI21X2 U7440 ( .D0(\u_DataPath/from_alu_data_out_i [18]), .D1(
        \u_DataPath/from_mem_data_out_i [18]), .S0(n3148), .Z(n8145) );
  HS65_LL_NOR2X5 U7441 ( .A(n6182), .B(n6187), .Z(n2821) );
  HS65_LL_NOR2X3 U7442 ( .A(n6187), .B(n6184), .Z(n6340) );
  HS65_LHS_XNOR2X6 U7443 ( .A(n7331), .B(n7458), .Z(\u_DataPath/pc_4_i [4]) );
  HS65_LL_NOR2AX3 U7444 ( .A(n8463), .B(n3148), .Z(n2952) );
  HS65_LH_NOR2X5 U7445 ( .A(n5544), .B(n5574), .Z(n5546) );
  HS65_LH_NAND2X7 U7446 ( .A(\u_DataPath/jaddr_i [18]), .B(n5949), .Z(n5962)
         );
  HS65_LH_BFX9 U7449 ( .A(n6348), .Z(n6943) );
  HS65_LHS_XNOR2X6 U7451 ( .A(n9221), .B(n9058), .Z(n6478) );
  HS65_LHS_XNOR2X6 U7452 ( .A(n9168), .B(n9059), .Z(n6483) );
  HS65_LL_NOR2X3 U7453 ( .A(n6186), .B(n6187), .Z(n6347) );
  HS65_LHS_XNOR2X6 U7454 ( .A(n9467), .B(n9092), .Z(n6481) );
  HS65_LL_MUXI21X2 U7456 ( .D0(\u_DataPath/from_alu_data_out_i [19]), .D1(
        \u_DataPath/from_mem_data_out_i [19]), .S0(n3148), .Z(n8144) );
  HS65_LH_NAND2X4 U7457 ( .A(n5677), .B(n5676), .Z(n5679) );
  HS65_LH_NAND2X4 U7459 ( .A(n5559), .B(n5558), .Z(n5561) );
  HS65_LH_NAND2X4 U7460 ( .A(n5603), .B(n5606), .Z(n5588) );
  HS65_LH_AOI21X2 U7461 ( .A(n5575), .B(n5542), .C(n5541), .Z(n5543) );
  HS65_LH_NAND2X4 U7462 ( .A(n5602), .B(n5601), .Z(n5608) );
  HS65_LH_NAND2X4 U7463 ( .A(n5591), .B(n5590), .Z(n5599) );
  HS65_LH_NAND2X4 U7464 ( .A(n5631), .B(n5630), .Z(n5637) );
  HS65_LH_NAND2X4 U7465 ( .A(n5685), .B(n5684), .Z(n5687) );
  HS65_LL_NOR2X3 U7466 ( .A(n2909), .B(n2770), .Z(n2911) );
  HS65_LH_IVX4 U7467 ( .A(n5594), .Z(n5595) );
  HS65_LH_NAND2X4 U7468 ( .A(n5690), .B(n5689), .Z(n5694) );
  HS65_LL_AND2X4 U7469 ( .A(n3184), .B(n9431), .Z(n2836) );
  HS65_LH_NAND2X4 U7470 ( .A(n5691), .B(n5643), .Z(n5644) );
  HS65_LH_NAND2X4 U7471 ( .A(n5640), .B(n5639), .Z(n5642) );
  HS65_LH_NAND2X4 U7472 ( .A(n5652), .B(n5651), .Z(n5656) );
  HS65_LH_NAND2X4 U7473 ( .A(n5704), .B(n5703), .Z(n5706) );
  HS65_LH_NAND2X4 U7474 ( .A(n5618), .B(n5617), .Z(n5622) );
  HS65_LH_NAND2X4 U7475 ( .A(n5681), .B(n5680), .Z(n5683) );
  HS65_LL_AND2X4 U7476 ( .A(n3184), .B(n9427), .Z(n4878) );
  HS65_LH_NAND2X4 U7477 ( .A(n5662), .B(n5661), .Z(n5663) );
  HS65_LH_IVX4 U7478 ( .A(n5658), .Z(n5711) );
  HS65_LH_NAND2X4 U7479 ( .A(n5710), .B(n5657), .Z(n5659) );
  HS65_LH_NAND2X4 U7480 ( .A(n5853), .B(n5852), .Z(n5857) );
  HS65_LHS_XNOR2X6 U7481 ( .A(n9046), .B(n9465), .Z(n7202) );
  HS65_LH_NAND2X4 U7482 ( .A(n5762), .B(n5761), .Z(n5764) );
  HS65_LH_NAND2X4 U7483 ( .A(n5810), .B(n5809), .Z(n5816) );
  HS65_LH_NAND2X4 U7484 ( .A(n5900), .B(n5899), .Z(n5905) );
  HS65_LH_NAND2X4 U7485 ( .A(n5811), .B(n5814), .Z(n5791) );
  HS65_LH_NAND2X5 U7486 ( .A(n5737), .B(n5849), .Z(n5739) );
  HS65_LH_NAND2X4 U7487 ( .A(n5887), .B(n5886), .Z(n5889) );
  HS65_LH_NAND2X4 U7489 ( .A(n5799), .B(n5798), .Z(n5807) );
  HS65_LH_NAND2X4 U7490 ( .A(n5871), .B(n5870), .Z(n5873) );
  HS65_LH_IVX4 U7491 ( .A(n5802), .Z(n5803) );
  HS65_LH_CNIVX3 U7493 ( .A(n2804), .Z(n7931) );
  HS65_LH_NAND2X4 U7494 ( .A(n5901), .B(n5846), .Z(n5850) );
  HS65_LH_NOR2X3 U7495 ( .A(n9384), .B(rst), .Z(\u_DataPath/idex_rt_i [4]) );
  HS65_LH_NAND2X4 U7496 ( .A(n5877), .B(n5792), .Z(n5796) );
  HS65_LH_NAND2X4 U7497 ( .A(n5834), .B(n5833), .Z(n5838) );
  HS65_LH_BFX9 U7498 ( .A(n7688), .Z(n7691) );
  HS65_LH_BFX9 U7499 ( .A(n7688), .Z(n7689) );
  HS65_LH_NAND2X4 U7500 ( .A(n5825), .B(n5824), .Z(n5831) );
  HS65_LH_BFX9 U7501 ( .A(n7688), .Z(n7690) );
  HS65_LH_NAND2X4 U7502 ( .A(n5893), .B(n5844), .Z(n5845) );
  HS65_LH_NAND2AX7 U7503 ( .A(n2818), .B(n6169), .Z(n6176) );
  HS65_LH_NOR2X3 U7504 ( .A(\u_DataPath/immediate_ext_dec_i [0]), .B(n8053), 
        .Z(n7995) );
  HS65_LH_NAND2AX7 U7505 ( .A(n7712), .B(n9446), .Z(n8127) );
  HS65_LH_NAND2AX7 U7506 ( .A(n7714), .B(n8804), .Z(n8036) );
  HS65_LH_NAND2AX7 U7507 ( .A(n7712), .B(n8686), .Z(n8154) );
  HS65_LH_OAI12X3 U7508 ( .A(n5871), .B(n5770), .C(n5772), .Z(n5742) );
  HS65_LH_OAI12X3 U7510 ( .A(n5603), .B(n5600), .C(n5602), .Z(n5575) );
  HS65_LL_AND2X4 U7511 ( .A(n2906), .B(n2905), .Z(n2913) );
  HS65_LH_IVX4 U7512 ( .A(n5800), .Z(n5886) );
  HS65_LH_OAI12X3 U7513 ( .A(n5883), .B(n5832), .C(n5834), .Z(n5794) );
  HS65_LH_OAI12X3 U7514 ( .A(n5691), .B(n5688), .C(n5690), .Z(n5594) );
  HS65_LH_NAND2X4 U7515 ( .A(\u_DataPath/immediate_ext_dec_i [5]), .B(
        \u_DataPath/immediate_ext_dec_i [4]), .Z(n7412) );
  HS65_LH_OR2X4 U7516 ( .A(opcode_i[0]), .B(opcode_i[2]), .Z(n2819) );
  HS65_LH_BFX9 U7517 ( .A(n8181), .Z(n7681) );
  HS65_LH_OAI12X3 U7518 ( .A(n5865), .B(n5861), .C(n5863), .Z(n5859) );
  HS65_LH_NAND2X4 U7519 ( .A(n5724), .B(n5723), .Z(n5726) );
  HS65_LH_NAND2X4 U7520 ( .A(n5716), .B(n5715), .Z(n5718) );
  HS65_LH_OAI12X3 U7521 ( .A(n5907), .B(n5851), .C(n5853), .Z(n5848) );
  HS65_LH_NAND2X4 U7522 ( .A(n5610), .B(n5609), .Z(n5615) );
  HS65_LH_OAI12X3 U7523 ( .A(n5901), .B(n5898), .C(n5900), .Z(n5736) );
  HS65_LL_NOR2AX6 U7524 ( .A(n7647), .B(n2865), .Z(n3528) );
  HS65_LH_NAND2X4 U7525 ( .A(n5624), .B(n5623), .Z(n5628) );
  HS65_LH_OAI12X3 U7526 ( .A(n5681), .B(n5616), .C(n5618), .Z(n5625) );
  HS65_LH_OAI12X3 U7528 ( .A(n5887), .B(n5797), .C(n5799), .Z(n5740) );
  HS65_LL_IVX2 U7529 ( .A(n2908), .Z(n2909) );
  HS65_LH_OAI12X3 U7530 ( .A(n5677), .B(n5567), .C(n5569), .Z(n5541) );
  HS65_LH_OAI12X3 U7532 ( .A(n5704), .B(n5650), .C(n5652), .Z(n5647) );
  HS65_LL_NAND3X2 U7533 ( .A(\u_DataPath/cw_to_ex_i [0]), .B(n5329), .C(n5015), 
        .Z(n3213) );
  HS65_LH_BFX9 U7534 ( .A(n8184), .Z(n7688) );
  HS65_LH_NOR2X3 U7535 ( .A(n9168), .B(rst), .Z(\u_DataPath/rs_ex_i [2]) );
  HS65_LL_NOR2X2 U7536 ( .A(\u_DataPath/cw_to_ex_i [4]), .B(n3283), .Z(n3301)
         );
  HS65_LH_OAI12X3 U7538 ( .A(n5698), .B(n5695), .C(n5697), .Z(n5535) );
  HS65_LH_CNIVX3 U7539 ( .A(\u_DataPath/pc_4_to_ex_i [22]), .Z(n7306) );
  HS65_LH_OR2X9 U7540 ( .A(n8526), .B(\u_DataPath/pc_4_to_ex_i [29]), .Z(n5672) );
  HS65_LH_NOR2X3 U7541 ( .A(n8498), .B(\u_DataPath/u_execute/link_value_i [1]), 
        .Z(n5660) );
  HS65_LH_OR2X4 U7542 ( .A(n8500), .B(\u_DataPath/u_execute/link_value_i [0]), 
        .Z(n5531) );
  HS65_LH_OR2X9 U7543 ( .A(n8526), .B(\u_DataPath/pc_4_to_ex_i [27]), .Z(n5719) );
  HS65_LLS_XNOR2X3 U7544 ( .A(\u_DataPath/RFaddr_out_memwb_i [2]), .B(
        \u_DataPath/rs_ex_i [2]), .Z(n2875) );
  HS65_LLS_XNOR2X3 U7545 ( .A(\u_DataPath/rs_ex_i [0]), .B(
        \u_DataPath/RFaddr_out_memwb_i [0]), .Z(n2876) );
  HS65_LH_NOR2X5 U7546 ( .A(n8508), .B(\u_DataPath/pc_4_to_ex_i [12]), .Z(
        n5586) );
  HS65_LH_IVX7 U7547 ( .A(\u_DataPath/rs_ex_i [3]), .Z(n2872) );
  HS65_LH_NOR2X5 U7548 ( .A(n8526), .B(\u_DataPath/pc_4_to_ex_i [16]), .Z(
        n5619) );
  HS65_LH_IVX9 U7549 ( .A(n7649), .Z(\u_DataPath/regfile_addr_out_towb_i [4])
         );
  HS65_LH_OR2X9 U7550 ( .A(n8526), .B(\u_DataPath/pc_4_to_ex_i [18]), .Z(n5623) );
  HS65_LL_NAND2X2 U7551 ( .A(\u_DataPath/cw_to_ex_i [0]), .B(
        \u_DataPath/cw_to_ex_i [1]), .Z(n5328) );
  HS65_LH_IVX4 U7552 ( .A(\u_DataPath/pc_4_to_ex_i [18]), .Z(n7640) );
  HS65_LH_CNIVX3 U7553 ( .A(\u_DataPath/pc_4_to_ex_i [15]), .Z(n7430) );
  HS65_LH_OR2X9 U7554 ( .A(n8526), .B(\u_DataPath/pc_4_to_ex_i [20]), .Z(n5609) );
  HS65_LH_IVX9 U7555 ( .A(\u_DataPath/RFaddr_out_memwb_i [3]), .Z(n8027) );
  HS65_LLS_XNOR2X3 U7556 ( .A(\u_DataPath/idex_rt_i [4]), .B(
        \u_DataPath/RFaddr_out_memwb_i [4]), .Z(n2908) );
  HS65_LLS_XNOR2X3 U7557 ( .A(\u_DataPath/idex_rt_i [1]), .B(
        \u_DataPath/RFaddr_out_memwb_i [1]), .Z(n2906) );
  HS65_LH_OR2X9 U7558 ( .A(n8526), .B(\u_DataPath/pc_4_to_ex_i [23]), .Z(n5723) );
  HS65_LH_NOR2X5 U7559 ( .A(\u_DataPath/idex_rt_i [0]), .B(
        \u_DataPath/pc_4_to_ex_i [16]), .Z(n5835) );
  HS65_LH_IVX9 U7560 ( .A(\u_DataPath/data_read_ex_2_i [2]), .Z(n8378) );
  HS65_LH_NOR2X5 U7561 ( .A(n8524), .B(\u_DataPath/pc_4_to_ex_i [8]), .Z(n5895) );
  HS65_LH_NOR2X5 U7562 ( .A(n8465), .B(\u_DataPath/pc_4_to_ex_i [2]), .Z(n5915) );
  HS65_LH_NOR2X5 U7563 ( .A(n8522), .B(\u_DataPath/pc_4_to_ex_i [5]), .Z(n5851) );
  HS65_LH_NOR2X5 U7564 ( .A(n8504), .B(\u_DataPath/pc_4_to_ex_i [14]), .Z(
        n5773) );
  HS65_LH_NOR2X5 U7565 ( .A(n8469), .B(\u_DataPath/pc_4_to_ex_i [10]), .Z(
        n5800) );
  HS65_LH_NOR2X5 U7568 ( .A(\u_DataPath/idex_rt_i [2]), .B(
        \u_DataPath/pc_4_to_ex_i [18]), .Z(n5879) );
  HS65_LL_NOR2AX6 U7569 ( .A(n2891), .B(n2890), .Z(\lte_x_57/B[30] ) );
  HS65_LL_AO22X4 U7571 ( .A(\lte_x_57/B[4] ), .B(n7680), .C(n7682), .D(
        \u_DataPath/u_execute/resAdd1_i [4]), .Z(
        \u_DataPath/jump_address_i [4]) );
  HS65_LL_NOR2AX3 U7573 ( .A(n4256), .B(n4255), .Z(n4267) );
  HS65_LH_CBI4I1X3 U7574 ( .A(n5296), .B(n5295), .C(n5294), .D(n5293), .Z(
        n5307) );
  HS65_LL_MUXI21X2 U7575 ( .D0(\u_DataPath/from_alu_data_out_i [8]), .D1(
        \u_DataPath/from_mem_data_out_i [8]), .S0(n3235), .Z(n8228) );
  HS65_LL_NOR2AX3 U7576 ( .A(n8280), .B(n8339), .Z(n7669) );
  HS65_LLS_XNOR2X3 U7577 ( .A(n3894), .B(n3893), .Z(n3895) );
  HS65_LH_CNIVX3 U7578 ( .A(\u_DataPath/RFaddr_out_memwb_i [4]), .Z(n7941) );
  HS65_LL_AOI12X2 U7581 ( .A(n5423), .B(n5422), .C(n5421), .Z(n5431) );
  HS65_LL_NAND3X5 U7582 ( .A(n3484), .B(n3823), .C(n3483), .Z(n4573) );
  HS65_LL_NOR2AX3 U7585 ( .A(n2786), .B(\sub_x_51/A[13] ), .Z(n4077) );
  HS65_LLS_XNOR2X3 U7586 ( .A(n4096), .B(n4095), .Z(n4097) );
  HS65_LL_NAND4ABX3 U7587 ( .A(n3955), .B(n3947), .C(n3946), .D(n3945), .Z(
        n3968) );
  HS65_LL_CBI4I1X3 U7589 ( .A(n5227), .B(n5408), .C(n5384), .D(n4895), .Z(
        n4896) );
  HS65_LL_OAI13X1 U7590 ( .A(n3039), .B(n3073), .C(n5375), .D(n5376), .Z(n5026) );
  HS65_LL_AOI12X2 U7591 ( .A(n5118), .B(n5117), .C(n5116), .Z(n5119) );
  HS65_LL_NOR2AX3 U7593 ( .A(n3940), .B(n9538), .Z(n5343) );
  HS65_LL_AO12X4 U7596 ( .A(n3796), .B(n4842), .C(n3746), .Z(n3747) );
  HS65_LL_AOI12X2 U7597 ( .A(\sub_x_51/A[18] ), .B(n3742), .C(n3723), .Z(n3726) );
  HS65_LL_AND2X4 U7598 ( .A(n2804), .B(\u_DataPath/jaddr_i [18]), .Z(n5938) );
  HS65_LL_NOR3AX2 U7599 ( .A(n3574), .B(n3825), .C(n3820), .Z(n3576) );
  HS65_LL_NOR2AX3 U7600 ( .A(n3093), .B(n3092), .Z(n3094) );
  HS65_LL_NOR2X2 U7601 ( .A(n5304), .B(n5004), .Z(n4920) );
  HS65_LH_NOR2AX3 U7604 ( .A(n5426), .B(n5372), .Z(n4895) );
  HS65_LL_AND2X4 U7607 ( .A(n3184), .B(n9137), .Z(n3219) );
  HS65_LH_NOR3X1 U7610 ( .A(n4879), .B(n4878), .C(n4877), .Z(n4882) );
  HS65_LH_AOI21X2 U7611 ( .A(n5103), .B(n5102), .C(n5101), .Z(n5104) );
  HS65_LH_AOI21X2 U7612 ( .A(n5144), .B(n5143), .C(n5142), .Z(n5153) );
  HS65_LL_NOR2AX3 U7614 ( .A(n3958), .B(n3957), .Z(n3959) );
  HS65_LL_NAND2AX4 U7615 ( .A(n3972), .B(n3956), .Z(n3957) );
  HS65_LH_NAND2X2 U7616 ( .A(n5043), .B(n5347), .Z(n3944) );
  HS65_LHS_XNOR2X3 U7617 ( .A(\lte_x_57/B[11] ), .B(n5077), .Z(n4971) );
  HS65_LL_NOR2AX3 U7618 ( .A(n3694), .B(n4203), .Z(n3695) );
  HS65_LH_OAI21X2 U7619 ( .A(n4794), .B(n3075), .C(n3379), .Z(n3694) );
  HS65_LL_NAND4ABX3 U7620 ( .A(n8435), .B(n3184), .C(n3183), .D(n8437), .Z(
        n3185) );
  HS65_LH_AOI22X1 U7621 ( .A(\sub_x_51/A[18] ), .B(n2792), .C(n5498), .D(
        \sub_x_51/A[20] ), .Z(n3383) );
  HS65_LLS_XNOR2X3 U7623 ( .A(\sub_x_51/A[5] ), .B(n3949), .Z(n4954) );
  HS65_LH_AO22X4 U7624 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][27] ), .B(n9010), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][27] ), .D(
        n9189), .Z(n6324) );
  HS65_LH_AOI22X1 U7625 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][27] ), .B(n8865), 
        .C(n9256), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][27] ), .Z(n7165)
         );
  HS65_LH_AOI22X1 U7626 ( .A(n8868), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][27] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][27] ), .D(n9197), 
        .Z(n7162) );
  HS65_LH_AOI22X1 U7627 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][14] ), .B(n8884), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][14] ), .D(
        n9193), .Z(n6875) );
  HS65_LH_AOI22X1 U7628 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][14] ), .B(n9259), 
        .C(n9256), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][14] ), .Z(n6089)
         );
  HS65_LH_AOI22X1 U7629 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][15] ), .B(n9259), 
        .C(n8864), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][15] ), .Z(n7267)
         );
  HS65_LH_AOI22X1 U7630 ( .A(n9243), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][15] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][15] ), .D(n9197), 
        .Z(n7264) );
  HS65_LH_AO22X4 U7631 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][11] ), .B(n9187), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][11] ), .D(
        n8852), .Z(n6504) );
  HS65_LH_AOI22X1 U7632 ( .A(n8868), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][11] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][11] ), .D(n9197), 
        .Z(n6807) );
  HS65_LH_AO22X4 U7633 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][19] ), .B(n9154), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][19] ), .D(
        n9194), .Z(n6291) );
  HS65_LH_AO22X4 U7634 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][19] ), .B(n9010), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][19] ), .D(
        n9189), .Z(n6303) );
  HS65_LH_AOI22X1 U7635 ( .A(n9243), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][19] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][19] ), .D(n9009), 
        .Z(n6767) );
  HS65_LH_AOI22X1 U7636 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][3] ), .B(n9259), 
        .C(n8864), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][3] ), .Z(n6124)
         );
  HS65_LH_AOI22X1 U7637 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][10] ), .B(n8884), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][10] ), .D(
        n9193), .Z(n6717) );
  HS65_LH_AOI22X1 U7638 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][10] ), .B(n9259), 
        .C(n9256), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][10] ), .Z(n7045)
         );
  HS65_LH_AOI22X1 U7639 ( .A(n9243), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][10] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][10] ), .D(n9009), 
        .Z(n7042) );
  HS65_LH_AOI22X1 U7640 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][26] ), .B(n8884), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][26] ), .D(
        n9193), .Z(n6945) );
  HS65_LH_AOI22X1 U7641 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][26] ), .B(n8865), 
        .C(n9256), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][26] ), .Z(n6790)
         );
  HS65_LH_AOI22X1 U7642 ( .A(n8868), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][26] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][26] ), .D(n9197), 
        .Z(n6787) );
  HS65_LH_AO22X4 U7643 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][23] ), .B(n9187), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][23] ), .D(
        n8852), .Z(n6334) );
  HS65_LH_AOI22X1 U7644 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][23] ), .B(n8865), 
        .C(n9256), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][23] ), .Z(n7125)
         );
  HS65_LH_AOI22X1 U7645 ( .A(n8868), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][23] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][23] ), .D(n9197), 
        .Z(n7122) );
  HS65_LH_AOI22X1 U7646 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][30] ), .B(n9159), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][30] ), .D(
        n8862), .Z(n7533) );
  HS65_LH_AOI22X1 U7647 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][12] ), .B(n8884), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][12] ), .D(
        n9193), .Z(n6697) );
  HS65_LH_AOI22X1 U7648 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][12] ), .B(n8865), 
        .C(n9256), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][12] ), .Z(n7145)
         );
  HS65_LH_AOI22X1 U7649 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][7] ), .B(n8884), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][7] ), .D(n9193), .Z(n6471) );
  HS65_LH_AO22X4 U7650 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][7] ), .B(n9187), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][7] ), .D(
        n8852), .Z(n6462) );
  HS65_LH_AOI22X1 U7651 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][7] ), .B(n9259), 
        .C(n8864), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][7] ), .Z(n6049)
         );
  HS65_LH_AOI22X1 U7652 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][13] ), .B(n9226), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][13] ), .D(
        n9193), .Z(n6410) );
  HS65_LH_AOI22X1 U7653 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][13] ), .B(n9259), 
        .C(n8864), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][13] ), .Z(n7025)
         );
  HS65_LH_AOI22X1 U7654 ( .A(n9243), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][13] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][13] ), .D(n9009), 
        .Z(n7022) );
  HS65_LH_AOI22X1 U7655 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][29] ), .B(n9259), 
        .C(n8864), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][29] ), .Z(n7561)
         );
  HS65_LH_AOI22X1 U7656 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][21] ), .B(n8865), 
        .C(n9256), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][21] ), .Z(n6003)
         );
  HS65_LH_AOI22X1 U7657 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][5] ), .B(n8865), 
        .C(n9256), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][5] ), .Z(n7085)
         );
  HS65_LH_AOI22X1 U7658 ( .A(n8868), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][5] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][5] ), .D(n9197), 
        .Z(n7082) );
  HS65_LH_AOI22X1 U7659 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][25] ), .B(n8884), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][25] ), .D(
        n9193), .Z(n6965) );
  HS65_LH_AOI22X1 U7660 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][25] ), .B(n9259), 
        .C(n8864), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][25] ), .Z(n7485)
         );
  HS65_LH_AOI22X1 U7661 ( .A(n9243), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][25] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][25] ), .D(n9009), 
        .Z(n7482) );
  HS65_LH_AOI22X1 U7662 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][9] ), .B(n8884), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][9] ), .D(n9193), .Z(n7005) );
  HS65_LH_AOI22X1 U7663 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][9] ), .B(n8865), 
        .C(n9256), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][9] ), .Z(n7065)
         );
  HS65_LH_AOI22X1 U7664 ( .A(n8868), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][9] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][9] ), .D(n9197), 
        .Z(n7062) );
  HS65_LH_AOI22X1 U7665 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][24] ), .B(n9226), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][24] ), .D(
        n9193), .Z(n6280) );
  HS65_LH_AO22X4 U7666 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][24] ), .B(n9154), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][24] ), .D(
        n9194), .Z(n6268) );
  HS65_LH_AOI22X1 U7667 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][24] ), .B(n9259), 
        .C(n8864), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][24] ), .Z(n5983)
         );
  HS65_LH_AOI22X1 U7668 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][28] ), .B(n8865), 
        .C(n9256), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][28] ), .Z(n7596)
         );
  HS65_LH_AOI22X1 U7669 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][28] ), .B(n9159), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][28] ), .D(
        n8862), .Z(n7583) );
  HS65_LH_AOI22X1 U7670 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][22] ), .B(n9259), 
        .C(n8864), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][22] ), .Z(n7185)
         );
  HS65_LH_AOI22X1 U7671 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][4] ), .B(n9259), 
        .C(n8864), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][4] ), .Z(n6029)
         );
  HS65_LH_AOI22X1 U7672 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][8] ), .B(n8884), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][8] ), .D(n9193), .Z(n6657) );
  HS65_LH_AOI22X1 U7673 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][8] ), .B(n8865), 
        .C(n9256), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][8] ), .Z(n6850)
         );
  HS65_LH_AOI22X1 U7674 ( .A(n8868), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][8] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][8] ), .D(n9197), 
        .Z(n6847) );
  HS65_LH_AOI22X1 U7675 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][20] ), .B(n9259), 
        .C(n8864), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][20] ), .Z(n7105)
         );
  HS65_LH_AOI22X1 U7676 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][17] ), .B(n8865), 
        .C(n9256), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][17] ), .Z(n5954)
         );
  HS65_LH_AOI22X1 U7677 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][2] ), .B(n9259), 
        .C(n8864), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][2] ), .Z(n6151)
         );
  HS65_LH_AOI22X1 U7678 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][18] ), .B(n8884), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][18] ), .D(
        n9193), .Z(n6677) );
  HS65_LH_AOI22X1 U7679 ( .A(n9243), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][18] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][18] ), .D(n9009), 
        .Z(n7224) );
  HS65_LH_AOI22X1 U7680 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][6] ), .B(n8884), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][6] ), .D(n9193), .Z(n6741) );
  HS65_LH_AOI22X1 U7681 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][6] ), .B(n8865), 
        .C(n9256), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][6] ), .Z(n6830)
         );
  HS65_LH_AOI22X1 U7682 ( .A(n8868), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][6] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][6] ), .D(n9197), 
        .Z(n6827) );
  HS65_LH_AOI22X1 U7683 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][1] ), .B(n9226), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][1] ), .D(n9193), .Z(n6251) );
  HS65_LH_BFX9 U7684 ( .A(n6122), .Z(n7500) );
  HS65_LH_AOI22X1 U7685 ( .A(n9243), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][1] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][1] ), .D(n9009), 
        .Z(n7244) );
  HS65_LH_BFX9 U7686 ( .A(n7003), .Z(n6635) );
  HS65_LH_NOR2X6 U7687 ( .A(n6188), .B(n6164), .Z(n6977) );
  HS65_LH_NOR2X2 U7688 ( .A(\sub_x_51/A[13] ), .B(n2786), .Z(n5083) );
  HS65_LL_NOR2X2 U7689 ( .A(n4709), .B(n4458), .Z(n5068) );
  HS65_LH_OAI21X2 U7690 ( .A(n5030), .B(n5364), .C(n5367), .Z(n5031) );
  HS65_LL_NOR2AX3 U7691 ( .A(n5027), .B(n5366), .Z(n5394) );
  HS65_LH_NAND3X2 U7692 ( .A(n5417), .B(n5043), .C(n5416), .Z(n5046) );
  HS65_LL_NAND2X2 U7693 ( .A(n5412), .B(n5044), .Z(n5045) );
  HS65_LH_AOI21X2 U7697 ( .A(n3963), .B(n5360), .C(n5366), .Z(n3964) );
  HS65_LL_NAND4ABX3 U7698 ( .A(n8403), .B(n3184), .C(n8405), .D(n8404), .Z(
        n3011) );
  HS65_LH_AOI21X2 U7700 ( .A(n4781), .B(n5201), .C(n4309), .Z(n4285) );
  HS65_LLS_XNOR2X3 U7701 ( .A(n5187), .B(n4910), .Z(n4946) );
  HS65_LL_NAND4ABX3 U7704 ( .A(n4317), .B(n4316), .C(n4315), .D(n4314), .Z(
        n4793) );
  HS65_LL_NOR2AX3 U7709 ( .A(n2968), .B(n4871), .Z(n2969) );
  HS65_LH_NOR3X1 U7710 ( .A(opcode_i[1]), .B(opcode_i[0]), .C(n7608), .Z(n7609) );
  HS65_LH_AOI22X1 U7712 ( .A(n8868), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][3] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][3] ), .D(n9197), 
        .Z(n6117) );
  HS65_LLS_XNOR2X3 U7713 ( .A(n4494), .B(n4493), .Z(n4495) );
  HS65_LH_AOI22X1 U7715 ( .A(n8868), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][2] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][2] ), .D(n9197), 
        .Z(n6148) );
  HS65_LH_OAI21X2 U7718 ( .A(opcode_i[5]), .B(n7966), .C(n7615), .Z(n7394) );
  HS65_LH_CNIVX3 U7719 ( .A(n5879), .Z(n5792) );
  HS65_LH_CNIVX3 U7720 ( .A(n5832), .Z(n5833) );
  HS65_LH_CNIVX3 U7721 ( .A(n5895), .Z(n5844) );
  HS65_LH_CNIVX3 U7722 ( .A(n5808), .Z(n5809) );
  HS65_LH_CNIVX3 U7723 ( .A(n5898), .Z(n5899) );
  HS65_LH_CNIVX3 U7724 ( .A(n5797), .Z(n5798) );
  HS65_LH_AOI22X1 U7725 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][27] ), .B(n8859), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][27] ), .D(
        n9116), .Z(n6310) );
  HS65_LH_AOI22X1 U7726 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][27] ), .B(n8851), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][27] ), .D(
        n8850), .Z(n6318) );
  HS65_LH_AOI22X1 U7727 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][27] ), .B(n9162), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][27] ), .D(
        n8854), .Z(n6315) );
  HS65_LH_AO22X4 U7728 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][27] ), .B(n9160), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][27] ), .D(
        n9267), .Z(n6323) );
  HS65_LH_AOI22X1 U7729 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][27] ), .B(n9226), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][27] ), .D(
        n8848), .Z(n6322) );
  HS65_LH_AOI22X1 U7730 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][27] ), .B(n9159), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][27] ), .D(
        n8862), .Z(n7169) );
  HS65_LH_AOI22X1 U7731 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][27] ), .B(n9113), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][27] ), .D(
        n8861), .Z(n7168) );
  HS65_LH_AOI22X1 U7732 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][27] ), .B(n9096), 
        .C(n9158), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][27] ), .Z(n7158)
         );
  HS65_LH_AO22X4 U7733 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][27] ), .B(n8947), 
        .C(n8946), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][27] ), .Z(n7157)
         );
  HS65_LH_AO22X4 U7734 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][27] ), .B(n8948), 
        .C(n8951), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][27] ), .Z(n7156)
         );
  HS65_LH_AOI22X1 U7735 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][27] ), .B(n9062), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][27] ), .D(
        n8863), .Z(n7164) );
  HS65_LH_AO22X4 U7736 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][27] ), .B(n9165), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][27] ), .D(
        n9065), .Z(n7160) );
  HS65_LH_AO22X4 U7737 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][27] ), .B(n9153), 
        .C(n9068), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][27] ), .Z(n7161)
         );
  HS65_LH_AOI22X1 U7738 ( .A(n9161), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][27] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][27] ), .D(n9095), 
        .Z(n7163) );
  HS65_LH_AOI22X1 U7739 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][14] ), .B(n8937), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][14] ), .D(
        n9067), .Z(n6870) );
  HS65_LH_AOI22X1 U7740 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][14] ), .B(n8860), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][14] ), .D(
        n9157), .Z(n6865) );
  HS65_LH_AO22X4 U7741 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][14] ), .B(n8885), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][14] ), .D(
        n8856), .Z(n6862) );
  HS65_LH_AOI22X1 U7742 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][14] ), .B(n8933), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][14] ), .D(
        n9240), .Z(n6874) );
  HS65_LH_AO22X4 U7743 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][14] ), .B(n9010), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][14] ), .D(
        n9189), .Z(n6877) );
  HS65_LH_AOI22X1 U7744 ( .A(n9243), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][14] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][14] ), .D(n9009), 
        .Z(n6086) );
  HS65_LH_AO22X4 U7745 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][14] ), .B(n8947), 
        .C(n8946), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][14] ), .Z(n6081)
         );
  HS65_LH_AOI22X1 U7746 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][14] ), .B(n9096), 
        .C(n9158), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][14] ), .Z(n6082)
         );
  HS65_LH_AOI22X1 U7747 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][14] ), .B(n9098), 
        .C(n9100), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][14] ), .Z(n6083)
         );
  HS65_LH_AO22X4 U7748 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][14] ), .B(n9070), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][14] ), .D(
        n9064), .Z(n6094) );
  HS65_LH_AOI22X1 U7749 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][15] ), .B(n9246), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][15] ), .D(
        n9067), .Z(n6891) );
  HS65_LH_AOI22X1 U7750 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][15] ), .B(n8860), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][15] ), .D(
        n9157), .Z(n6885) );
  HS65_LH_AO22X4 U7751 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][15] ), .B(n8885), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][15] ), .D(
        n8856), .Z(n6882) );
  HS65_LH_AOI22X1 U7752 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][15] ), .B(n8884), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][15] ), .D(
        n8848), .Z(n6897) );
  HS65_LH_AO22X4 U7753 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][15] ), .B(n9260), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][15] ), .D(
        n9189), .Z(n6899) );
  HS65_LH_AO22X4 U7754 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][15] ), .B(n9070), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][15] ), .D(
        n9064), .Z(n7272) );
  HS65_LH_AOI22X1 U7755 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][15] ), .B(n9098), 
        .C(n9200), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][15] ), .Z(n7261)
         );
  HS65_LH_AO22X4 U7756 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][15] ), .B(n9206), 
        .C(n9205), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][15] ), .Z(n7259)
         );
  HS65_LH_AO22X4 U7757 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][15] ), .B(n9204), 
        .C(n9203), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][15] ), .Z(n7258)
         );
  HS65_LH_AOI22X1 U7758 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][15] ), .B(n9062), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][15] ), .D(
        n8863), .Z(n7266) );
  HS65_LH_AO22X4 U7759 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][15] ), .B(n9165), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][15] ), .D(
        n9245), .Z(n7262) );
  HS65_LH_AOI22X1 U7760 ( .A(n9161), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][15] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][15] ), .D(n9095), 
        .Z(n7265) );
  HS65_LH_AOI22X1 U7761 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][11] ), .B(n8937), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][11] ), .D(
        n9262), .Z(n6508) );
  HS65_LH_AOI22X1 U7762 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][11] ), .B(n8933), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][11] ), .D(
        n9163), .Z(n6512) );
  HS65_LH_AO22X4 U7763 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][11] ), .B(n9260), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][11] ), .D(
        n9189), .Z(n6515) );
  HS65_LH_AO22X4 U7764 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][11] ), .B(n9469), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][11] ), .D(
        n8853), .Z(n6505) );
  HS65_LH_AOI22X1 U7765 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][11] ), .B(n9159), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][11] ), .D(
        n8862), .Z(n6814) );
  HS65_LH_AOI22X1 U7766 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][11] ), .B(n9098), 
        .C(n9200), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][11] ), .Z(n6804)
         );
  HS65_LH_AO22X4 U7767 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][11] ), .B(n9206), 
        .C(n8946), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][11] ), .Z(n6802)
         );
  HS65_LH_AO22X4 U7768 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][11] ), .B(n9204), 
        .C(n8951), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][11] ), .Z(n6801)
         );
  HS65_LH_AOI22X1 U7769 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][11] ), .B(n9062), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][11] ), .D(
        n8863), .Z(n6809) );
  HS65_LH_AO22X4 U7770 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][11] ), .B(n9165), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][11] ), .D(
        n9065), .Z(n6805) );
  HS65_LH_AO22X4 U7771 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][11] ), .B(n9153), 
        .C(n9068), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][11] ), .Z(n6806)
         );
  HS65_LH_AOI22X1 U7772 ( .A(n9161), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][11] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][11] ), .D(n9095), 
        .Z(n6808) );
  HS65_LH_AOI22X1 U7773 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][19] ), .B(n9246), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][19] ), .D(
        n9067), .Z(n6295) );
  HS65_LH_AOI22X1 U7774 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][19] ), .B(n9162), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][19] ), .D(
        n8854), .Z(n6293) );
  HS65_LH_AOI22X1 U7775 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][19] ), .B(n9191), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][19] ), .D(
        n8855), .Z(n6294) );
  HS65_LH_AO22X4 U7776 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][19] ), .B(n9160), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][19] ), .D(
        n9267), .Z(n6302) );
  HS65_LH_AOI22X1 U7777 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][19] ), .B(n9226), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][19] ), .D(
        n8848), .Z(n6301) );
  HS65_LH_AOI22X1 U7778 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][19] ), .B(n9096), 
        .C(n9158), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][19] ), .Z(n6763)
         );
  HS65_LH_AO22X4 U7779 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][19] ), .B(n8947), 
        .C(n8946), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][19] ), .Z(n6762)
         );
  HS65_LH_AO22X4 U7780 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][19] ), .B(n8948), 
        .C(n8951), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][19] ), .Z(n6761)
         );
  HS65_LH_AO22X4 U7781 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][19] ), .B(n9070), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][19] ), .D(
        n9064), .Z(n6775) );
  HS65_LH_AO22X4 U7782 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][19] ), .B(n9152), 
        .C(n9097), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][19] ), .Z(n6776)
         );
  HS65_LH_AOI22X1 U7783 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][19] ), .B(n9113), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][19] ), .D(
        n8861), .Z(n6773) );
  HS65_LH_AO22X4 U7784 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][19] ), .B(n8867), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][19] ), .D(
        n8866), .Z(n6771) );
  HS65_LH_AO22X4 U7785 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][19] ), .B(n9102), 
        .C(n9101), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][19] ), .Z(n6772)
         );
  HS65_LH_AO22X4 U7786 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][3] ), .B(n8939), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][3] ), .D(
        n9155), .Z(n6447) );
  HS65_LH_AOI22X1 U7787 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][3] ), .B(n9246), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][3] ), .D(n9067), .Z(n6445) );
  HS65_LH_AOI22X1 U7788 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][3] ), .B(n8859), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][3] ), .D(
        n9116), .Z(n6439) );
  HS65_LH_AOI22X1 U7789 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][3] ), .B(n8950), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][3] ), .D(
        n8855), .Z(n6444) );
  HS65_LH_AOI22X1 U7790 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][3] ), .B(n9159), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][3] ), .D(n8862), .Z(n6135) );
  HS65_LH_AOI22X1 U7791 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][3] ), .B(n9098), 
        .C(n9200), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][3] ), .Z(n6107)
         );
  HS65_LH_AO22X4 U7792 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][3] ), .B(n9206), 
        .C(n9205), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][3] ), .Z(n6105)
         );
  HS65_LH_AO22X4 U7793 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][3] ), .B(n9204), 
        .C(n9203), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][3] ), .Z(n6104)
         );
  HS65_LH_AOI22X1 U7794 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][3] ), .B(n9062), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][3] ), .D(n8863), .Z(n6123) );
  HS65_LH_AO22X4 U7795 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][10] ), .B(n9154), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][10] ), .D(
        n8852), .Z(n6708) );
  HS65_LH_AO22X4 U7796 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][10] ), .B(n9156), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][10] ), .D(
        n8853), .Z(n6709) );
  HS65_LH_AOI22X1 U7797 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][10] ), .B(n8933), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][10] ), .D(
        n9240), .Z(n6716) );
  HS65_LH_AO22X4 U7798 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][10] ), .B(n9260), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][10] ), .D(
        n9189), .Z(n6719) );
  HS65_LH_AOI22X1 U7799 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][10] ), .B(n8937), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][10] ), .D(
        n9262), .Z(n6712) );
  HS65_LH_AO22X4 U7800 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][10] ), .B(n8940), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][10] ), .D(
        n8949), .Z(n6715) );
  HS65_LH_AOI22X1 U7801 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][10] ), .B(n9096), 
        .C(n9158), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][10] ), .Z(n7038)
         );
  HS65_LH_AO22X4 U7802 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][10] ), .B(n8947), 
        .C(n8946), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][10] ), .Z(n7037)
         );
  HS65_LH_AO22X4 U7803 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][10] ), .B(n8948), 
        .C(n8951), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][10] ), .Z(n7036)
         );
  HS65_LH_AO22X4 U7804 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][10] ), .B(n9070), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][10] ), .D(
        n9064), .Z(n7050) );
  HS65_LH_AO22X4 U7805 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][10] ), .B(n9152), 
        .C(n9097), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][10] ), .Z(n7051)
         );
  HS65_LH_AO22X4 U7806 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][10] ), .B(n8867), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][10] ), .D(
        n8866), .Z(n7046) );
  HS65_LH_AO22X4 U7807 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][10] ), .B(n9102), 
        .C(n9101), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][10] ), .Z(n7047)
         );
  HS65_LH_AOI22X1 U7808 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][26] ), .B(n8937), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][26] ), .D(
        n9067), .Z(n6939) );
  HS65_LH_AOI22X1 U7809 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][26] ), .B(n8860), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][26] ), .D(
        n9157), .Z(n6934) );
  HS65_LH_AO22X4 U7810 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][26] ), .B(n8885), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][26] ), .D(
        n8856), .Z(n6931) );
  HS65_LH_AOI22X1 U7811 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][26] ), .B(n8933), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][26] ), .D(
        n9240), .Z(n6944) );
  HS65_LH_AO22X4 U7812 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][26] ), .B(n9260), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][26] ), .D(
        n9189), .Z(n6947) );
  HS65_LH_AO22X4 U7813 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][26] ), .B(n9154), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][26] ), .D(
        n8852), .Z(n6935) );
  HS65_LH_AOI22X1 U7814 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][26] ), .B(n9159), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][26] ), .D(
        n8862), .Z(n6794) );
  HS65_LH_AOI22X1 U7815 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][26] ), .B(n9098), 
        .C(n9200), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][26] ), .Z(n6784)
         );
  HS65_LH_AO22X4 U7816 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][26] ), .B(n9206), 
        .C(n9205), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][26] ), .Z(n6782)
         );
  HS65_LH_AO22X4 U7817 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][26] ), .B(n9204), 
        .C(n9203), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][26] ), .Z(n6781)
         );
  HS65_LH_AOI22X1 U7818 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][26] ), .B(n9062), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][26] ), .D(
        n8863), .Z(n6789) );
  HS65_LH_AO22X4 U7819 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][26] ), .B(n9165), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][26] ), .D(
        n9065), .Z(n6785) );
  HS65_LH_AO22X4 U7820 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][26] ), .B(n9153), 
        .C(n9068), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][26] ), .Z(n6786)
         );
  HS65_LH_AOI22X1 U7821 ( .A(n9161), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][26] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][26] ), .D(n9095), 
        .Z(n6788) );
  HS65_LH_AOI22X1 U7822 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][23] ), .B(n8937), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][23] ), .D(
        n9262), .Z(n6341) );
  HS65_LH_AOI22X1 U7823 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][23] ), .B(n8859), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][23] ), .D(
        n9116), .Z(n6331) );
  HS65_LH_AOI22X1 U7824 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][23] ), .B(n8933), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][23] ), .D(
        n9163), .Z(n6349) );
  HS65_LH_AO22X4 U7825 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][23] ), .B(n9260), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][23] ), .D(
        n9189), .Z(n6352) );
  HS65_LH_AO22X4 U7826 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][23] ), .B(n9469), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][23] ), .D(
        n8853), .Z(n6335) );
  HS65_LH_AOI22X1 U7827 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][23] ), .B(n9159), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][23] ), .D(
        n8862), .Z(n7129) );
  HS65_LH_AOI22X1 U7828 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][23] ), .B(n9096), 
        .C(n9158), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][23] ), .Z(n7118)
         );
  HS65_LH_AO22X4 U7829 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][23] ), .B(n8947), 
        .C(n8946), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][23] ), .Z(n7117)
         );
  HS65_LH_AO22X4 U7830 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][23] ), .B(n8948), 
        .C(n8951), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][23] ), .Z(n7116)
         );
  HS65_LH_AOI22X1 U7831 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][23] ), .B(n9062), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][23] ), .D(
        n8863), .Z(n7124) );
  HS65_LH_AO22X4 U7832 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][23] ), .B(n9165), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][23] ), .D(
        n9065), .Z(n7120) );
  HS65_LH_AO22X4 U7833 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][23] ), .B(n9153), 
        .C(n9068), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][23] ), .Z(n7121)
         );
  HS65_LH_AOI22X1 U7834 ( .A(n9161), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][23] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][23] ), .D(n9095), 
        .Z(n7123) );
  HS65_LH_AOI22X1 U7835 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][30] ), .B(n9246), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][30] ), .D(
        n9067), .Z(n6571) );
  HS65_LH_AOI22X1 U7836 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][30] ), .B(n8938), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][30] ), .D(
        n8850), .Z(n6572) );
  HS65_LH_AOI22X1 U7837 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][30] ), .B(n9226), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][30] ), .D(
        n8848), .Z(n6576) );
  HS65_LH_AO22X4 U7838 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][30] ), .B(n9160), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][30] ), .D(
        n9164), .Z(n6577) );
  HS65_LH_AOI22X1 U7839 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][30] ), .B(n9248), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][30] ), .D(
        n9163), .Z(n6575) );
  HS65_LH_AO22X4 U7840 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][30] ), .B(n9010), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][30] ), .D(
        n8849), .Z(n6578) );
  HS65_LH_AO22X4 U7841 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][30] ), .B(n8885), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][30] ), .D(
        n8856), .Z(n6563) );
  HS65_LH_AOI22X1 U7842 ( .A(n8868), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][30] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][30] ), .D(n9197), 
        .Z(n7535) );
  HS65_LH_AOI22X1 U7843 ( .A(n9161), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][30] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][30] ), .D(n9095), 
        .Z(n7536) );
  HS65_LH_AO22X4 U7844 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][30] ), .B(n9166), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[9][30] ), .D(
        n9113), .Z(n7537) );
  HS65_LH_AO22X4 U7845 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][30] ), .B(n9153), 
        .C(n9068), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][30] ), .Z(n7542)
         );
  HS65_LH_AOI22X1 U7846 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][30] ), .B(n8865), 
        .C(n8864), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][30] ), .Z(n7539)
         );
  HS65_LH_AO22X4 U7847 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][30] ), .B(n9165), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][30] ), .D(
        n9065), .Z(n7541) );
  HS65_LH_AOI22X1 U7848 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][30] ), .B(n9062), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][30] ), .D(
        n8863), .Z(n7534) );
  HS65_LH_AO22X4 U7849 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][30] ), .B(n9102), 
        .C(n9101), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][30] ), .Z(n7532)
         );
  HS65_LH_AO22X4 U7850 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][12] ), .B(n9154), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][12] ), .D(
        n8852), .Z(n6688) );
  HS65_LH_AO22X4 U7851 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][12] ), .B(n9156), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][12] ), .D(
        n8853), .Z(n6689) );
  HS65_LH_AOI22X1 U7852 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][12] ), .B(n8933), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][12] ), .D(
        n9240), .Z(n6696) );
  HS65_LH_AO22X4 U7853 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][12] ), .B(n9260), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][12] ), .D(
        n9189), .Z(n6699) );
  HS65_LH_AOI22X1 U7854 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][12] ), .B(n8937), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][12] ), .D(
        n9262), .Z(n6692) );
  HS65_LH_AO22X4 U7855 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][12] ), .B(n8940), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][12] ), .D(
        n8949), .Z(n6695) );
  HS65_LH_AOI22X1 U7856 ( .A(n8868), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][12] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][12] ), .D(n9009), 
        .Z(n7142) );
  HS65_LH_AOI22X1 U7857 ( .A(n9161), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][12] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][12] ), .D(n9095), 
        .Z(n7143) );
  HS65_LH_AO22X4 U7858 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][12] ), .B(n9153), 
        .C(n9068), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][12] ), .Z(n7141)
         );
  HS65_LH_AO22X4 U7859 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][12] ), .B(n9165), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][12] ), .D(
        n9065), .Z(n7140) );
  HS65_LH_AOI22X1 U7860 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][12] ), .B(n9098), 
        .C(n9200), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][12] ), .Z(n7139)
         );
  HS65_LH_AOI22X1 U7861 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][12] ), .B(n9062), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][12] ), .D(
        n8863), .Z(n7144) );
  HS65_LH_AOI22X1 U7862 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][12] ), .B(n9159), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][12] ), .D(
        n8862), .Z(n7149) );
  HS65_LH_AOI22X1 U7863 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][7] ), .B(n8937), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][7] ), .D(n9262), .Z(n6466) );
  HS65_LH_AOI22X1 U7864 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][7] ), .B(n8859), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][7] ), .D(
        n9116), .Z(n6460) );
  HS65_LH_AOI22X1 U7865 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][7] ), .B(n8933), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][7] ), .D(
        n9240), .Z(n6470) );
  HS65_LH_AO22X4 U7866 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][7] ), .B(n9260), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][7] ), .D(n9189), .Z(n6473) );
  HS65_LH_AOI22X1 U7867 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][7] ), .B(n9096), 
        .C(n9158), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][7] ), .Z(n6042)
         );
  HS65_LH_AO22X4 U7868 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][7] ), .B(n8947), 
        .C(n8946), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][7] ), .Z(n6041)
         );
  HS65_LH_AO22X4 U7869 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][7] ), .B(n8948), 
        .C(n8951), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][7] ), .Z(n6040)
         );
  HS65_LH_AO22X4 U7870 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][7] ), .B(n9070), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][7] ), .D(
        n9064), .Z(n6054) );
  HS65_LH_AOI22X1 U7871 ( .A(n9243), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][7] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][7] ), .D(n9009), 
        .Z(n6046) );
  HS65_LH_AO22X4 U7872 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][13] ), .B(n9251), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][13] ), .D(
        n9155), .Z(n6407) );
  HS65_LH_AOI22X1 U7873 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][13] ), .B(n9246), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][13] ), .D(
        n9067), .Z(n6405) );
  HS65_LH_AOI22X1 U7874 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][13] ), .B(n8859), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][13] ), .D(
        n9116), .Z(n6399) );
  HS65_LH_AOI22X1 U7875 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][13] ), .B(n9248), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][13] ), .D(
        n9240), .Z(n6409) );
  HS65_LH_AO22X4 U7876 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][13] ), .B(n9160), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][13] ), .D(
        n9267), .Z(n6411) );
  HS65_LH_AO22X4 U7877 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][13] ), .B(n9010), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][13] ), .D(
        n9189), .Z(n6412) );
  HS65_LH_AOI22X1 U7878 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][13] ), .B(n9096), 
        .C(n9158), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][13] ), .Z(n7018)
         );
  HS65_LH_AO22X4 U7879 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][13] ), .B(n8947), 
        .C(n8946), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][13] ), .Z(n7017)
         );
  HS65_LH_AO22X4 U7880 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][13] ), .B(n8948), 
        .C(n8951), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][13] ), .Z(n7016)
         );
  HS65_LH_AO22X4 U7881 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][13] ), .B(n9070), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][13] ), .D(
        n9064), .Z(n7030) );
  HS65_LH_AO22X4 U7882 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][13] ), .B(n9152), 
        .C(n9097), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][13] ), .Z(n7031)
         );
  HS65_LH_AOI22X1 U7883 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][13] ), .B(n9113), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][13] ), .D(
        n8861), .Z(n7028) );
  HS65_LH_AO22X4 U7884 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][13] ), .B(n8867), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][13] ), .D(
        n8866), .Z(n7026) );
  HS65_LH_AO22X4 U7885 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][13] ), .B(n9102), 
        .C(n9101), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][13] ), .Z(n7027)
         );
  HS65_LH_AOI22X1 U7886 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][29] ), .B(n8851), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][29] ), .D(
        n8850), .Z(n6920) );
  HS65_LH_AOI22X1 U7887 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][29] ), .B(n8937), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][29] ), .D(
        n9067), .Z(n6919) );
  HS65_LH_AOI22X1 U7888 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][29] ), .B(n8860), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][29] ), .D(
        n9157), .Z(n6907) );
  HS65_LH_AO22X4 U7889 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][29] ), .B(n8885), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][29] ), .D(
        n8856), .Z(n6904) );
  HS65_LH_AOI22X1 U7890 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][29] ), .B(n8933), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][29] ), .D(
        n9163), .Z(n6923) );
  HS65_LH_AOI22X1 U7891 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][29] ), .B(n8884), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][29] ), .D(
        n8848), .Z(n6924) );
  HS65_LH_AO22X4 U7892 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][29] ), .B(n9260), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][29] ), .D(
        n9189), .Z(n6926) );
  HS65_LH_AOI22X1 U7893 ( .A(n8868), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][29] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][29] ), .D(n9197), 
        .Z(n7556) );
  HS65_LH_AO22X4 U7894 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][29] ), .B(n9152), 
        .C(n9097), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][29] ), .Z(n7559)
         );
  HS65_LH_AOI22X1 U7895 ( .A(n9161), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][29] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][29] ), .D(n9095), 
        .Z(n7557) );
  HS65_LH_AO22X4 U7896 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][29] ), .B(n9166), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[9][29] ), .D(
        n9113), .Z(n7558) );
  HS65_LH_AO22X4 U7897 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][29] ), .B(n9096), 
        .C(n9198), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][29] ), .Z(n7547)
         );
  HS65_LH_AO22X4 U7898 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][29] ), .B(n9165), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][29] ), .D(
        n9065), .Z(n7563) );
  HS65_LH_AO22X4 U7899 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][29] ), .B(n9153), 
        .C(n9068), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][29] ), .Z(n7564)
         );
  HS65_LH_AOI22X1 U7900 ( .A(n9201), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][29] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][29] ), .D(n9202), 
        .Z(n7562) );
  HS65_LH_AOI22X1 U7901 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][21] ), .B(n8859), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][21] ), .D(
        n9116), .Z(n6379) );
  HS65_LH_AOI22X1 U7902 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][21] ), .B(n9226), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][21] ), .D(
        n8848), .Z(n6390) );
  HS65_LH_AO22X4 U7903 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][21] ), .B(n9160), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][21] ), .D(
        n9164), .Z(n6391) );
  HS65_LH_AO22X4 U7904 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][21] ), .B(n9010), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][21] ), .D(
        n8849), .Z(n6392) );
  HS65_LH_AOI22X1 U7905 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][21] ), .B(n9246), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][21] ), .D(
        n9262), .Z(n6385) );
  HS65_LH_AO22X4 U7906 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][21] ), .B(n9251), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][21] ), .D(
        n9155), .Z(n6387) );
  HS65_LH_AOI22X1 U7907 ( .A(n9243), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][21] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][21] ), .D(n9009), 
        .Z(n6000) );
  HS65_LH_AO22X4 U7908 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][21] ), .B(n9165), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][21] ), .D(
        n9065), .Z(n5998) );
  HS65_LH_AOI22X1 U7909 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][21] ), .B(n9096), 
        .C(n9158), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][21] ), .Z(n5996)
         );
  HS65_LH_AO22X4 U7910 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][21] ), .B(n8947), 
        .C(n8946), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][21] ), .Z(n5995)
         );
  HS65_LH_AO22X4 U7911 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][21] ), .B(n8948), 
        .C(n8951), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][21] ), .Z(n5994)
         );
  HS65_LH_AOI22X1 U7912 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][5] ), .B(n9246), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][5] ), .D(n9067), .Z(n6631) );
  HS65_LH_AOI22X1 U7913 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][5] ), .B(n8938), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][5] ), .D(n8850), .Z(n6632) );
  HS65_LH_AOI22X1 U7914 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][5] ), .B(n9226), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][5] ), .D(n8848), .Z(n6637) );
  HS65_LH_AO22X4 U7915 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][5] ), .B(n9160), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][5] ), .D(n9164), .Z(n6638) );
  HS65_LH_AOI22X1 U7916 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][5] ), .B(n9248), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][5] ), .D(
        n9163), .Z(n6636) );
  HS65_LH_AO22X4 U7917 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][5] ), .B(n9010), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][5] ), .D(n8849), .Z(n6639) );
  HS65_LH_AO22X4 U7918 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][5] ), .B(n8885), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][5] ), .D(
        n8856), .Z(n6623) );
  HS65_LH_AOI22X1 U7919 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][5] ), .B(n9098), 
        .C(n9200), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][5] ), .Z(n7079)
         );
  HS65_LH_AO22X4 U7920 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][5] ), .B(n9206), 
        .C(n9205), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][5] ), .Z(n7077)
         );
  HS65_LH_AO22X4 U7921 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][5] ), .B(n9204), 
        .C(n9203), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][5] ), .Z(n7076)
         );
  HS65_LH_AO22X4 U7922 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][5] ), .B(n9165), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][5] ), .D(
        n9065), .Z(n7080) );
  HS65_LH_AO22X4 U7923 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][5] ), .B(n9153), 
        .C(n9068), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][5] ), .Z(n7081)
         );
  HS65_LH_AOI22X1 U7924 ( .A(n9161), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][5] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][5] ), .D(n9095), 
        .Z(n7083) );
  HS65_LH_AOI22X1 U7925 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][25] ), .B(n8860), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][25] ), .D(
        n9157), .Z(n6955) );
  HS65_LH_AO22X4 U7926 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][25] ), .B(n8885), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][25] ), .D(
        n8856), .Z(n6952) );
  HS65_LH_AO22X4 U7927 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][25] ), .B(n9154), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][25] ), .D(
        n8852), .Z(n6956) );
  HS65_LH_AO22X4 U7928 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][25] ), .B(n9156), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][25] ), .D(
        n8853), .Z(n6957) );
  HS65_LH_AOI22X1 U7929 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][25] ), .B(n8933), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][25] ), .D(
        n9163), .Z(n6964) );
  HS65_LH_AO22X4 U7930 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][25] ), .B(n9260), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][25] ), .D(
        n9189), .Z(n6967) );
  HS65_LH_AOI22X1 U7931 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][25] ), .B(n8937), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][25] ), .D(
        n9067), .Z(n6960) );
  HS65_LH_AO22X4 U7932 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][25] ), .B(n8940), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][25] ), .D(
        n8949), .Z(n6963) );
  HS65_LH_AOI22X1 U7933 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][25] ), .B(n9096), 
        .C(n9158), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][25] ), .Z(n7478)
         );
  HS65_LH_AO22X4 U7934 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][25] ), .B(n8947), 
        .C(n8946), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][25] ), .Z(n7477)
         );
  HS65_LH_AO22X4 U7935 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][25] ), .B(n8948), 
        .C(n8951), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][25] ), .Z(n7476)
         );
  HS65_LH_AO22X4 U7936 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][25] ), .B(n9070), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][25] ), .D(
        n9064), .Z(n7490) );
  HS65_LH_AO22X4 U7937 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][25] ), .B(n9152), 
        .C(n9097), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][25] ), .Z(n7491)
         );
  HS65_LH_AO22X4 U7938 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][25] ), .B(n8867), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][25] ), .D(
        n8866), .Z(n7486) );
  HS65_LH_AO22X4 U7939 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][25] ), .B(n9102), 
        .C(n9101), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][25] ), .Z(n7487)
         );
  HS65_LH_AOI22X1 U7940 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][9] ), .B(n8860), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][9] ), .D(
        n9157), .Z(n6981) );
  HS65_LH_AO22X4 U7941 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][9] ), .B(n8885), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][9] ), .D(
        n8856), .Z(n6978) );
  HS65_LH_AO22X4 U7942 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][9] ), .B(n9154), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][9] ), .D(
        n8852), .Z(n6987) );
  HS65_LH_AO22X4 U7943 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][9] ), .B(n9156), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][9] ), .D(
        n8853), .Z(n6988) );
  HS65_LH_AOI22X1 U7944 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][9] ), .B(n8933), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][9] ), .D(
        n9163), .Z(n7004) );
  HS65_LH_AO22X4 U7945 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][9] ), .B(n9260), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][9] ), .D(n9189), .Z(n7007) );
  HS65_LH_AOI22X1 U7946 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][9] ), .B(n8937), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][9] ), .D(n9067), .Z(n6994) );
  HS65_LH_AO22X4 U7947 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][9] ), .B(n8940), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][9] ), .D(
        n8949), .Z(n6997) );
  HS65_LH_AOI22X1 U7948 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][9] ), .B(n9159), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][9] ), .D(n8862), .Z(n7069) );
  HS65_LH_AOI22X1 U7949 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][9] ), .B(n9098), 
        .C(n9200), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][9] ), .Z(n7059)
         );
  HS65_LH_AO22X4 U7950 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][9] ), .B(n9206), 
        .C(n9205), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][9] ), .Z(n7057)
         );
  HS65_LH_AO22X4 U7951 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][9] ), .B(n9204), 
        .C(n9203), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][9] ), .Z(n7056)
         );
  HS65_LH_AOI22X1 U7952 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][9] ), .B(n9062), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][9] ), .D(n8863), .Z(n7064) );
  HS65_LH_AO22X4 U7953 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][9] ), .B(n9165), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][9] ), .D(
        n9065), .Z(n7060) );
  HS65_LH_AO22X4 U7954 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][9] ), .B(n9153), 
        .C(n9068), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][9] ), .Z(n7061)
         );
  HS65_LH_AOI22X1 U7955 ( .A(n9161), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][9] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][9] ), .D(n9095), 
        .Z(n7063) );
  HS65_LH_AO22X4 U7956 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][24] ), .B(n9251), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][24] ), .D(
        n9155), .Z(n6275) );
  HS65_LH_AOI22X1 U7957 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][24] ), .B(n9246), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][24] ), .D(
        n9067), .Z(n6273) );
  HS65_LH_AO22X4 U7958 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][24] ), .B(n9160), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][24] ), .D(
        n9267), .Z(n6281) );
  HS65_LH_AO22X4 U7959 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][24] ), .B(n9010), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][24] ), .D(
        n9189), .Z(n6282) );
  HS65_LH_AO22X4 U7960 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][24] ), .B(n9469), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][24] ), .D(
        n8853), .Z(n6269) );
  HS65_LH_AOI22X1 U7961 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][24] ), .B(n9096), 
        .C(n9158), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][24] ), .Z(n5974)
         );
  HS65_LH_AO22X4 U7962 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][24] ), .B(n8947), 
        .C(n8946), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][24] ), .Z(n5973)
         );
  HS65_LH_AO22X4 U7963 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][24] ), .B(n8948), 
        .C(n8951), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][24] ), .Z(n5972)
         );
  HS65_LH_AOI22X1 U7964 ( .A(n9243), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][24] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][24] ), .D(n9009), 
        .Z(n5978) );
  HS65_LH_AO22X4 U7965 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][28] ), .B(n8885), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][28] ), .D(
        n8856), .Z(n6520) );
  HS65_LH_AOI22X1 U7966 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][28] ), .B(n9246), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][28] ), .D(
        n9067), .Z(n6531) );
  HS65_LH_AOI22X1 U7967 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][28] ), .B(n8938), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][28] ), .D(
        n8850), .Z(n6532) );
  HS65_LH_AO22X4 U7968 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][28] ), .B(n9010), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][28] ), .D(
        n8849), .Z(n6538) );
  HS65_LH_AOI22X1 U7969 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][28] ), .B(n9226), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][28] ), .D(
        n8848), .Z(n6536) );
  HS65_LH_AOI22X1 U7970 ( .A(n9243), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][28] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][28] ), .D(n9009), 
        .Z(n7589) );
  HS65_LH_AO22X4 U7971 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][28] ), .B(n9166), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[9][28] ), .D(
        n9113), .Z(n7591) );
  HS65_LH_AO22X4 U7972 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][28] ), .B(n9165), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][28] ), .D(
        n9065), .Z(n7598) );
  HS65_LH_AO22X4 U7973 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][28] ), .B(n9153), 
        .C(n9068), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][28] ), .Z(n7599)
         );
  HS65_LH_AOI22X1 U7975 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][22] ), .B(n9246), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][22] ), .D(
        n9067), .Z(n6551) );
  HS65_LH_AOI22X1 U7976 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][22] ), .B(n8938), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][22] ), .D(
        n8850), .Z(n6552) );
  HS65_LH_AOI22X1 U7977 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][22] ), .B(n9226), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][22] ), .D(
        n8848), .Z(n6556) );
  HS65_LH_AO22X4 U7978 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][22] ), .B(n9160), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][22] ), .D(
        n9164), .Z(n6557) );
  HS65_LH_AOI22X1 U7979 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][22] ), .B(n9248), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][22] ), .D(
        n9163), .Z(n6555) );
  HS65_LH_AO22X4 U7980 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][22] ), .B(n9010), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][22] ), .D(
        n8849), .Z(n6558) );
  HS65_LH_AO22X4 U7981 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][22] ), .B(n8885), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][22] ), .D(
        n8856), .Z(n6543) );
  HS65_LH_AOI22X1 U7982 ( .A(n9243), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][22] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][22] ), .D(n9197), 
        .Z(n7182) );
  HS65_LH_AOI22X1 U7983 ( .A(n9207), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][22] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][22] ), .D(n9095), 
        .Z(n7183) );
  HS65_LH_AOI22X1 U7984 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][22] ), .B(n9098), 
        .C(n9200), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][22] ), .Z(n7179)
         );
  HS65_LH_AO22X4 U7985 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][22] ), .B(n9206), 
        .C(n9205), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][22] ), .Z(n7177)
         );
  HS65_LH_AO22X4 U7986 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][22] ), .B(n9204), 
        .C(n9203), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][22] ), .Z(n7176)
         );
  HS65_LH_AOI22X1 U7987 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][22] ), .B(n9062), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][22] ), .D(
        n8863), .Z(n7184) );
  HS65_LH_AO22X4 U7988 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][22] ), .B(n9102), 
        .C(n9101), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][22] ), .Z(n7187)
         );
  HS65_LH_AO22X4 U7989 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][22] ), .B(n9070), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][22] ), .D(
        n9244), .Z(n7190) );
  HS65_LH_AOI22X1 U7990 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][22] ), .B(n9250), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][22] ), .D(
        n8862), .Z(n7189) );
  HS65_LH_AOI22X1 U7991 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][4] ), .B(n9246), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][4] ), .D(n9067), .Z(n6425) );
  HS65_LH_AOI22X1 U7992 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][4] ), .B(n8859), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][4] ), .D(
        n9116), .Z(n6419) );
  HS65_LH_AO22X4 U7993 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][4] ), .B(n9010), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][4] ), .D(n8849), .Z(n6432) );
  HS65_LH_AO22X4 U7994 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][4] ), .B(n9160), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][4] ), .D(n9164), .Z(n6431) );
  HS65_LH_AOI22X1 U7995 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][4] ), .B(n9162), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][4] ), .D(
        n8854), .Z(n6423) );
  HS65_LH_AOI22X1 U7996 ( .A(n9243), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][4] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][4] ), .D(n9009), 
        .Z(n6024) );
  HS65_LH_AO22X4 U7997 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][4] ), .B(n9096), 
        .C(n9158), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][4] ), .Z(n6018)
         );
  HS65_LH_AO22X4 U7998 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][4] ), .B(n9098), 
        .C(n9100), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][4] ), .Z(n6019)
         );
  HS65_LH_AO22X4 U7999 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][4] ), .B(n9102), 
        .C(n9101), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][4] ), .Z(n6031) );
  HS65_LH_AO22X4 U8000 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][4] ), .B(n9070), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][4] ), .D(
        n9064), .Z(n6034) );
  HS65_LH_AO22X4 U8001 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][8] ), .B(n9469), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][8] ), .D(
        n8853), .Z(n6649) );
  HS65_LH_AO22X4 U8002 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][8] ), .B(n9154), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][8] ), .D(
        n8852), .Z(n6648) );
  HS65_LH_AOI22X1 U8003 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][8] ), .B(n8933), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][8] ), .D(
        n9240), .Z(n6656) );
  HS65_LH_AO22X4 U8004 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][8] ), .B(n9260), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][8] ), .D(n9189), .Z(n6659) );
  HS65_LH_AOI22X1 U8005 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][8] ), .B(n8937), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][8] ), .D(n9262), .Z(n6652) );
  HS65_LH_AO22X4 U8006 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][8] ), .B(n8940), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][8] ), .D(
        n8949), .Z(n6655) );
  HS65_LH_AOI22X1 U8007 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][8] ), .B(n9159), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][8] ), .D(n8862), .Z(n6854) );
  HS65_LH_AOI22X1 U8008 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][8] ), .B(n9098), 
        .C(n9200), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][8] ), .Z(n6844)
         );
  HS65_LH_AO22X4 U8009 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][8] ), .B(n9206), 
        .C(n9205), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][8] ), .Z(n6842)
         );
  HS65_LH_AO22X4 U8010 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][8] ), .B(n9204), 
        .C(n9203), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][8] ), .Z(n6841)
         );
  HS65_LH_AOI22X1 U8011 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][8] ), .B(n9062), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][8] ), .D(n8863), .Z(n6849) );
  HS65_LH_AO22X4 U8012 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][8] ), .B(n9165), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][8] ), .D(
        n9065), .Z(n6845) );
  HS65_LH_AO22X4 U8013 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][8] ), .B(n9153), 
        .C(n9068), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][8] ), .Z(n6846)
         );
  HS65_LH_AO22X4 U8014 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][20] ), .B(n8885), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][20] ), .D(
        n8856), .Z(n6583) );
  HS65_LH_AOI22X1 U8015 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][20] ), .B(n9226), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][20] ), .D(
        n8848), .Z(n6596) );
  HS65_LH_AO22X4 U8016 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][20] ), .B(n9160), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][20] ), .D(
        n9164), .Z(n6597) );
  HS65_LH_AOI22X1 U8017 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][20] ), .B(n9248), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][20] ), .D(
        n9163), .Z(n6595) );
  HS65_LH_AO22X4 U8018 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][20] ), .B(n9260), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][20] ), .D(
        n8849), .Z(n6598) );
  HS65_LH_AOI22X1 U8019 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][20] ), .B(n8938), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][20] ), .D(
        n8850), .Z(n6592) );
  HS65_LH_AOI22X1 U8020 ( .A(n9243), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][20] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][20] ), .D(n9197), 
        .Z(n7102) );
  HS65_LH_AO22X4 U8021 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][20] ), .B(n9165), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][20] ), .D(
        n9245), .Z(n7100) );
  HS65_LH_AOI22X1 U8022 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][20] ), .B(n9096), 
        .C(n9158), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][20] ), .Z(n7098)
         );
  HS65_LH_AOI22X1 U8023 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][20] ), .B(n9247), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][20] ), .D(
        n8863), .Z(n7104) );
  HS65_LH_AO22X4 U8024 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][20] ), .B(n9102), 
        .C(n9101), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][20] ), .Z(n7107)
         );
  HS65_LH_AOI22X1 U8025 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][20] ), .B(n9113), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][20] ), .D(
        n8861), .Z(n7108) );
  HS65_LH_AOI22X1 U8026 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][20] ), .B(n9159), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][20] ), .D(
        n8862), .Z(n7109) );
  HS65_LH_AO22X4 U8027 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][20] ), .B(n9070), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][20] ), .D(
        n9064), .Z(n7110) );
  HS65_LH_AOI22X1 U8028 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][16] ), .B(n8859), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][16] ), .D(
        n9195), .Z(n6167) );
  HS65_LH_AO22X4 U8029 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][16] ), .B(n9260), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][16] ), .D(
        n8849), .Z(n6192) );
  HS65_LH_AOI22X1 U8030 ( .A(n9243), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][16] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][16] ), .D(n9009), 
        .Z(n6066) );
  HS65_LH_AOI22X1 U8031 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][16] ), .B(n9096), 
        .C(n9158), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][16] ), .Z(n6062)
         );
  HS65_LH_AO22X4 U8032 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][16] ), .B(n8947), 
        .C(n8946), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][16] ), .Z(n6061)
         );
  HS65_LH_AO22X4 U8033 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][16] ), .B(n8948), 
        .C(n8951), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][16] ), .Z(n6060)
         );
  HS65_LH_AOI22X1 U8034 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][17] ), .B(n8859), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][17] ), .D(
        n9116), .Z(n6359) );
  HS65_LH_AOI22X1 U8035 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][17] ), .B(n9226), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][17] ), .D(
        n8848), .Z(n6370) );
  HS65_LH_AO22X4 U8036 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][17] ), .B(n9160), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][17] ), .D(
        n9164), .Z(n6371) );
  HS65_LH_AO22X4 U8037 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][17] ), .B(n9010), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][17] ), .D(
        n8849), .Z(n6372) );
  HS65_LH_AOI22X1 U8038 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][17] ), .B(n9246), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][17] ), .D(
        n9262), .Z(n6365) );
  HS65_LH_AO22X4 U8039 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][17] ), .B(n9251), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][17] ), .D(
        n9155), .Z(n6367) );
  HS65_LH_AO22X4 U8040 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][17] ), .B(n9165), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][17] ), .D(
        n9065), .Z(n5945) );
  HS65_LH_AOI22X1 U8041 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][17] ), .B(n9096), 
        .C(n9158), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][17] ), .Z(n5942)
         );
  HS65_LH_AO22X4 U8042 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][17] ), .B(n8947), 
        .C(n8946), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][17] ), .Z(n5941)
         );
  HS65_LH_AO22X4 U8043 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][17] ), .B(n8948), 
        .C(n8951), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][17] ), .Z(n5940)
         );
  HS65_LH_AOI22X1 U8044 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][2] ), .B(n8859), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][2] ), .D(
        n9195), .Z(n6219) );
  HS65_LH_AOI22X1 U8045 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][2] ), .B(n8851), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][2] ), .D(n8850), .Z(n6226) );
  HS65_LH_AO22X4 U8046 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][2] ), .B(n9010), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][2] ), .D(n8849), .Z(n6232) );
  HS65_LH_AO22X4 U8047 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][2] ), .B(n9160), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][2] ), .D(n9164), .Z(n6231) );
  HS65_LH_AOI22X1 U8048 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][2] ), .B(n9159), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][2] ), .D(n8862), .Z(n6155) );
  HS65_LH_AO22X4 U8049 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][2] ), .B(n9206), 
        .C(n9205), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][2] ), .Z(n6143)
         );
  HS65_LH_AO22X4 U8050 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][2] ), .B(n9204), 
        .C(n9203), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][2] ), .Z(n6142)
         );
  HS65_LH_AOI22X1 U8051 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][2] ), .B(n9062), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][2] ), .D(n8863), .Z(n6150) );
  HS65_LH_AO22X4 U8052 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][18] ), .B(n9154), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][18] ), .D(
        n8852), .Z(n6668) );
  HS65_LH_AO22X4 U8053 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][18] ), .B(n9156), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][18] ), .D(
        n8853), .Z(n6669) );
  HS65_LH_AOI22X1 U8054 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][18] ), .B(n8933), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][18] ), .D(
        n9240), .Z(n6676) );
  HS65_LH_AO22X4 U8055 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][18] ), .B(n9260), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][18] ), .D(
        n9189), .Z(n6679) );
  HS65_LH_AOI22X1 U8056 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][18] ), .B(n8937), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][18] ), .D(
        n9262), .Z(n6672) );
  HS65_LH_AO22X4 U8057 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][18] ), .B(n8940), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][18] ), .D(
        n8949), .Z(n6675) );
  HS65_LH_AO22X4 U8058 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][18] ), .B(n8947), 
        .C(n8946), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][18] ), .Z(n7219)
         );
  HS65_LH_AO22X4 U8059 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][18] ), .B(n8948), 
        .C(n8951), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][18] ), .Z(n7218)
         );
  HS65_LH_AO22X4 U8060 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][18] ), .B(n9070), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][18] ), .D(
        n9064), .Z(n7232) );
  HS65_LH_AO22X4 U8061 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][18] ), .B(n9152), 
        .C(n9097), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][18] ), .Z(n7233)
         );
  HS65_LH_AO22X4 U8062 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][18] ), .B(n8867), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][18] ), .D(
        n8866), .Z(n7228) );
  HS65_LH_AO22X4 U8063 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][18] ), .B(n9102), 
        .C(n9101), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][18] ), .Z(n7229)
         );
  HS65_LH_AO22X4 U8064 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][6] ), .B(n9154), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][6] ), .D(
        n8852), .Z(n6732) );
  HS65_LH_AO22X4 U8065 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][6] ), .B(n9156), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][6] ), .D(
        n8853), .Z(n6733) );
  HS65_LH_AOI22X1 U8066 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][6] ), .B(n8933), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][6] ), .D(
        n9240), .Z(n6740) );
  HS65_LH_AO22X4 U8067 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][6] ), .B(n9260), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][6] ), .D(n9189), .Z(n6743) );
  HS65_LH_AOI22X1 U8068 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][6] ), .B(n8937), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][6] ), .D(n9262), .Z(n6736) );
  HS65_LH_AO22X4 U8069 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][6] ), .B(n8940), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][6] ), .D(
        n8949), .Z(n6739) );
  HS65_LH_AOI22X1 U8070 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][6] ), .B(n9159), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][6] ), .D(n8862), .Z(n6834) );
  HS65_LH_AOI22X1 U8071 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][6] ), .B(n9098), 
        .C(n9200), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][6] ), .Z(n6824)
         );
  HS65_LH_AO22X4 U8072 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][6] ), .B(n9206), 
        .C(n9205), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][6] ), .Z(n6822)
         );
  HS65_LH_AO22X4 U8073 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][6] ), .B(n9204), 
        .C(n9203), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][6] ), .Z(n6821)
         );
  HS65_LH_AOI22X1 U8074 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][6] ), .B(n9062), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][6] ), .D(n8863), .Z(n6829) );
  HS65_LH_AO22X4 U8075 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][6] ), .B(n9165), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][6] ), .D(
        n9065), .Z(n6825) );
  HS65_LH_AO22X4 U8076 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][6] ), .B(n9153), 
        .C(n9068), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][6] ), .Z(n6826)
         );
  HS65_LH_AO22X4 U8077 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][1] ), .B(n9251), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][1] ), .D(
        n9155), .Z(n6248) );
  HS65_LH_AOI22X1 U8078 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][1] ), .B(n9246), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][1] ), .D(n9262), .Z(n6246) );
  HS65_LH_AO22X4 U8079 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][1] ), .B(n8859), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][1] ), .D(
        n9195), .Z(n6237) );
  HS65_LH_AO22X4 U8080 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][1] ), .B(n9010), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][1] ), .D(n8849), .Z(n6253) );
  HS65_LH_AOI22X1 U8081 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][1] ), .B(n9248), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][1] ), .D(
        n9240), .Z(n6250) );
  HS65_LH_AO22X4 U8082 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][1] ), .B(n9160), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][1] ), .D(n9164), .Z(n6252) );
  HS65_LH_AO22X4 U8083 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][1] ), .B(n9070), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][1] ), .D(
        n9064), .Z(n7252) );
  HS65_LH_AO22X4 U8084 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][1] ), .B(n9152), 
        .C(n9097), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][1] ), .Z(n7253) );
  HS65_LH_AO22X4 U8085 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][1] ), .B(n8867), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][1] ), .D(
        n8866), .Z(n7248) );
  HS65_LH_AO22X4 U8086 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][1] ), .B(n9102), 
        .C(n9101), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][1] ), .Z(n7249) );
  HS65_LH_AOI22X1 U8087 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][0] ), .B(n8859), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][0] ), .D(
        n9195), .Z(n6199) );
  HS65_LH_AO22X4 U8088 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][0] ), .B(n9260), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][0] ), .D(n8849), .Z(n6212) );
  HS65_LH_AO22X4 U8094 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][0] ), .B(n9165), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][0] ), .D(
        n9065), .Z(n7285) );
  HS65_LH_AO22X4 U8095 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][0] ), .B(n9153), 
        .C(n9068), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][0] ), .Z(n7286)
         );
  HS65_LH_AOI22X1 U8097 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][31] ), .B(n9246), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][31] ), .D(
        n9067), .Z(n6611) );
  HS65_LH_AOI22X1 U8098 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][31] ), .B(n8938), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][31] ), .D(
        n8850), .Z(n6612) );
  HS65_LH_AOI22X1 U8099 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][31] ), .B(n9226), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][31] ), .D(
        n8848), .Z(n6616) );
  HS65_LH_AO22X4 U8100 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][31] ), .B(n9160), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][31] ), .D(
        n9164), .Z(n6617) );
  HS65_LH_AOI22X1 U8101 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][31] ), .B(n9248), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][31] ), .D(
        n9163), .Z(n6615) );
  HS65_LH_AO22X4 U8102 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][31] ), .B(n9010), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][31] ), .D(
        n8849), .Z(n6618) );
  HS65_LH_AO22X4 U8103 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][31] ), .B(n8885), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][31] ), .D(
        n8856), .Z(n6603) );
  HS65_LH_BFX9 U8104 ( .A(n8368), .Z(n7716) );
  HS65_LH_CNIVX3 U8105 ( .A(n5629), .Z(n5630) );
  HS65_LH_CNIVX3 U8106 ( .A(n5589), .Z(n5590) );
  HS65_LH_CNIVX3 U8107 ( .A(n5688), .Z(n5689) );
  HS65_LH_CNIVX3 U8108 ( .A(n5695), .Z(n5696) );
  HS65_LH_CNIVX3 U8109 ( .A(n5650), .Z(n5651) );
  HS65_LH_NOR2AX3 U8113 ( .A(n5041), .B(n5040), .Z(n5042) );
  HS65_LH_CNIVX3 U8114 ( .A(n5349), .Z(n5406) );
  HS65_LH_OR2X4 U8115 ( .A(n5312), .B(n5311), .Z(n2856) );
  HS65_LH_AOI21X2 U8117 ( .A(n5417), .B(n5416), .C(n5415), .Z(n5419) );
  HS65_LH_OAI21X2 U8119 ( .A(n5111), .B(n5110), .C(n5109), .Z(n5112) );
  HS65_LH_AOI21X2 U8125 ( .A(n5095), .B(n5094), .C(n5093), .Z(n5096) );
  HS65_LH_OAI21X2 U8126 ( .A(n4767), .B(n5097), .C(n3842), .Z(n5098) );
  HS65_LH_NOR2X2 U8127 ( .A(n5091), .B(n5097), .Z(n5100) );
  HS65_LH_NOR2X2 U8128 ( .A(\lte_x_57/B[3] ), .B(n2789), .Z(n5091) );
  HS65_LH_OAI21X2 U8130 ( .A(n3767), .B(n4859), .C(n4861), .Z(n5102) );
  HS65_LH_NOR2X2 U8131 ( .A(n5088), .B(n4270), .Z(n5103) );
  HS65_LH_NOR2X2 U8132 ( .A(\lte_x_57/B[7] ), .B(n5207), .Z(n5088) );
  HS65_LL_NOR2X2 U8133 ( .A(n5218), .B(n4859), .Z(n5090) );
  HS65_LH_NOR2X2 U8135 ( .A(n5078), .B(n5110), .Z(n5114) );
  HS65_LH_OAI21X2 U8141 ( .A(n5127), .B(n5184), .C(n5433), .Z(n5128) );
  HS65_LH_NOR3AX2 U8148 ( .A(n4967), .B(n4966), .C(n4965), .Z(n4968) );
  HS65_LH_NAND3X2 U8156 ( .A(n4910), .B(n5187), .C(n5125), .Z(n4911) );
  HS65_LH_IVX2 U8157 ( .A(n5286), .Z(n4922) );
  HS65_LH_NAND3X2 U8158 ( .A(n5311), .B(n5446), .C(n5312), .Z(n4926) );
  HS65_LH_AOI21X2 U8160 ( .A(n5036), .B(n5333), .C(n5336), .Z(n3952) );
  HS65_LH_NAND2X2 U8161 ( .A(n2774), .B(n5508), .Z(n5040) );
  HS65_LH_NAND2X2 U8162 ( .A(n9538), .B(n4871), .Z(n3941) );
  HS65_LH_NAND2X2 U8163 ( .A(n3090), .B(n8721), .Z(n3091) );
  HS65_LH_AOI21X2 U8170 ( .A(n5396), .B(n5027), .C(n5395), .Z(n5397) );
  HS65_LH_AOI22X1 U8172 ( .A(n5386), .B(n5385), .C(n5426), .D(n5384), .Z(n5389) );
  HS65_LH_NAND2X2 U8173 ( .A(\u_DataPath/cw_to_ex_i [0]), .B(n5446), .Z(n5447)
         );
  HS65_LH_OAI22X1 U8174 ( .A(\lte_x_57/B[30] ), .B(n2790), .C(n5445), .D(n5444), .Z(n5448) );
  HS65_LH_AOI21X2 U8175 ( .A(n5337), .B(n5336), .C(n5335), .Z(n5338) );
  HS65_LH_AOI21X2 U8179 ( .A(n5292), .B(n5291), .C(n5290), .Z(n5308) );
  HS65_LH_NAND2X2 U8180 ( .A(n5298), .B(n5297), .Z(n5300) );
  HS65_LH_AOI21X2 U8181 ( .A(n5329), .B(n5328), .C(n5161), .Z(n5171) );
  HS65_LH_OAI21X2 U8182 ( .A(n5288), .B(n5294), .C(n5295), .Z(n5465) );
  HS65_LH_AOI21X2 U8184 ( .A(n5427), .B(n5026), .C(n5025), .Z(n5034) );
  HS65_LH_AOI21X2 U8185 ( .A(n5032), .B(n5394), .C(n5031), .Z(n5033) );
  HS65_LH_AOI312X2 U8187 ( .A(n5450), .B(n5315), .C(n5019), .D(n5453), .E(
        n5438), .F(n5018), .Z(n5020) );
  HS65_LH_NAND3X2 U8188 ( .A(n5072), .B(n5016), .C(n4594), .Z(n5019) );
  HS65_LH_CBI4I6X2 U8189 ( .A(n5445), .B(n5444), .C(n5309), .D(n5014), .Z(
        n5022) );
  HS65_LH_OAI21X2 U8190 ( .A(n5450), .B(n5317), .C(n5455), .Z(n4934) );
  HS65_LL_OAI13X1 U8192 ( .A(n5192), .B(n5316), .C(n3200), .D(n5452), .Z(n4936) );
  HS65_LH_OA112X4 U8193 ( .A(n4918), .B(n5066), .C(n2824), .D(n5064), .Z(n4921) );
  HS65_LH_AOI21X2 U8194 ( .A(n4930), .B(n4929), .C(n4928), .Z(n4938) );
  HS65_LH_NAND3X2 U8196 ( .A(n4927), .B(n5449), .C(n4926), .Z(n4928) );
  HS65_LH_NAND3X2 U8198 ( .A(n5192), .B(n5452), .C(n3200), .Z(n4004) );
  HS65_LH_AOI21X2 U8200 ( .A(n5288), .B(n5364), .C(n5296), .Z(n3996) );
  HS65_LH_AOI21X2 U8202 ( .A(n5356), .B(n5335), .C(n5424), .Z(n3971) );
  HS65_LHS_XNOR2X3 U8203 ( .A(n5211), .B(\lte_x_57/B[3] ), .Z(n4972) );
  HS65_LHS_XNOR2X3 U8204 ( .A(n5386), .B(n5385), .Z(n4974) );
  HS65_LLS_XOR2X3 U8205 ( .A(\add_x_50/A[23] ), .B(n5252), .Z(n4961) );
  HS65_LH_CBI4I1X3 U8206 ( .A(n2802), .B(n5203), .C(n4149), .D(n2793), .Z(
        n4152) );
  HS65_LH_OAI21X3 U8207 ( .A(n5529), .B(n2829), .C(n3627), .Z(n3924) );
  HS65_LH_CBI4I1X3 U8213 ( .A(n5507), .B(n5064), .C(n5506), .D(
        \sub_x_51/A[20] ), .Z(n3468) );
  HS65_LH_OAI21X2 U8218 ( .A(n4203), .B(n2829), .C(n4202), .Z(n4207) );
  HS65_LH_OAI22X1 U8219 ( .A(n3054), .B(n3322), .C(n5385), .D(n2829), .Z(n3738) );
  HS65_LH_OAI21X2 U8226 ( .A(n5078), .B(n5426), .C(n5228), .Z(n5229) );
  HS65_LH_OAI21X2 U8227 ( .A(n5233), .B(n5391), .C(n5232), .Z(n5236) );
  HS65_LL_NOR2X2 U8229 ( .A(n4270), .B(n5080), .Z(n5202) );
  HS65_LH_NOR2X2 U8230 ( .A(n5204), .B(n5391), .Z(n5205) );
  HS65_LH_OAI21X2 U8232 ( .A(n5213), .B(n3779), .C(n3777), .Z(n5216) );
  HS65_LH_NAND2X2 U8233 ( .A(n5223), .B(n5210), .Z(n5226) );
  HS65_LH_NOR2X2 U8234 ( .A(n5218), .B(n5209), .Z(n5210) );
  HS65_LL_AND2X4 U8237 ( .A(n5486), .B(n5485), .Z(n5521) );
  HS65_LL_NOR2AX3 U8239 ( .A(n5383), .B(n5382), .Z(n5476) );
  HS65_LH_CBI4I1X3 U8241 ( .A(n5052), .B(n5465), .C(n5463), .D(n5461), .Z(
        n5013) );
  HS65_LH_AOI21X2 U8242 ( .A(n5259), .B(n4004), .C(n4003), .Z(n4007) );
  HS65_LH_OAI21X2 U8243 ( .A(n5297), .B(n3991), .C(n5255), .Z(n4001) );
  HS65_LH_AOI21X2 U8245 ( .A(n5354), .B(n5375), .C(n5372), .Z(n3970) );
  HS65_LH_NOR2X2 U8246 ( .A(\u_DataPath/cw_to_ex_i [2]), .B(n5062), .Z(n4019)
         );
  HS65_LH_NOR2X2 U8247 ( .A(\u_DataPath/cw_to_ex_i [3]), .B(n4018), .Z(n5327)
         );
  HS65_LH_AOI21X2 U8248 ( .A(n5778), .B(n5743), .C(n5742), .Z(n5744) );
  HS65_LHS_XNOR2X3 U8252 ( .A(n5392), .B(n5393), .Z(n3579) );
  HS65_LH_AOI21X2 U8258 ( .A(n4323), .B(n4322), .C(n4792), .Z(n3930) );
  HS65_LHS_XNOR2X3 U8260 ( .A(n5084), .B(n3962), .Z(n4962) );
  HS65_LH_AOI21X2 U8262 ( .A(n3916), .B(n3915), .C(n4659), .Z(n3921) );
  HS65_LH_AOI21X2 U8263 ( .A(n4324), .B(n4325), .C(n4292), .Z(n3922) );
  HS65_LH_NOR2AX3 U8264 ( .A(n3465), .B(n4971), .Z(n3699) );
  HS65_LH_NAND2X2 U8266 ( .A(n4257), .B(n4259), .Z(n3679) );
  HS65_LH_AOI21X2 U8268 ( .A(\lte_x_57/B[10] ), .B(n4247), .C(n4246), .Z(n4248) );
  HS65_LL_OAI22X1 U8269 ( .A(n4846), .B(n3074), .C(n4784), .D(n4284), .Z(n4246) );
  HS65_LH_OAI21X2 U8270 ( .A(n4794), .B(n3074), .C(n3379), .Z(n4247) );
  HS65_LLS_XNOR2X3 U8271 ( .A(\u_DataPath/u_execute/A_inALU_i[26] ), .B(n5190), 
        .Z(n4967) );
  HS65_LH_CBI4I1X3 U8274 ( .A(n5507), .B(n5312), .C(n4500), .D(
        \lte_x_57/B[30] ), .Z(n3300) );
  HS65_LH_AOI21X2 U8275 ( .A(n4781), .B(n5312), .C(n4502), .Z(n3291) );
  HS65_LH_OAI21X2 U8276 ( .A(n4113), .B(n4112), .C(n4743), .Z(n3290) );
  HS65_LH_CBI4I1X3 U8281 ( .A(n5507), .B(n5082), .C(n5506), .D(
        \sub_x_51/A[13] ), .Z(n4060) );
  HS65_LL_NOR2AX3 U8283 ( .A(n4528), .B(n4527), .Z(n4529) );
  HS65_LH_AOI22X1 U8286 ( .A(n4671), .B(n4063), .C(n4842), .D(n3390), .Z(n4065) );
  HS65_LH_AOI22X1 U8291 ( .A(n4673), .B(n4478), .C(n4225), .D(n4477), .Z(n4483) );
  HS65_LH_AOI21X2 U8292 ( .A(n3128), .B(n3826), .C(n3724), .Z(n3725) );
  HS65_LH_NOR2X2 U8293 ( .A(n2824), .B(n3338), .Z(n3723) );
  HS65_LH_AOI21X2 U8297 ( .A(n4781), .B(n5079), .C(n4028), .Z(n4029) );
  HS65_LH_NAND2X2 U8299 ( .A(n2802), .B(n5079), .Z(n4027) );
  HS65_LH_AOI222X2 U8300 ( .A(n4573), .B(n4673), .C(\u_DataPath/cw_to_ex_i [0]), .D(n4619), .E(n4572), .F(n4225), .Z(n4574) );
  HS65_LH_CNIVX3 U8303 ( .A(n3827), .Z(n3828) );
  HS65_LL_NOR2X3 U8307 ( .A(n5184), .B(n4458), .Z(n4704) );
  HS65_LLS_XNOR2X3 U8308 ( .A(n2825), .B(n5251), .Z(n4986) );
  HS65_LH_CBI4I1X3 U8309 ( .A(n5507), .B(n5251), .C(n4149), .D(
        \sub_x_51/A[22] ), .Z(n4130) );
  HS65_LH_AOI21X2 U8310 ( .A(n5517), .B(n4987), .C(n3858), .Z(n3870) );
  HS65_LH_CBI4I1X3 U8316 ( .A(n5507), .B(n5187), .C(n5506), .D(n3128), .Z(
        n4435) );
  HS65_LH_AOI21X2 U8318 ( .A(n5092), .B(n4194), .C(n4193), .Z(n4195) );
  HS65_LH_NOR2X2 U8319 ( .A(n4794), .B(n4192), .Z(n4194) );
  HS65_LL_AOI22X1 U8323 ( .A(n4829), .B(n4828), .C(n5510), .D(n4827), .Z(n4835) );
  HS65_LH_NAND2X2 U8324 ( .A(n4832), .B(n5505), .Z(n4833) );
  HS65_LL_NAND2X2 U8325 ( .A(n4831), .B(n4830), .Z(n4834) );
  HS65_LL_CBI4I1X3 U8326 ( .A(n5507), .B(n5089), .C(n5506), .D(\lte_x_57/B[6] ), .Z(n4845) );
  HS65_LH_NAND2X2 U8329 ( .A(n2802), .B(n7321), .Z(n4652) );
  HS65_LLS_XNOR2X3 U8332 ( .A(\u_DataPath/RFaddr_out_memwb_i [1]), .B(
        \u_DataPath/rs_ex_i [1]), .Z(n2878) );
  HS65_LLS_XNOR2X3 U8333 ( .A(\u_DataPath/rs_ex_i [3]), .B(
        \u_DataPath/RFaddr_out_memwb_i [3]), .Z(n2879) );
  HS65_LH_AOI21X2 U8334 ( .A(n5507), .B(n9538), .C(n4149), .Z(n3805) );
  HS65_LH_OAI21X2 U8335 ( .A(n2829), .B(n4192), .C(n3807), .Z(n3808) );
  HS65_LH_NOR2X2 U8337 ( .A(n4427), .B(n5245), .Z(n5188) );
  HS65_LH_CNIVX3 U8338 ( .A(n7647), .Z(n7015) );
  HS65_LHS_XNOR2X3 U8343 ( .A(\add_x_50/A[19] ), .B(n5246), .Z(n4951) );
  HS65_LH_OA12X4 U8345 ( .A(n4798), .B(n5481), .C(n4797), .Z(n4809) );
  HS65_LL_NOR4ABX2 U8347 ( .A(n4252), .B(n4251), .C(n4250), .D(n4249), .Z(
        n4256) );
  HS65_LLS_XNOR2X3 U8348 ( .A(n4608), .B(n4607), .Z(n4633) );
  HS65_LL_CBI4I1X3 U8349 ( .A(n2802), .B(n5190), .C(n5506), .D(
        \u_DataPath/u_execute/A_inALU_i[26] ), .Z(n4612) );
  HS65_LL_NOR4ABX2 U8351 ( .A(n4757), .B(n4756), .C(n4755), .D(n4754), .Z(
        n4758) );
  HS65_LH_AOI21X2 U8352 ( .A(n5517), .B(n4956), .C(n4158), .Z(n4164) );
  HS65_LH_AOI21X2 U8353 ( .A(n4411), .B(n4162), .C(n4161), .Z(n4163) );
  HS65_LHS_XOR2X3 U8355 ( .A(n4344), .B(n4343), .Z(n4345) );
  HS65_LL_NAND2AX4 U8356 ( .A(n3589), .B(n3588), .Z(n4812) );
  HS65_LH_NOR2X6 U8359 ( .A(n6184), .B(n6183), .Z(n7003) );
  HS65_LLS_XNOR2X3 U8362 ( .A(n3424), .B(n3423), .Z(n3425) );
  HS65_LH_IVX4 U8363 ( .A(n4146), .Z(n3837) );
  HS65_LL_AOI22X1 U8364 ( .A(n4673), .B(n4569), .C(n4842), .D(n4570), .Z(n3831) );
  HS65_LH_NAND2X2 U8367 ( .A(n4673), .B(n4849), .Z(n4121) );
  HS65_LL_NOR3AX2 U8371 ( .A(n3481), .B(n3480), .C(n3479), .Z(n3498) );
  HS65_LH_NOR3AX2 U8372 ( .A(n4438), .B(n4437), .C(n4436), .Z(n4439) );
  HS65_LHS_XOR2X3 U8374 ( .A(n8797), .B(n9316), .Z(n6492) );
  HS65_LL_NAND2X2 U8375 ( .A(n7669), .B(n8325), .Z(n7668) );
  HS65_LH_NAND3X2 U8376 ( .A(n3527), .B(n7216), .C(n7647), .Z(n7643) );
  HS65_LH_NAND3X2 U8377 ( .A(n9334), .B(n9209), .C(n9172), .Z(n7644) );
  HS65_LH_NAND3X2 U8378 ( .A(n9210), .B(n9335), .C(n9172), .Z(n8010) );
  HS65_LH_CNIVX3 U8379 ( .A(n5903), .Z(n5846) );
  HS65_LH_CNIVX3 U8381 ( .A(n5890), .Z(n5891) );
  HS65_LH_CNIVX3 U8383 ( .A(n5851), .Z(n5852) );
  HS65_LH_CNIVX3 U8384 ( .A(n5760), .Z(n5761) );
  HS65_LH_CNIVX3 U8385 ( .A(n5770), .Z(n5771) );
  HS65_LH_CNIVX3 U8387 ( .A(\u_DataPath/pc_4_to_ex_i [19]), .Z(n7444) );
  HS65_LH_CNIVX3 U8388 ( .A(n5910), .Z(n5911) );
  HS65_LLS_XNOR2X3 U8389 ( .A(n4465), .B(n4464), .Z(n4499) );
  HS65_LH_CNIVX3 U8390 ( .A(\u_DataPath/pc_4_to_ex_i [24]), .Z(n6759) );
  HS65_LL_NAND2X2 U8391 ( .A(n3834), .B(n4410), .Z(n3840) );
  HS65_LH_CNIVX3 U8394 ( .A(\u_DataPath/data_read_ex_2_i [0]), .Z(n2956) );
  HS65_LH_CNIVX3 U8395 ( .A(n7351), .Z(n7354) );
  HS65_LH_CBI4I1X3 U8396 ( .A(n7607), .B(n7411), .C(n7410), .D(n7409), .Z(
        n7958) );
  HS65_LH_AOI22X1 U8397 ( .A(n9243), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][31] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][31] ), .D(n9009), 
        .Z(n7511) );
  HS65_LH_AO22X4 U8398 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][31] ), .B(n9152), 
        .C(n9097), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][31] ), .Z(n7514)
         );
  HS65_LH_AO22X4 U8399 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][31] ), .B(n9166), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[9][31] ), .D(
        n9113), .Z(n7513) );
  HS65_LH_AO22X4 U8400 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][31] ), .B(n9098), 
        .C(n9100), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][31] ), .Z(n7497)
         );
  HS65_LH_AO22X4 U8401 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][31] ), .B(n9070), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][31] ), .D(
        n9064), .Z(n7504) );
  HS65_LH_AO22X4 U8402 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][31] ), .B(n9102), 
        .C(n9101), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][31] ), .Z(n7505)
         );
  HS65_LH_NAND3X2 U8403 ( .A(n8021), .B(n7402), .C(n7401), .Z(n8022) );
  HS65_LH_AOI21X2 U8404 ( .A(n8019), .B(n7403), .C(n7405), .Z(n7402) );
  HS65_LH_OR2X4 U8405 ( .A(n8515), .B(\u_DataPath/pc_4_to_ex_i [31]), .Z(n5732) );
  HS65_LH_IVX9 U8406 ( .A(\u_DataPath/jaddr_i [24]), .Z(n8015) );
  HS65_LHS_XOR2X6 U8407 ( .A(n7469), .B(n7468), .Z(\u_DataPath/pc_4_i [23]) );
  HS65_LH_OAI12X3 U8408 ( .A(n9104), .B(n7311), .C(n8787), .Z(n8459) );
  HS65_LH_CNIVX3 U8410 ( .A(n5600), .Z(n5601) );
  HS65_LH_CNIVX3 U8411 ( .A(n5707), .Z(n5708) );
  HS65_LL_OR2ABX27 U8413 ( .A(n9241), .B(n3450), .Z(write_op) );
  HS65_LH_CNIVX3 U8414 ( .A(n8459), .Z(n8460) );
  HS65_LH_CNIVX3 U8415 ( .A(\u_DataPath/RFaddr_out_memwb_i [0]), .Z(n8026) );
  HS65_LH_NAND2AX4 U8416 ( .A(iram_data[28]), .B(n7706), .Z(opcode_i[2]) );
  HS65_LH_NAND2AX4 U8417 ( .A(iram_data[26]), .B(n7705), .Z(opcode_i[0]) );
  HS65_LH_CNIVX3 U8418 ( .A(\u_DataPath/RFaddr_out_memwb_i [1]), .Z(n7937) );
  HS65_LH_CNIVX3 U8419 ( .A(\u_DataPath/RFaddr_out_memwb_i [2]), .Z(n7940) );
  HS65_LH_AO222X4 U8420 ( .A(n7706), .B(n9019), .C(n7690), .D(n8613), .E(n9319), .F(n7686), .Z(addr_to_iram_14) );
  HS65_LH_NAND2AX4 U8421 ( .A(n7712), .B(n9344), .Z(n8126) );
  HS65_LH_NAND2AX4 U8422 ( .A(n7712), .B(n8788), .Z(n8117) );
  HS65_LH_NAND2X2 U8423 ( .A(n1885), .B(n9313), .Z(n8366) );
  HS65_LH_OAI12X24 U8424 ( .A(n8004), .B(n8726), .C(n1885), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N149 ) );
  HS65_LH_OAI12X24 U8425 ( .A(n8004), .B(n8720), .C(n1885), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N148 ) );
  HS65_LL_OAI21X12 U8426 ( .A(n8005), .B(n2720), .C(n1885), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N143 ) );
  HS65_LL_OAI21X12 U8427 ( .A(n8010), .B(n8014), .C(n1885), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N127 ) );
  HS65_LH_OAI12X24 U8428 ( .A(n8004), .B(n3532), .C(n1885), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N152 ) );
  HS65_LL_OAI21X12 U8429 ( .A(n8720), .B(n8014), .C(n1885), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N92 ) );
  HS65_LH_NOR4ABX4 U8430 ( .A(n7987), .B(n8513), .C(n9090), .D(n8901), .Z(
        n7988) );
  HS65_LH_CBI4I1X3 U8431 ( .A(n7613), .B(n7967), .C(opcode_i[0]), .D(n7396), 
        .Z(n7970) );
  HS65_LHS_XOR2X3 U8432 ( .A(n8907), .B(n5902), .Z(
        \u_DataPath/u_execute/resAdd1_i [6]) );
  HS65_LHS_XOR2X3 U8433 ( .A(n8905), .B(n5878), .Z(
        \u_DataPath/u_execute/resAdd1_i [18]) );
  HS65_LHS_XOR2X3 U8434 ( .A(n8904), .B(n5837), .Z(
        \u_DataPath/u_execute/resAdd1_i [17]) );
  HS65_LHS_XOR2X3 U8435 ( .A(n8903), .B(n5830), .Z(
        \u_DataPath/u_execute/resAdd1_i [20]) );
  HS65_LHS_XOR2X3 U8436 ( .A(n8902), .B(n5894), .Z(
        \u_DataPath/u_execute/resAdd1_i [8]) );
  HS65_LH_NAND2X2 U8437 ( .A(n5931), .B(n5930), .Z(n5933) );
  HS65_LHS_XOR2X3 U8439 ( .A(n8916), .B(n5856), .Z(
        \u_DataPath/u_execute/resAdd1_i [5]) );
  HS65_LHS_XOR2X3 U8440 ( .A(n9039), .B(n5821), .Z(
        \u_DataPath/u_execute/resAdd1_i [21]) );
  HS65_LHS_XOR2X3 U8441 ( .A(n8914), .B(n5815), .Z(
        \u_DataPath/u_execute/resAdd1_i [13]) );
  HS65_LH_AOI21X2 U8442 ( .A(n2797), .B(n9332), .C(n8408), .Z(
        \u_DataPath/mem_writedata_out_i [12]) );
  HS65_LH_NAND2X2 U8443 ( .A(n5919), .B(n5918), .Z(n5921) );
  HS65_LHS_XNOR2X3 U8444 ( .A(n8910), .B(n5888), .Z(
        \u_DataPath/u_execute/resAdd1_i [10]) );
  HS65_LHS_XOR2X3 U8445 ( .A(n8909), .B(n5806), .Z(
        \u_DataPath/u_execute/resAdd1_i [11]) );
  HS65_LH_NOR4ABX2 U8446 ( .A(n6328), .B(n6327), .C(n6326), .D(n6325), .Z(
        n8207) );
  HS65_LH_AOI22X1 U8447 ( .A(n8313), .B(n9436), .C(n7693), .D(
        \u_DataPath/u_execute/link_value_i [27]), .Z(n8206) );
  HS65_LH_NOR4ABX2 U8448 ( .A(n6099), .B(n6098), .C(n6097), .D(n6096), .Z(
        n8060) );
  HS65_LH_NOR4ABX2 U8449 ( .A(n6519), .B(n6518), .C(n6517), .D(n6516), .Z(
        n8217) );
  HS65_LH_CNIVX3 U8451 ( .A(\u_DataPath/pc_4_to_ex_i [11]), .Z(n7626) );
  HS65_LH_NOR4ABX2 U8452 ( .A(n6307), .B(n6306), .C(n6305), .D(n6304), .Z(
        n8198) );
  HS65_LH_AOI22X1 U8453 ( .A(n8313), .B(n9134), .C(n7693), .D(
        \u_DataPath/u_execute/link_value_i [19]), .Z(n8195) );
  HS65_LH_NOR4ABX2 U8454 ( .A(n6456), .B(n6455), .C(n6454), .D(n6453), .Z(
        n8057) );
  HS65_LH_NOR4ABX2 U8455 ( .A(n6141), .B(n6140), .C(n6139), .D(n6138), .Z(
        n8297) );
  HS65_LH_CNIVX3 U8456 ( .A(\u_DataPath/pc_4_to_ex_i [3]), .Z(n7420) );
  HS65_LH_NOR4ABX2 U8457 ( .A(n6723), .B(n6722), .C(n6721), .D(n6720), .Z(
        n8235) );
  HS65_LH_CNIVX3 U8458 ( .A(\u_DataPath/pc_4_to_ex_i [10]), .Z(n7427) );
  HS65_LL_AOI22X1 U8459 ( .A(n8687), .B(n9432), .C(n9252), .D(n9105), .Z(n8249) );
  HS65_LH_CNIVX3 U8460 ( .A(\u_DataPath/pc_4_to_ex_i [26]), .Z(n7304) );
  HS65_LH_NOR4ABX2 U8461 ( .A(n6356), .B(n6355), .C(n6354), .D(n6353), .Z(
        n8211) );
  HS65_LH_AOI22X1 U8462 ( .A(n8313), .B(n9428), .C(n7693), .D(
        \u_DataPath/u_execute/link_value_i [23]), .Z(n8210) );
  HS65_LH_NOR4ABX2 U8463 ( .A(n6582), .B(n6581), .C(n6580), .D(n6579), .Z(
        n8289) );
  HS65_LH_NOR4ABX2 U8464 ( .A(n6703), .B(n6702), .C(n6701), .D(n6700), .Z(
        n8240) );
  HS65_LH_NOR4ABX2 U8465 ( .A(n6477), .B(n6476), .C(n6475), .D(n6474), .Z(
        n8225) );
  HS65_LH_NOR4ABX2 U8466 ( .A(n6059), .B(n6058), .C(n6057), .D(n6056), .Z(
        n8064) );
  HS65_LH_CNIVX3 U8467 ( .A(\u_DataPath/pc_4_to_ex_i [7]), .Z(n7419) );
  HS65_LH_NOR4ABX2 U8468 ( .A(n6416), .B(n6415), .C(n6414), .D(n6413), .Z(
        n8168) );
  HS65_LH_CNIVX3 U8469 ( .A(\u_DataPath/pc_4_to_ex_i [13]), .Z(n7434) );
  HS65_LH_AOI22X1 U8470 ( .A(n8313), .B(n9435), .C(n7695), .D(
        \u_DataPath/u_execute/link_value_i [29]), .Z(n7656) );
  HS65_LH_NOR4ABX2 U8471 ( .A(n6396), .B(n6395), .C(n6394), .D(n6393), .Z(
        n8203) );
  HS65_LH_NOR4ABX2 U8472 ( .A(n6013), .B(n6012), .C(n6011), .D(n6010), .Z(
        n8199) );
  HS65_LH_AOI22X1 U8473 ( .A(n8313), .B(n9143), .C(n7693), .D(
        \u_DataPath/u_execute/link_value_i [21]), .Z(n8201) );
  HS65_LH_NOR4ABX2 U8474 ( .A(n6643), .B(n6642), .C(n6641), .D(n6640), .Z(
        n8265) );
  HS65_LH_CNIVX3 U8475 ( .A(\u_DataPath/pc_4_to_ex_i [5]), .Z(n7620) );
  HS65_LL_AOI22X1 U8476 ( .A(n8687), .B(n9430), .C(n9252), .D(n8844), .Z(n8255) );
  HS65_LH_CNIVX3 U8477 ( .A(\u_DataPath/pc_4_to_ex_i [9]), .Z(n7623) );
  HS65_LH_NOR4ABX2 U8478 ( .A(n6286), .B(n6285), .C(n6284), .D(n6283), .Z(
        n8189) );
  HS65_LH_NOR4ABX2 U8479 ( .A(n5993), .B(n5992), .C(n5991), .D(n5990), .Z(
        n8068) );
  HS65_LH_NOR4ABX2 U8480 ( .A(n6542), .B(n6541), .C(n6540), .D(n6539), .Z(
        n8295) );
  HS65_LH_AOI22X1 U8481 ( .A(n8313), .B(n9452), .C(n7693), .D(
        \u_DataPath/u_execute/link_value_i [28]), .Z(n8293) );
  HS65_LH_NOR4ABX2 U8482 ( .A(n6562), .B(n6561), .C(n6560), .D(n6559), .Z(
        n8285) );
  HS65_LHS_XNOR2X3 U8483 ( .A(n9006), .B(n5908), .Z(
        \u_DataPath/u_execute/resAdd1_i [4]) );
  HS65_LH_NOR4ABX2 U8484 ( .A(n6436), .B(n6435), .C(n6434), .D(n6433), .Z(
        n8054) );
  HS65_LH_NOR4ABX2 U8485 ( .A(n6039), .B(n6038), .C(n6037), .D(n6036), .Z(
        n8018) );
  HS65_LH_NOR4ABX2 U8486 ( .A(n6663), .B(n6662), .C(n6661), .D(n6660), .Z(
        n8232) );
  HS65_LH_NOR4ABX2 U8487 ( .A(n6602), .B(n6601), .C(n6600), .D(n6599), .Z(
        n8292) );
  HS65_LH_AOI22X1 U8488 ( .A(n8313), .B(n8818), .C(n7693), .D(
        \u_DataPath/u_execute/link_value_i [20]), .Z(n8290) );
  HS65_LH_NOR4ABX2 U8489 ( .A(n6196), .B(n6195), .C(n6194), .D(n6193), .Z(
        n8188) );
  HS65_LH_NOR4ABX2 U8490 ( .A(n6079), .B(n6078), .C(n6077), .D(n6076), .Z(
        n8069) );
  HS65_LHS_XOR2X3 U8491 ( .A(n9408), .B(n7641), .Z(
        \u_DataPath/u_execute/link_value_i [16]) );
  HS65_LH_NOR4ABX2 U8492 ( .A(n6376), .B(n6375), .C(n6374), .D(n6373), .Z(
        n8194) );
  HS65_LH_NOR4ABX2 U8493 ( .A(n5971), .B(n5970), .C(n5969), .D(n5968), .Z(
        n8190) );
  HS65_LH_AOI22X1 U8494 ( .A(n8313), .B(n9135), .C(n7693), .D(
        \u_DataPath/u_execute/link_value_i [17]), .Z(n8192) );
  HS65_LH_AOI21X2 U8495 ( .A(n2797), .B(n9229), .C(n8377), .Z(
        \u_DataPath/mem_writedata_out_i [2]) );
  HS65_LH_AO112X4 U8496 ( .A(n8376), .B(n2798), .C(n8375), .D(rst), .Z(n8377)
         );
  HS65_LH_AO22X9 U8497 ( .A(n7682), .B(\u_DataPath/u_execute/resAdd1_i [2]), 
        .C(n7680), .D(\lte_x_57/B[2] ), .Z(\u_DataPath/jump_address_i [2]) );
  HS65_LHS_XOR2X3 U8498 ( .A(n9004), .B(n5914), .Z(
        \u_DataPath/u_execute/resAdd1_i [2]) );
  HS65_LH_NOR4ABX2 U8499 ( .A(n6236), .B(n6235), .C(n6234), .D(n6233), .Z(
        n8056) );
  HS65_LH_NOR4ABX2 U8500 ( .A(n6161), .B(n6160), .C(n6159), .D(n6158), .Z(
        n8281) );
  HS65_LH_NOR4ABX2 U8501 ( .A(n6683), .B(n6682), .C(n6681), .D(n6680), .Z(
        n8243) );
  HS65_LH_NOR4ABX2 U8502 ( .A(n6747), .B(n6746), .C(n6745), .D(n6744), .Z(
        n8247) );
  HS65_LH_AO22X9 U8504 ( .A(n7682), .B(n8869), .C(n7680), .D(n5497), .Z(
        \u_DataPath/jump_address_i [1]) );
  HS65_LH_CNIVX3 U8505 ( .A(n5861), .Z(n5862) );
  HS65_LH_NOR4ABX2 U8506 ( .A(n6257), .B(n6256), .C(n6255), .D(n6254), .Z(
        n8050) );
  HS65_LH_AO22X9 U8507 ( .A(n7683), .B(n8870), .C(n7680), .D(n2780), .Z(
        \u_DataPath/jump_address_i [0]) );
  HS65_LH_OR2X4 U8508 ( .A(n8500), .B(\u_DataPath/u_execute/link_value_i [0]), 
        .Z(n5731) );
  HS65_LH_NOR4ABX2 U8509 ( .A(n6216), .B(n6215), .C(n6214), .D(n6213), .Z(
        n8059) );
  HS65_LH_CNIVX3 U8510 ( .A(n7974), .Z(n7976) );
  HS65_LH_AOI22X1 U8511 ( .A(n8313), .B(n9360), .C(n7693), .D(
        \u_DataPath/u_execute/link_value_i [31]), .Z(n8309) );
  HS65_LH_NOR4ABX2 U8512 ( .A(n6622), .B(n6621), .C(n6620), .D(n6619), .Z(
        n8312) );
  HS65_LH_NAND2X2 U8513 ( .A(n9118), .B(n8468), .Z(n8073) );
  HS65_LH_NOR4ABX2 U8514 ( .A(n8737), .B(n9040), .C(n9303), .D(n8071), .Z(
        \u_DataPath/cw_exmem_i [3]) );
  HS65_LH_NAND2AX4 U8515 ( .A(n7712), .B(n9443), .Z(n8360) );
  HS65_LH_NAND2AX4 U8516 ( .A(n7712), .B(n8963), .Z(n8129) );
  HS65_LH_NAND3X2 U8517 ( .A(opcode_i[1]), .B(n7411), .C(n8070), .Z(n8072) );
  HS65_LH_NAND2AX4 U8518 ( .A(n7712), .B(n8879), .Z(n8185) );
  HS65_LH_AND2X4 U8519 ( .A(n1885), .B(n8969), .Z(
        \u_DataPath/pc4_to_idexreg_i [31]) );
  HS65_LH_NAND2AX4 U8520 ( .A(n7712), .B(n9441), .Z(n8115) );
  HS65_LH_NAND2AX4 U8521 ( .A(n7712), .B(n8830), .Z(n8116) );
  HS65_LH_NAND2AX4 U8522 ( .A(n7712), .B(n9439), .Z(n8119) );
  HS65_LH_NAND2AX4 U8523 ( .A(n7712), .B(n9399), .Z(n8121) );
  HS65_LH_NAND2AX4 U8524 ( .A(n7712), .B(n8833), .Z(n8122) );
  HS65_LH_NAND2AX4 U8525 ( .A(n7712), .B(n9345), .Z(n8124) );
  HS65_LH_NOR2X2 U8526 ( .A(n8045), .B(rst), .Z(n8461) );
  HS65_LH_AND2X4 U8527 ( .A(n1885), .B(\u_DataPath/toPC2_i [28]), .Z(
        \u_DataPath/branch_target_i [28]) );
  HS65_LH_CNIVX3 U8528 ( .A(n5557), .Z(n5558) );
  HS65_LH_AND2X4 U8529 ( .A(n1885), .B(\u_DataPath/toPC2_i [26]), .Z(
        \u_DataPath/branch_target_i [26]) );
  HS65_LHS_XOR2X3 U8530 ( .A(n8895), .B(n5614), .Z(\u_DataPath/toPC2_i [20])
         );
  HS65_LHS_XOR2X3 U8531 ( .A(n8927), .B(n5636), .Z(\u_DataPath/toPC2_i [19])
         );
  HS65_LHS_XOR2X3 U8532 ( .A(n8894), .B(n5627), .Z(\u_DataPath/toPC2_i [18])
         );
  HS65_LHS_XOR2X3 U8533 ( .A(n8919), .B(n5621), .Z(\u_DataPath/toPC2_i [17])
         );
  HS65_LHS_XOR2X3 U8534 ( .A(n9091), .B(n5579), .Z(\u_DataPath/toPC2_i [15])
         );
  HS65_LHS_XOR2X3 U8536 ( .A(n8929), .B(n5607), .Z(\u_DataPath/toPC2_i [13])
         );
  HS65_LHS_XOR2X3 U8537 ( .A(n8928), .B(n5598), .Z(\u_DataPath/toPC2_i [11])
         );
  HS65_LHS_XOR2X3 U8539 ( .A(n8923), .B(n2799), .Z(\u_DataPath/toPC2_i [8]) );
  HS65_LH_CNIVX3 U8540 ( .A(n5692), .Z(n5643) );
  HS65_LHS_XOR2X3 U8541 ( .A(n9057), .B(n5699), .Z(\u_DataPath/toPC2_i [6]) );
  HS65_LH_CNIVX3 U8542 ( .A(n5700), .Z(n5645) );
  HS65_LHS_XOR2X3 U8543 ( .A(n8921), .B(n5655), .Z(\u_DataPath/toPC2_i [5]) );
  HS65_LH_CNIVX3 U8544 ( .A(n5712), .Z(n5657) );
  HS65_LH_CNIVX3 U8545 ( .A(n5660), .Z(n5661) );
  HS65_LLS_XNOR2X3 U8546 ( .A(n3671), .B(n3670), .Z(n3672) );
  HS65_LH_IVX9 U8547 ( .A(n5014), .Z(n5446) );
  HS65_LH_AOI22X1 U8548 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][19] ), .B(n8851), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][19] ), .D(
        n8850), .Z(n6296) );
  HS65_LH_AOI22X1 U8549 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][16] ), .B(n8851), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][16] ), .D(
        n8850), .Z(n6178) );
  HS65_LH_AOI22X1 U8550 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][0] ), .B(n8851), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][0] ), .D(n8850), .Z(n6206) );
  HS65_LL_NAND3X5 U8551 ( .A(n2840), .B(n3041), .C(n3040), .Z(n3962) );
  HS65_LL_AND2X4 U8552 ( .A(n3174), .B(n8730), .Z(n2841) );
  HS65_LL_AND2X4 U8553 ( .A(n8702), .B(n2712), .Z(n2842) );
  HS65_LL_AND2X4 U8554 ( .A(n3174), .B(n8730), .Z(n2845) );
  HS65_LH_AND2X4 U8555 ( .A(n3184), .B(n8730), .Z(n2846) );
  HS65_LH_AND2X4 U8556 ( .A(n4446), .B(n4445), .Z(n2847) );
  HS65_LL_AO31X4 U8557 ( .A(n5418), .B(n5344), .C(n5046), .D(n5045), .Z(n2859)
         );
  HS65_LL_NOR2AX3 U8558 ( .A(n3188), .B(\sub_x_51/A[18] ), .Z(n3539) );
  HS65_LL_NAND2AX7 U8559 ( .A(n3098), .B(n3097), .Z(n5529) );
  HS65_LL_NOR2AX3 U8560 ( .A(\u_DataPath/from_alu_data_out_i [30]), .B(n3148), 
        .Z(n2863) );
  HS65_LLS_XNOR2X3 U8561 ( .A(n2867), .B(n8029), .Z(n2870) );
  HS65_LLS_XNOR2X3 U8562 ( .A(n2868), .B(n6488), .Z(n2869) );
  HS65_LH_NOR2X6 U8563 ( .A(\u_DataPath/dataOut_exe_i [6]), .B(n3178), .Z(
        n4879) );
  HS65_LL_MUXI21X2 U8565 ( .D0(n8795), .D1(\u_DataPath/from_mem_data_out_i [5]), .S0(n9415), .Z(n8263) );
  HS65_LH_NOR2X6 U8566 ( .A(n2938), .B(n2794), .Z(n5934) );
  HS65_LH_NOR2X6 U8569 ( .A(n2780), .B(n5487), .Z(n3779) );
  HS65_LL_MUXI21X2 U8570 ( .D0(n8878), .D1(\u_DataPath/from_mem_data_out_i [1]), .S0(n9415), .Z(n8157) );
  HS65_LH_NOR2X2 U8571 ( .A(\u_DataPath/dataOut_exe_i [1]), .B(n9012), .Z(
        n2965) );
  HS65_LH_OAI12X6 U8572 ( .A(n3779), .B(n3775), .C(n3777), .Z(n4184) );
  HS65_LH_IVX9 U8574 ( .A(n4346), .Z(n5207) );
  HS65_LH_NOR2X6 U8575 ( .A(n8668), .B(n3181), .Z(n3006) );
  HS65_LH_NOR2AX3 U8576 ( .A(n3008), .B(n3980), .Z(n3009) );
  HS65_LH_IVX9 U8577 ( .A(n5386), .Z(n3074) );
  HS65_LH_MUXI21X2 U8578 ( .D0(\u_DataPath/from_alu_data_out_i [9]), .D1(
        \u_DataPath/from_mem_data_out_i [9]), .S0(n3148), .Z(n8399) );
  HS65_LH_MUXI21X2 U8579 ( .D0(\u_DataPath/from_alu_data_out_i [15]), .D1(
        \u_DataPath/from_mem_data_out_i [15]), .S0(n3148), .Z(n8277) );
  HS65_LH_MUXI21X2 U8580 ( .D0(\u_DataPath/from_alu_data_out_i [14]), .D1(
        \u_DataPath/from_mem_data_out_i [14]), .S0(n3235), .Z(n8151) );
  HS65_LH_NOR2X6 U8581 ( .A(\lte_x_57/B[14] ), .B(n3079), .Z(n3888) );
  HS65_LH_MUXI21X2 U8582 ( .D0(\u_DataPath/from_alu_data_out_i [12]), .D1(
        \u_DataPath/from_mem_data_out_i [12]), .S0(n3235), .Z(n8237) );
  HS65_LH_NOR2AX3 U8583 ( .A(n8662), .B(n3980), .Z(n3056) );
  HS65_LH_MUXI21X2 U8584 ( .D0(\u_DataPath/from_alu_data_out_i [13]), .D1(
        \u_DataPath/from_mem_data_out_i [13]), .S0(n3235), .Z(n8410) );
  HS65_LH_MUXI21X2 U8585 ( .D0(\u_DataPath/from_alu_data_out_i [24]), .D1(
        \u_DataPath/from_mem_data_out_i [24]), .S0(n3148), .Z(n8138) );
  HS65_LH_MUXI21X2 U8586 ( .D0(\u_DataPath/from_alu_data_out_i [27]), .D1(
        \u_DataPath/from_mem_data_out_i [27]), .S0(n3235), .Z(n8205) );
  HS65_LH_MUXI21X2 U8587 ( .D0(\u_DataPath/from_alu_data_out_i [29]), .D1(
        \u_DataPath/from_mem_data_out_i [29]), .S0(n3235), .Z(n8270) );
  HS65_LH_MUXI21X2 U8588 ( .D0(\u_DataPath/from_alu_data_out_i [17]), .D1(
        \u_DataPath/from_mem_data_out_i [17]), .S0(n3235), .Z(n8191) );
  HS65_LH_MUXI21X2 U8589 ( .D0(\u_DataPath/from_alu_data_out_i [16]), .D1(
        \u_DataPath/from_mem_data_out_i [16]), .S0(n3235), .Z(n8148) );
  HS65_LH_NOR2X6 U8591 ( .A(\sub_x_51/A[16] ), .B(n2795), .Z(n4427) );
  HS65_LL_NOR2X3 U8592 ( .A(n5245), .B(n4427), .Z(n4368) );
  HS65_LL_NOR2X3 U8593 ( .A(\sub_x_51/A[18] ), .B(n3188), .Z(n3633) );
  HS65_LH_MUXI21X2 U8594 ( .D0(\u_DataPath/from_alu_data_out_i [23]), .D1(
        \u_DataPath/from_mem_data_out_i [23]), .S0(n3235), .Z(n8209) );
  HS65_LH_NOR2AX3 U8595 ( .A(n3161), .B(n3980), .Z(n3162) );
  HS65_LH_MUXI21X2 U8597 ( .D0(\u_DataPath/from_alu_data_out_i [20]), .D1(
        \u_DataPath/from_mem_data_out_i [20]), .S0(n3235), .Z(n8275) );
  HS65_LH_MUXI21X2 U8598 ( .D0(\u_DataPath/from_alu_data_out_i [21]), .D1(
        \u_DataPath/from_mem_data_out_i [21]), .S0(n3235), .Z(n8200) );
  HS65_LH_NAND2X7 U8599 ( .A(\sub_x_51/A[16] ), .B(n2795), .Z(n4426) );
  HS65_LL_NAND2X4 U8600 ( .A(\sub_x_51/A[20] ), .B(n3192), .Z(n5433) );
  HS65_LLS_XNOR2X3 U8601 ( .A(n3212), .B(n3211), .Z(n3309) );
  HS65_LL_NOR2X3 U8605 ( .A(\sub_x_51/A[22] ), .B(n5251), .Z(n4727) );
  HS65_LH_OAI22X1 U8608 ( .A(n3103), .B(n3322), .C(n3225), .D(n4901), .Z(n3287) );
  HS65_LH_OAI22X1 U8610 ( .A(n3993), .B(n3322), .C(n4918), .D(n2829), .Z(n3297) );
  HS65_LL_NAND3X2 U8611 ( .A(\u_DataPath/cw_to_ex_i [1]), .B(n5062), .C(n5329), 
        .Z(n3302) );
  HS65_LLS_XNOR2X3 U8612 ( .A(n3318), .B(n3317), .Z(n3371) );
  HS65_LH_CBI4I1X3 U8616 ( .A(n2802), .B(\sub_x_51/A[27] ), .C(n4781), .D(
        n3106), .Z(n3336) );
  HS65_LH_IVX9 U8617 ( .A(n4743), .Z(n4665) );
  HS65_LLS_XNOR2X3 U8620 ( .A(n3378), .B(n3377), .Z(n3428) );
  HS65_LH_CBI4I1X3 U8621 ( .A(n5507), .B(n5072), .C(n5506), .D(
        \lte_x_57/B[25] ), .Z(n3381) );
  HS65_LH_AOI22X1 U8623 ( .A(\sub_x_51/A[22] ), .B(n2792), .C(n5498), .D(n5192), .Z(n3406) );
  HS65_LH_IVX9 U8624 ( .A(\u_DataPath/cw_tomem_i [5]), .Z(n3434) );
  HS65_LH_IVX9 U8625 ( .A(\u_DataPath/cw_tomem_i [4]), .Z(n3438) );
  HS65_LL_AND2ABX18 U8626 ( .A(n7351), .B(n3430), .Z(write_byte_snps_wire) );
  HS65_LH_NAND2X7 U8627 ( .A(n8163), .B(n3432), .Z(n3563) );
  HS65_LL_NOR2AX25 U8628 ( .A(n9330), .B(n3567), .Z(Address_toRAM[9]) );
  HS65_LL_NOR2AX25 U8629 ( .A(\u_DataPath/dataOut_exe_i [12]), .B(n3567), .Z(
        Address_toRAM[10]) );
  HS65_LL_NOR2AX25 U8630 ( .A(n8734), .B(n3567), .Z(Address_toRAM[7]) );
  HS65_LL_NOR2AX25 U8632 ( .A(\u_DataPath/dataOut_exe_i [30]), .B(n3439), .Z(
        Address_toRAM[28]) );
  HS65_LL_NOR2AX25 U8633 ( .A(\u_DataPath/dataOut_exe_i [21]), .B(n3439), .Z(
        Address_toRAM[19]) );
  HS65_LL_NOR2AX25 U8634 ( .A(\u_DataPath/dataOut_exe_i [22]), .B(n3439), .Z(
        Address_toRAM[20]) );
  HS65_LL_NOR2AX25 U8635 ( .A(n9125), .B(n3439), .Z(Address_toRAM[22]) );
  HS65_LL_NOR2AX25 U8636 ( .A(\u_DataPath/dataOut_exe_i [28]), .B(n3439), .Z(
        Address_toRAM[26]) );
  HS65_LL_NOR2AX25 U8637 ( .A(\u_DataPath/dataOut_exe_i [15]), .B(n3567), .Z(
        Address_toRAM[13]) );
  HS65_LL_NOR2AX25 U8638 ( .A(\u_DataPath/dataOut_exe_i [27]), .B(n3439), .Z(
        Address_toRAM[25]) );
  HS65_LL_NOR2AX25 U8639 ( .A(\u_DataPath/dataOut_exe_i [23]), .B(n3439), .Z(
        Address_toRAM[21]) );
  HS65_LH_IVX9 U8641 ( .A(n4305), .Z(n5492) );
  HS65_LL_NOR2AX3 U8642 ( .A(n4214), .B(n3845), .Z(n3462) );
  HS65_LH_NAND2X2 U8643 ( .A(n4781), .B(n5064), .Z(n3469) );
  HS65_LH_NAND2X2 U8644 ( .A(n4620), .B(n5092), .Z(n3466) );
  HS65_LH_CNIVX3 U8646 ( .A(n4572), .Z(n3494) );
  HS65_LH_CNIVX3 U8658 ( .A(n7014), .Z(n3527) );
  HS65_LH_CNIVX3 U8659 ( .A(n6488), .Z(n7012) );
  HS65_LH_NAND3X2 U8660 ( .A(n7013), .B(n7012), .C(n7647), .Z(n7645) );
  HS65_LL_AND2X18 U8662 ( .A(n8564), .B(write_op), .Z(Data_in[6]) );
  HS65_LL_AND2X18 U8663 ( .A(n8584), .B(write_op), .Z(Data_in[5]) );
  HS65_LL_NOR2AX25 U8664 ( .A(n8553), .B(n3567), .Z(Address_toRAM[14]) );
  HS65_LL_NOR2AX25 U8665 ( .A(\u_DataPath/dataOut_exe_i [25]), .B(n3439), .Z(
        Address_toRAM[23]) );
  HS65_LL_NOR2AX25 U8666 ( .A(\u_DataPath/dataOut_exe_i [20]), .B(n3439), .Z(
        Address_toRAM[18]) );
  HS65_LL_NOR2AX25 U8669 ( .A(n8574), .B(n3450), .Z(Data_in[8]) );
  HS65_LL_NOR2AX25 U8671 ( .A(n8579), .B(n3450), .Z(Data_in[16]) );
  HS65_LL_AO112X18 U8672 ( .A(n8728), .B(n3564), .C(n8727), .D(n9438), .Z(
        read_op) );
  HS65_LL_OR2ABX18 U8673 ( .A(n2813), .B(n8456), .Z(nibble[1]) );
  HS65_LL_NOR2AX25 U8674 ( .A(n9541), .B(n3567), .Z(Address_toRAM[3]) );
  HS65_LL_NOR2AX25 U8675 ( .A(\u_DataPath/dataOut_exe_i [4]), .B(n3567), .Z(
        Address_toRAM[2]) );
  HS65_LL_NOR2AX25 U8676 ( .A(\u_DataPath/dataOut_exe_i [3]), .B(n3567), .Z(
        Address_toRAM[1]) );
  HS65_LL_NOR2AX25 U8677 ( .A(n9122), .B(n3568), .Z(Data_in[26]) );
  HS65_LL_NOR2AX25 U8678 ( .A(n8761), .B(n3568), .Z(Data_in[25]) );
  HS65_LL_NOR2AX25 U8679 ( .A(n9123), .B(n3568), .Z(Data_in[24]) );
  HS65_LL_AND2ABX18 U8680 ( .A(n9268), .B(n3439), .Z(Address_toRAM[5]) );
  HS65_LL_AND2X18 U8681 ( .A(n8567), .B(write_op), .Z(Data_in[4]) );
  HS65_LL_AND2X18 U8682 ( .A(n8565), .B(write_op), .Z(Data_in[0]) );
  HS65_LL_AND2X18 U8683 ( .A(n8572), .B(write_op), .Z(Data_in[3]) );
  HS65_LL_AND2X18 U8684 ( .A(n8704), .B(write_op), .Z(Data_in[2]) );
  HS65_LL_AND2X18 U8685 ( .A(n8568), .B(write_op), .Z(Data_in[1]) );
  HS65_LL_AND2X18 U8686 ( .A(n8578), .B(write_op), .Z(Data_in[7]) );
  HS65_LH_CBI4I1X3 U8688 ( .A(n5507), .B(n5392), .C(n5506), .D(
        \lte_x_57/B[14] ), .Z(n3577) );
  HS65_LH_NAND2X2 U8689 ( .A(\lte_x_57/B[30] ), .B(n4208), .Z(n3592) );
  HS65_LL_CBI4I1X3 U8691 ( .A(n5507), .B(n5186), .C(n5506), .D(
        \sub_x_51/A[16] ), .Z(n3641) );
  HS65_LHS_XNOR2X6 U8692 ( .A(n3138), .B(n5186), .Z(n4950) );
  HS65_LH_OAI21X3 U8699 ( .A(n3065), .B(n2829), .C(n3851), .Z(n3854) );
  HS65_LH_CBI4I1X3 U8701 ( .A(n5507), .B(n5208), .C(n5506), .D(\lte_x_57/B[4] ), .Z(n3857) );
  HS65_LH_NOR3X1 U8704 ( .A(n2776), .B(n4147), .C(n4332), .Z(n3931) );
  HS65_LH_NAND2X4 U8705 ( .A(n5354), .B(n5376), .Z(n3972) );
  HS65_LH_AOI21X2 U8706 ( .A(n5347), .B(n5415), .C(n5342), .Z(n3942) );
  HS65_LH_CNIVX3 U8709 ( .A(n8774), .Z(n3979) );
  HS65_LH_NOR2X6 U8710 ( .A(n3979), .B(n2794), .Z(n8451) );
  HS65_LH_NOR2X2 U8711 ( .A(n4383), .B(n5063), .Z(n3994) );
  HS65_LL_AOI12X3 U8712 ( .A(n4022), .B(n4021), .C(n4020), .Z(n8339) );
  HS65_LHS_XNOR2X3 U8713 ( .A(n5082), .B(n3065), .Z(n4957) );
  HS65_LLS_XNOR2X3 U8714 ( .A(n4086), .B(n4085), .Z(n4087) );
  HS65_LH_NAND2X2 U8717 ( .A(n4781), .B(n5203), .Z(n4151) );
  HS65_LHS_XNOR2X6 U8718 ( .A(n5203), .B(n3054), .Z(n4956) );
  HS65_LH_NAND2X2 U8719 ( .A(n4781), .B(n5092), .Z(n4191) );
  HS65_LLS_XNOR2X3 U8721 ( .A(n4243), .B(n4242), .Z(n4269) );
  HS65_LHS_XNOR2X6 U8722 ( .A(n5201), .B(n4283), .Z(n4975) );
  HS65_LL_CBI4I1X3 U8723 ( .A(n5507), .B(n5201), .C(n5506), .D(\sub_x_51/A[8] ), .Z(n4287) );
  HS65_LLS_XNOR2X3 U8726 ( .A(n4380), .B(n4379), .Z(n4395) );
  HS65_LLS_XNOR2X3 U8727 ( .A(n4383), .B(n5063), .Z(n4945) );
  HS65_LL_CBI4I1X3 U8728 ( .A(n5507), .B(n5063), .C(n5506), .D(
        \sub_x_51/A[18] ), .Z(n4384) );
  HS65_LLS_XNOR2X3 U8729 ( .A(n4404), .B(n4403), .Z(n4424) );
  HS65_LH_NAND2X2 U8731 ( .A(n3465), .B(n4946), .Z(n4434) );
  HS65_LH_CBI4I1X3 U8732 ( .A(n5507), .B(n5066), .C(n5506), .D(
        \sub_x_51/A[21] ), .Z(n4467) );
  HS65_LHS_XNOR2X3 U8733 ( .A(n4918), .B(n5066), .Z(n4952) );
  HS65_LH_NAND2X2 U8737 ( .A(n4604), .B(n4683), .Z(n4606) );
  HS65_LH_AOI22X1 U8740 ( .A(\lte_x_57/B[28] ), .B(n2792), .C(n2796), .D(
        \lte_x_57/B[29] ), .Z(n4660) );
  HS65_LLS_XNOR2X3 U8741 ( .A(n4717), .B(n4716), .Z(n4764) );
  HS65_LH_AND2X4 U8742 ( .A(n4730), .B(n4723), .Z(n4733) );
  HS65_LH_NAND2X2 U8745 ( .A(n4781), .B(n5211), .Z(n4782) );
  HS65_LH_OAI22X1 U8748 ( .A(n9538), .B(n4871), .C(n4870), .D(n2774), .Z(n4872) );
  HS65_LH_NAND2X2 U8749 ( .A(n4880), .B(n8388), .Z(n4881) );
  HS65_LH_NAND4ABX3 U8750 ( .A(n4892), .B(n4897), .C(n5039), .D(n4883), .Z(
        n4890) );
  HS65_LH_CBI4I6X2 U8751 ( .A(n5412), .B(n5334), .C(n5349), .D(n4892), .Z(
        n4893) );
  HS65_LH_OA112X9 U8752 ( .A(n5372), .B(n5376), .C(n5354), .D(n4896), .Z(n4898) );
  HS65_LH_NOR2X2 U8753 ( .A(n5529), .B(n5067), .Z(n4998) );
  HS65_LH_NAND4ABX3 U8754 ( .A(n5163), .B(n5162), .C(n5279), .D(n5164), .Z(
        n4995) );
  HS65_LH_NAND4ABX3 U8755 ( .A(n4956), .B(n4955), .C(n4954), .D(n4953), .Z(
        n4982) );
  HS65_LH_NAND4ABX3 U8756 ( .A(n4962), .B(n4961), .C(n4960), .D(n4959), .Z(
        n4969) );
  HS65_LHS_XNOR2X3 U8757 ( .A(\lte_x_57/B[14] ), .B(n5392), .Z(n4973) );
  HS65_LL_NOR3X1 U8759 ( .A(n4994), .B(n4993), .C(n4992), .Z(n5169) );
  HS65_LH_NAND3X2 U8760 ( .A(\u_DataPath/cw_to_ex_i [0]), .B(n5015), .C(n5449), 
        .Z(n5021) );
  HS65_LL_NAND2AX4 U8761 ( .A(n5029), .B(n5028), .Z(n5428) );
  HS65_LH_NOR4ABX2 U8762 ( .A(n5035), .B(n5427), .C(n5424), .D(n5428), .Z(
        n5050) );
  HS65_LH_CBI4I1X3 U8763 ( .A(n5406), .B(n5220), .C(n5404), .D(n5403), .Z(
        n5037) );
  HS65_LL_NOR2X2 U8766 ( .A(n3372), .B(n5139), .Z(n5074) );
  HS65_LL_NAND2X2 U8767 ( .A(n5103), .B(n5090), .Z(n5106) );
  HS65_LL_NOR2X2 U8768 ( .A(\lte_x_57/B[4] ), .B(n3241), .Z(n5097) );
  HS65_LH_AND2X4 U8769 ( .A(n2780), .B(n5487), .Z(n5095) );
  HS65_LH_AND2X4 U8770 ( .A(n3940), .B(n2968), .Z(n5093) );
  HS65_LH_AOI21X2 U8771 ( .A(n5100), .B(n5099), .C(n5098), .Z(n5105) );
  HS65_LH_AND2X4 U8774 ( .A(n7321), .B(n5148), .Z(n5149) );
  HS65_LL_NOR2X2 U8776 ( .A(\lte_x_57/B[4] ), .B(n3241), .Z(n5209) );
  HS65_LH_NOR2X2 U8777 ( .A(n2994), .B(\lte_x_57/B[2] ), .Z(n5212) );
  HS65_LH_NOR2X2 U8778 ( .A(n5212), .B(n5091), .Z(n5217) );
  HS65_LH_NAND2X2 U8780 ( .A(\lte_x_57/B[28] ), .B(n2791), .Z(n5265) );
  HS65_LH_NOR4ABX2 U8784 ( .A(n5356), .B(n5376), .C(n5373), .D(n5377), .Z(
        n5357) );
  HS65_LH_AOI22X1 U8786 ( .A(n5393), .B(n5392), .C(n3886), .D(n5391), .Z(n5399) );
  HS65_LH_AND2X4 U8788 ( .A(n5490), .B(n5489), .Z(n5491) );
  HS65_LH_AND2X4 U8789 ( .A(n5664), .B(n5531), .Z(\u_DataPath/toPC2_i [0]) );
  HS65_LH_CNIVX3 U8790 ( .A(n5581), .Z(n5582) );
  HS65_LH_CNIVX3 U8791 ( .A(n5616), .Z(n5617) );
  HS65_LHS_XOR2X3 U8793 ( .A(n5664), .B(n5663), .Z(\u_DataPath/toPC2_i [1]) );
  HS65_LH_OR2X4 U8794 ( .A(n8526), .B(\u_DataPath/pc_4_to_ex_i [31]), .Z(n5665) );
  HS65_LH_AND2X4 U8795 ( .A(n5865), .B(n5731), .Z(
        \u_DataPath/u_execute/resAdd1_i [0]) );
  HS65_LH_NAND2X7 U8797 ( .A(n8469), .B(\u_DataPath/pc_4_to_ex_i [10]), .Z(
        n5887) );
  HS65_LH_NAND2X7 U8798 ( .A(n8508), .B(\u_DataPath/pc_4_to_ex_i [12]), .Z(
        n5811) );
  HS65_LH_NAND2X7 U8799 ( .A(n8504), .B(\u_DataPath/pc_4_to_ex_i [14]), .Z(
        n5871) );
  HS65_LH_NAND2X7 U8800 ( .A(\u_DataPath/idex_rt_i [0]), .B(
        \u_DataPath/pc_4_to_ex_i [16]), .Z(n5883) );
  HS65_LH_NAND2X7 U8801 ( .A(\u_DataPath/idex_rt_i [1]), .B(
        \u_DataPath/pc_4_to_ex_i [17]), .Z(n5834) );
  HS65_LHS_XOR2X3 U8803 ( .A(n8915), .B(n5763), .Z(
        \u_DataPath/u_execute/resAdd1_i [29]) );
  HS65_LH_CNIVX3 U8804 ( .A(n5765), .Z(n5766) );
  HS65_LH_CNIVX3 U8805 ( .A(n5784), .Z(n5785) );
  HS65_LH_CNIVX3 U8806 ( .A(n5823), .Z(n5824) );
  HS65_LH_CNIVX3 U8807 ( .A(n5839), .Z(n5840) );
  HS65_LH_AOI21X2 U8808 ( .A(n9413), .B(n5908), .C(n9273), .Z(n5856) );
  HS65_LH_CNIVX3 U8809 ( .A(n5915), .Z(n5858) );
  HS65_LHS_XOR2X3 U8810 ( .A(n5865), .B(n5864), .Z(
        \u_DataPath/u_execute/resAdd1_i [1]) );
  HS65_LH_IVX9 U8811 ( .A(\u_DataPath/jaddr_i [17]), .Z(n5936) );
  HS65_LH_BFX9 U8812 ( .A(n6100), .Z(n7475) );
  HS65_LH_NOR4ABX2 U8813 ( .A(n5943), .B(n5942), .C(n5941), .D(n5940), .Z(
        n5971) );
  HS65_LH_NAND2X7 U8814 ( .A(n8016), .B(n5944), .Z(n5951) );
  HS65_LH_AOI22X1 U8815 ( .A(n9161), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][17] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][17] ), .D(n9095), 
        .Z(n5948) );
  HS65_LH_NOR2X6 U8816 ( .A(n5950), .B(n5961), .Z(n6109) );
  HS65_LH_NOR4ABX2 U8818 ( .A(n5948), .B(n5947), .C(n5946), .D(n5945), .Z(
        n5970) );
  HS65_LH_NAND2X7 U8819 ( .A(n8016), .B(n5949), .Z(n5957) );
  HS65_LH_NOR2X6 U8820 ( .A(n5961), .B(n5952), .Z(n6026) );
  HS65_LH_NOR2X6 U8821 ( .A(n5950), .B(n5963), .Z(n6027) );
  HS65_LH_AO22X4 U8822 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][17] ), .B(n8867), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][17] ), .D(
        n8866), .Z(n5955) );
  HS65_LH_NOR2X6 U8823 ( .A(n5961), .B(n5951), .Z(n5980) );
  HS65_LH_NOR2X6 U8824 ( .A(n5963), .B(n5952), .Z(n5981) );
  HS65_LH_NOR2X6 U8825 ( .A(n5963), .B(n5957), .Z(n6122) );
  HS65_LH_NAND4ABX3 U8826 ( .A(n5956), .B(n5955), .C(n5954), .D(n5953), .Z(
        n5969) );
  HS65_LH_NOR2X6 U8827 ( .A(n5959), .B(n5962), .Z(n6132) );
  HS65_LH_NOR2X6 U8828 ( .A(n5963), .B(n5962), .Z(n6133) );
  HS65_LH_AOI22X1 U8829 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][17] ), .B(n9113), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][17] ), .D(
        n9166), .Z(n5964) );
  HS65_LH_NAND4ABX3 U8830 ( .A(n5967), .B(n5966), .C(n5965), .D(n5964), .Z(
        n5968) );
  HS65_LH_NOR4ABX2 U8831 ( .A(n5975), .B(n5974), .C(n5973), .D(n5972), .Z(
        n5993) );
  HS65_LH_BFX9 U8832 ( .A(n6108), .Z(n7509) );
  HS65_LH_AO22X9 U8833 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][24] ), .B(n9364), 
        .C(n9253), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][24] ), .Z(n5977)
         );
  HS65_LH_NOR4ABX2 U8834 ( .A(n5979), .B(n5978), .C(n5977), .D(n5976), .Z(
        n5992) );
  HS65_LH_AO22X4 U8835 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][24] ), .B(n9102), 
        .C(n9101), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][24] ), .Z(n5985)
         );
  HS65_LH_AO22X4 U8836 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][24] ), .B(n8867), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][24] ), .D(
        n8866), .Z(n5984) );
  HS65_LH_NAND4ABX3 U8837 ( .A(n5985), .B(n5984), .C(n5983), .D(n5982), .Z(
        n5991) );
  HS65_LH_AO22X4 U8838 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][24] ), .B(n9152), 
        .C(n9097), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][24] ), .Z(n5989)
         );
  HS65_LH_AO22X4 U8839 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][24] ), .B(n9070), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][24] ), .D(
        n9064), .Z(n5988) );
  HS65_LH_AOI22X1 U8840 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][24] ), .B(n9113), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][24] ), .D(
        n8861), .Z(n5986) );
  HS65_LH_NAND4ABX3 U8841 ( .A(n5989), .B(n5988), .C(n5987), .D(n5986), .Z(
        n5990) );
  HS65_LH_NOR4ABX2 U8842 ( .A(n5997), .B(n5996), .C(n5995), .D(n5994), .Z(
        n6013) );
  HS65_LH_AOI22X1 U8843 ( .A(n9161), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][21] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][21] ), .D(n9095), 
        .Z(n6001) );
  HS65_LH_AO22X9 U8844 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][21] ), .B(n9364), 
        .C(n9068), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][21] ), .Z(n5999)
         );
  HS65_LH_NOR4ABX2 U8845 ( .A(n6001), .B(n6000), .C(n5999), .D(n5998), .Z(
        n6012) );
  HS65_LH_AO22X4 U8846 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][21] ), .B(n8867), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][21] ), .D(
        n8866), .Z(n6004) );
  HS65_LH_NAND4ABX3 U8847 ( .A(n6005), .B(n6004), .C(n6003), .D(n6002), .Z(
        n6011) );
  HS65_LH_AOI22X1 U8848 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][21] ), .B(n9113), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][21] ), .D(
        n9166), .Z(n6006) );
  HS65_LH_NAND4ABX3 U8849 ( .A(n6009), .B(n6008), .C(n6007), .D(n6006), .Z(
        n6010) );
  HS65_LH_BFX9 U8850 ( .A(n6014), .Z(n7570) );
  HS65_LH_BFX9 U8851 ( .A(n6015), .Z(n7569) );
  HS65_LH_BFX9 U8852 ( .A(n6016), .Z(n7572) );
  HS65_LH_BFX9 U8853 ( .A(n6017), .Z(n7571) );
  HS65_LH_NOR4ABX2 U8854 ( .A(n6021), .B(n6020), .C(n6019), .D(n6018), .Z(
        n6039) );
  HS65_LH_NOR4ABX2 U8856 ( .A(n6025), .B(n6024), .C(n6023), .D(n6022), .Z(
        n6038) );
  HS65_LH_BFX9 U8857 ( .A(n6026), .Z(n7593) );
  HS65_LH_BFX9 U8858 ( .A(n6027), .Z(n7594) );
  HS65_LH_NAND4ABX3 U8860 ( .A(n6031), .B(n6030), .C(n6029), .D(n6028), .Z(
        n6037) );
  HS65_LH_AO22X4 U8861 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][4] ), .B(n9152), 
        .C(n9097), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][4] ), .Z(n6035) );
  HS65_LH_NAND4ABX3 U8862 ( .A(n6035), .B(n6034), .C(n6033), .D(n6032), .Z(
        n6036) );
  HS65_LH_NOR4ABX2 U8863 ( .A(n6043), .B(n6042), .C(n6041), .D(n6040), .Z(
        n6059) );
  HS65_LH_AO22X4 U8864 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][7] ), .B(n9364), 
        .C(n9253), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][7] ), .Z(n6045)
         );
  HS65_LH_NOR4ABX2 U8865 ( .A(n6047), .B(n6046), .C(n6045), .D(n6044), .Z(
        n6058) );
  HS65_LH_AO22X4 U8866 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][7] ), .B(n9102), 
        .C(n9101), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][7] ), .Z(n6051) );
  HS65_LH_AO22X4 U8867 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][7] ), .B(n8867), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][7] ), .D(
        n8866), .Z(n6050) );
  HS65_LH_NAND4ABX3 U8868 ( .A(n6051), .B(n6050), .C(n6049), .D(n6048), .Z(
        n6057) );
  HS65_LH_AO22X4 U8869 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][7] ), .B(n9152), 
        .C(n9097), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][7] ), .Z(n6055) );
  HS65_LH_AOI22X1 U8870 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][7] ), .B(n9113), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][7] ), .D(n8861), .Z(n6052) );
  HS65_LH_NAND4ABX3 U8871 ( .A(n6055), .B(n6054), .C(n6053), .D(n6052), .Z(
        n6056) );
  HS65_LH_NOR4ABX2 U8872 ( .A(n6063), .B(n6062), .C(n6061), .D(n6060), .Z(
        n6079) );
  HS65_LH_NOR4ABX2 U8874 ( .A(n6067), .B(n6066), .C(n6065), .D(n6064), .Z(
        n6078) );
  HS65_LH_AO22X4 U8875 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][16] ), .B(n9102), 
        .C(n9101), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][16] ), .Z(n6071)
         );
  HS65_LH_AO22X4 U8876 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][16] ), .B(n8867), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][16] ), .D(
        n8866), .Z(n6070) );
  HS65_LH_NAND4ABX3 U8877 ( .A(n6071), .B(n6070), .C(n6069), .D(n6068), .Z(
        n6077) );
  HS65_LH_AO22X4 U8878 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][16] ), .B(n9070), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][16] ), .D(
        n9064), .Z(n6074) );
  HS65_LH_AOI22X1 U8879 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][16] ), .B(n9113), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][16] ), .D(
        n8861), .Z(n6072) );
  HS65_LH_NAND4ABX3 U8880 ( .A(n6075), .B(n6074), .C(n6073), .D(n6072), .Z(
        n6076) );
  HS65_LH_AO22X4 U8881 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][14] ), .B(n8948), 
        .C(n8951), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][14] ), .Z(n6080)
         );
  HS65_LH_NOR4ABX2 U8882 ( .A(n6083), .B(n6082), .C(n6081), .D(n6080), .Z(
        n6099) );
  HS65_LH_AO22X9 U8883 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][14] ), .B(n9364), 
        .C(n9253), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][14] ), .Z(n6085)
         );
  HS65_LH_NOR4ABX2 U8884 ( .A(n6087), .B(n6086), .C(n6085), .D(n6084), .Z(
        n6098) );
  HS65_LH_AO22X4 U8885 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][14] ), .B(n9102), 
        .C(n9101), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][14] ), .Z(n6091)
         );
  HS65_LH_AO22X4 U8886 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][14] ), .B(n8867), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][14] ), .D(
        n8866), .Z(n6090) );
  HS65_LH_NAND4ABX3 U8887 ( .A(n6091), .B(n6090), .C(n6089), .D(n6088), .Z(
        n6097) );
  HS65_LH_NAND4ABX3 U8888 ( .A(n6095), .B(n6094), .C(n6093), .D(n6092), .Z(
        n6096) );
  HS65_LH_BFX9 U8889 ( .A(n6101), .Z(n7278) );
  HS65_LH_BFX9 U8890 ( .A(n6102), .Z(n7280) );
  HS65_LH_BFX9 U8891 ( .A(n6103), .Z(n7279) );
  HS65_LH_NOR4ABX2 U8892 ( .A(n6107), .B(n6106), .C(n6105), .D(n6104), .Z(
        n6141) );
  HS65_LH_AOI22X1 U8893 ( .A(n9161), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][3] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][3] ), .D(n9095), 
        .Z(n6118) );
  HS65_LH_BFX9 U8894 ( .A(n6110), .Z(n7555) );
  HS65_LH_AO22X4 U8895 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][3] ), .B(n9153), 
        .C(n9068), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][3] ), .Z(n6116)
         );
  HS65_LH_AO22X4 U8896 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][3] ), .B(n9165), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][3] ), .D(
        n9065), .Z(n6115) );
  HS65_LH_NOR4ABX2 U8897 ( .A(n6118), .B(n6117), .C(n6116), .D(n6115), .Z(
        n6140) );
  HS65_LH_AO22X4 U8898 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][3] ), .B(n9102), 
        .C(n9101), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][3] ), .Z(n6126) );
  HS65_LH_NAND4ABX3 U8899 ( .A(n6126), .B(n6125), .C(n6124), .D(n6123), .Z(
        n6139) );
  HS65_LH_AO22X4 U8900 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][3] ), .B(n9152), 
        .C(n9097), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][3] ), .Z(n6137) );
  HS65_LH_AO22X4 U8901 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][3] ), .B(n9070), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][3] ), .D(
        n9064), .Z(n6136) );
  HS65_LH_NAND4ABX3 U8902 ( .A(n6137), .B(n6136), .C(n6135), .D(n6134), .Z(
        n6138) );
  HS65_LH_NOR4ABX2 U8903 ( .A(n6145), .B(n6144), .C(n6143), .D(n6142), .Z(
        n6161) );
  HS65_LH_AOI22X1 U8904 ( .A(n9161), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][2] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][2] ), .D(n9095), 
        .Z(n6149) );
  HS65_LH_AO22X4 U8905 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][2] ), .B(n9153), 
        .C(n9068), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][2] ), .Z(n6147)
         );
  HS65_LH_AO22X4 U8906 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][2] ), .B(n9165), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][2] ), .D(
        n9065), .Z(n6146) );
  HS65_LH_NOR4ABX2 U8907 ( .A(n6149), .B(n6148), .C(n6147), .D(n6146), .Z(
        n6160) );
  HS65_LH_AO22X4 U8908 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][2] ), .B(n9102), 
        .C(n9101), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][2] ), .Z(n6153) );
  HS65_LH_NAND4ABX3 U8910 ( .A(n6153), .B(n6152), .C(n6151), .D(n6150), .Z(
        n6159) );
  HS65_LH_AO22X4 U8911 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][2] ), .B(n9152), 
        .C(n9097), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][2] ), .Z(n6157) );
  HS65_LH_AO22X4 U8912 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][2] ), .B(n9070), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][2] ), .D(
        n9064), .Z(n6156) );
  HS65_LH_NAND4ABX3 U8913 ( .A(n6157), .B(n6156), .C(n6155), .D(n6154), .Z(
        n6158) );
  HS65_LH_NOR2X6 U8914 ( .A(n6188), .B(n6162), .Z(n6497) );
  HS65_LH_BFX9 U8915 ( .A(n6497), .Z(n6457) );
  HS65_LH_NOR2X6 U8916 ( .A(n6182), .B(n6162), .Z(n6498) );
  HS65_LH_BFX9 U8917 ( .A(n6259), .Z(n6972) );
  HS65_LH_NOR2X6 U8918 ( .A(n6186), .B(n6164), .Z(n6975) );
  HS65_LH_NOR2X6 U8919 ( .A(n6184), .B(n6164), .Z(n6499) );
  HS65_LH_AO22X9 U8920 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][16] ), .B(n9472), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][16] ), .D(
        n8857), .Z(n6166) );
  HS65_LH_NOR2X6 U8921 ( .A(n6182), .B(n6164), .Z(n6976) );
  HS65_LH_NOR4ABX2 U8923 ( .A(n6168), .B(n6167), .C(n6166), .D(n6165), .Z(
        n6196) );
  HS65_LH_NAND2X7 U8924 ( .A(n2818), .B(n6169), .Z(n6174) );
  HS65_LH_NOR2X6 U8925 ( .A(n6186), .B(n6174), .Z(n6265) );
  HS65_LH_AOI22X1 U8926 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][16] ), .B(n8950), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][16] ), .D(
        n8855), .Z(n6173) );
  HS65_LH_NOR2X6 U8927 ( .A(n6188), .B(n6176), .Z(n6266) );
  HS65_LH_AOI22X1 U8928 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][16] ), .B(n9162), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][16] ), .D(
        n8854), .Z(n6172) );
  HS65_LH_NOR2X6 U8929 ( .A(n6174), .B(n6184), .Z(n6267) );
  HS65_LH_NOR2X6 U8930 ( .A(n6184), .B(n6175), .Z(n6312) );
  HS65_LH_BFX9 U8931 ( .A(n6312), .Z(n6910) );
  HS65_LH_AO22X9 U8932 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][16] ), .B(n9187), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][16] ), .D(
        n9194), .Z(n6170) );
  HS65_LH_NOR4ABX2 U8933 ( .A(n6173), .B(n6172), .C(n6171), .D(n6170), .Z(
        n6195) );
  HS65_LH_AO22X9 U8934 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][16] ), .B(n9249), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][16] ), .D(
        n9185), .Z(n6180) );
  HS65_LH_NAND3X5 U8936 ( .A(\u_DataPath/jaddr_i [24]), .B(n2811), .C(n2817), 
        .Z(n6187) );
  HS65_LH_NOR2X6 U8937 ( .A(n6182), .B(n6187), .Z(n6339) );
  HS65_LH_NOR2X6 U8938 ( .A(n2812), .B(\u_DataPath/jaddr_i [24]), .Z(n6181) );
  HS65_LH_NAND2X7 U8939 ( .A(n2818), .B(n6181), .Z(n6185) );
  HS65_LH_NOR2X6 U8940 ( .A(n6186), .B(n6185), .Z(n6245) );
  HS65_LH_NAND4ABX3 U8941 ( .A(n6180), .B(n6179), .C(n6178), .D(n6177), .Z(
        n6194) );
  HS65_LH_NAND2X7 U8942 ( .A(n2817), .B(n6181), .Z(n6183) );
  HS65_LH_NOR2X6 U8943 ( .A(n6186), .B(n6183), .Z(n6277) );
  HS65_LH_AO22X9 U8944 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][16] ), .B(n9470), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][16] ), .D(
        n9164), .Z(n6191) );
  HS65_LH_NOR2X6 U8945 ( .A(n6188), .B(n6185), .Z(n6299) );
  HS65_LH_BFX9 U8946 ( .A(n6299), .Z(n7002) );
  HS65_LH_NAND4ABX3 U8947 ( .A(n6192), .B(n6191), .C(n6190), .D(n6189), .Z(
        n6193) );
  HS65_LH_AO22X9 U8948 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][0] ), .B(n9472), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][0] ), .D(
        n8857), .Z(n6198) );
  HS65_LH_NOR4ABX2 U8950 ( .A(n6200), .B(n6199), .C(n6198), .D(n6197), .Z(
        n6216) );
  HS65_LH_AOI22X1 U8951 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][0] ), .B(n8950), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][0] ), .D(
        n8855), .Z(n6204) );
  HS65_LH_AOI22X1 U8952 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][0] ), .B(n9162), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][0] ), .D(
        n8854), .Z(n6203) );
  HS65_LH_AO22X9 U8953 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][0] ), .B(n9156), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][0] ), .D(
        n9475), .Z(n6202) );
  HS65_LH_AO22X9 U8954 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][0] ), .B(n9187), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][0] ), .D(
        n9194), .Z(n6201) );
  HS65_LH_NOR4ABX2 U8955 ( .A(n6204), .B(n6203), .C(n6202), .D(n6201), .Z(
        n6215) );
  HS65_LH_AO22X9 U8956 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][0] ), .B(n9249), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][0] ), .D(
        n9185), .Z(n6208) );
  HS65_LH_NAND4ABX3 U8957 ( .A(n6208), .B(n6207), .C(n6206), .D(n6205), .Z(
        n6214) );
  HS65_LH_AO22X9 U8958 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][0] ), .B(n9470), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][0] ), .D(n9164), .Z(n6211) );
  HS65_LH_NAND4ABX3 U8959 ( .A(n6212), .B(n6211), .C(n6210), .D(n6209), .Z(
        n6213) );
  HS65_LH_AO22X9 U8960 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][2] ), .B(n9472), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][2] ), .D(
        n8857), .Z(n6218) );
  HS65_LH_AO22X9 U8961 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][2] ), .B(n9473), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][2] ), .D(
        n9474), .Z(n6217) );
  HS65_LH_NOR4ABX2 U8962 ( .A(n6220), .B(n6219), .C(n6218), .D(n6217), .Z(
        n6236) );
  HS65_LH_AOI22X1 U8963 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][2] ), .B(n8950), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][2] ), .D(
        n8855), .Z(n6224) );
  HS65_LH_AOI22X1 U8964 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][2] ), .B(n9162), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][2] ), .D(
        n8854), .Z(n6223) );
  HS65_LH_AO22X9 U8965 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][2] ), .B(n9156), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][2] ), .D(
        n9475), .Z(n6222) );
  HS65_LH_NOR4ABX2 U8967 ( .A(n6224), .B(n6223), .C(n6222), .D(n6221), .Z(
        n6235) );
  HS65_LH_AO22X9 U8968 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][2] ), .B(n9249), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][2] ), .D(
        n9185), .Z(n6228) );
  HS65_LH_NAND4ABX3 U8969 ( .A(n6228), .B(n6227), .C(n6226), .D(n6225), .Z(
        n6234) );
  HS65_LH_NAND4ABX3 U8970 ( .A(n6232), .B(n6231), .C(n6230), .D(n6229), .Z(
        n6233) );
  HS65_LH_AO22X9 U8971 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][1] ), .B(n9196), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][1] ), .D(
        n9157), .Z(n6238) );
  HS65_LH_NOR4ABX2 U8972 ( .A(n6240), .B(n6239), .C(n6238), .D(n6237), .Z(
        n6257) );
  HS65_LH_AOI22X1 U8973 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][1] ), .B(n8950), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][1] ), .D(
        n8855), .Z(n6244) );
  HS65_LH_AOI22X1 U8974 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][1] ), .B(n9162), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][1] ), .D(
        n8854), .Z(n6243) );
  HS65_LH_AO22X9 U8975 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][1] ), .B(n9156), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][1] ), .D(
        n9475), .Z(n6242) );
  HS65_LH_NOR4ABX2 U8977 ( .A(n6244), .B(n6243), .C(n6242), .D(n6241), .Z(
        n6256) );
  HS65_LH_AO22X9 U8978 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][1] ), .B(n9249), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][1] ), .D(
        n9185), .Z(n6249) );
  HS65_LH_NAND4ABX3 U8979 ( .A(n6249), .B(n6248), .C(n6247), .D(n6246), .Z(
        n6255) );
  HS65_LH_NAND4ABX3 U8980 ( .A(n6253), .B(n6252), .C(n6251), .D(n6250), .Z(
        n6254) );
  HS65_LH_BFX9 U8981 ( .A(n6258), .Z(n6724) );
  HS65_LH_NOR4ABX2 U8984 ( .A(n6263), .B(n6262), .C(n6261), .D(n6260), .Z(
        n6286) );
  HS65_LH_BFX9 U8985 ( .A(n6264), .Z(n6982) );
  HS65_LH_BFX9 U8986 ( .A(n6266), .Z(n6983) );
  HS65_LH_NOR4ABX2 U8987 ( .A(n6271), .B(n6270), .C(n6269), .D(n6268), .Z(
        n6285) );
  HS65_LH_NAND4ABX3 U8989 ( .A(n6276), .B(n6275), .C(n6274), .D(n6273), .Z(
        n6284) );
  HS65_LH_BFX9 U8990 ( .A(n6277), .Z(n6998) );
  HS65_LH_NAND4ABX3 U8991 ( .A(n6282), .B(n6281), .C(n6280), .D(n6279), .Z(
        n6283) );
  HS65_LH_NOR4ABX2 U8994 ( .A(n6290), .B(n6289), .C(n6288), .D(n6287), .Z(
        n6307) );
  HS65_LH_NOR4ABX2 U8995 ( .A(n6294), .B(n6293), .C(n6292), .D(n6291), .Z(
        n6306) );
  HS65_LH_AO22X9 U8996 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][19] ), .B(n9249), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][19] ), .D(
        n9185), .Z(n6298) );
  HS65_LH_NAND4ABX3 U8997 ( .A(n6298), .B(n6297), .C(n6296), .D(n6295), .Z(
        n6305) );
  HS65_LH_NAND4ABX3 U8998 ( .A(n6303), .B(n6302), .C(n6301), .D(n6300), .Z(
        n6304) );
  HS65_LH_AO22X9 U9000 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][27] ), .B(n9473), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][27] ), .D(
        n9474), .Z(n6308) );
  HS65_LH_NOR4ABX2 U9001 ( .A(n6311), .B(n6310), .C(n6309), .D(n6308), .Z(
        n6328) );
  HS65_LH_NOR4ABX2 U9002 ( .A(n6316), .B(n6315), .C(n6314), .D(n6313), .Z(
        n6327) );
  HS65_LH_AO22X9 U9003 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][27] ), .B(n9249), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][27] ), .D(
        n9185), .Z(n6320) );
  HS65_LH_NAND4ABX3 U9004 ( .A(n6320), .B(n6319), .C(n6318), .D(n6317), .Z(
        n6326) );
  HS65_LH_NAND4ABX3 U9005 ( .A(n6324), .B(n6323), .C(n6322), .D(n6321), .Z(
        n6325) );
  HS65_LH_AO22X9 U9006 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][23] ), .B(n9472), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][23] ), .D(
        n8857), .Z(n6330) );
  HS65_LH_AO22X9 U9007 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][23] ), .B(n9473), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][23] ), .D(
        n9474), .Z(n6329) );
  HS65_LH_NOR4ABX2 U9008 ( .A(n6332), .B(n6331), .C(n6330), .D(n6329), .Z(
        n6356) );
  HS65_LH_BFX9 U9009 ( .A(n6333), .Z(n6984) );
  HS65_LH_BFX9 U9010 ( .A(n6986), .Z(n6911) );
  HS65_LH_NOR4ABX2 U9011 ( .A(n6337), .B(n6336), .C(n6335), .D(n6334), .Z(
        n6355) );
  HS65_LH_AO22X9 U9012 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][23] ), .B(n8940), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][23] ), .D(
        n8949), .Z(n6344) );
  HS65_LH_BFX9 U9013 ( .A(n6338), .Z(n6991) );
  HS65_LH_AO22X9 U9014 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][23] ), .B(n8939), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][23] ), .D(
        n9186), .Z(n6343) );
  HS65_LH_NAND4ABX3 U9015 ( .A(n6344), .B(n6343), .C(n6342), .D(n6341), .Z(
        n6354) );
  HS65_LH_AO22X9 U9016 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][23] ), .B(n9470), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][23] ), .D(
        n9267), .Z(n6351) );
  HS65_LH_NAND4ABX3 U9017 ( .A(n6352), .B(n6351), .C(n6350), .D(n6349), .Z(
        n6353) );
  HS65_LH_AO22X9 U9018 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][17] ), .B(n9472), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][17] ), .D(
        n8857), .Z(n6358) );
  HS65_LH_AO22X9 U9019 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][17] ), .B(n9473), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][17] ), .D(
        n9474), .Z(n6357) );
  HS65_LH_NOR4ABX2 U9020 ( .A(n6360), .B(n6359), .C(n6358), .D(n6357), .Z(
        n6376) );
  HS65_LH_AO22X9 U9021 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][17] ), .B(n9156), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][17] ), .D(
        n9475), .Z(n6362) );
  HS65_LH_AO22X9 U9022 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][17] ), .B(n9154), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][17] ), .D(
        n9194), .Z(n6361) );
  HS65_LH_NOR4ABX2 U9023 ( .A(n6364), .B(n6363), .C(n6362), .D(n6361), .Z(
        n6375) );
  HS65_LH_AO22X9 U9024 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][17] ), .B(n9249), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][17] ), .D(
        n9185), .Z(n6368) );
  HS65_LH_NAND4ABX3 U9025 ( .A(n6368), .B(n6367), .C(n6366), .D(n6365), .Z(
        n6374) );
  HS65_LH_NAND4ABX3 U9026 ( .A(n6372), .B(n6371), .C(n6370), .D(n6369), .Z(
        n6373) );
  HS65_LH_AO22X9 U9027 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][21] ), .B(n9472), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][21] ), .D(
        n8857), .Z(n6378) );
  HS65_LH_NOR4ABX2 U9029 ( .A(n6380), .B(n6379), .C(n6378), .D(n6377), .Z(
        n6396) );
  HS65_LH_AOI22X1 U9030 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][21] ), .B(n8950), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][21] ), .D(
        n8855), .Z(n6384) );
  HS65_LH_AO22X9 U9031 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][21] ), .B(n9154), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][21] ), .D(
        n9194), .Z(n6381) );
  HS65_LH_NOR4ABX2 U9032 ( .A(n6384), .B(n6383), .C(n6382), .D(n6381), .Z(
        n6395) );
  HS65_LH_AO22X9 U9033 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][21] ), .B(n9249), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][21] ), .D(
        n9185), .Z(n6388) );
  HS65_LH_NAND4ABX3 U9034 ( .A(n6388), .B(n6387), .C(n6386), .D(n6385), .Z(
        n6394) );
  HS65_LH_NAND4ABX3 U9035 ( .A(n6392), .B(n6391), .C(n6390), .D(n6389), .Z(
        n6393) );
  HS65_LH_AO22X9 U9037 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][13] ), .B(n9473), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][13] ), .D(
        n9474), .Z(n6397) );
  HS65_LH_NOR4ABX2 U9038 ( .A(n6400), .B(n6399), .C(n6398), .D(n6397), .Z(
        n6416) );
  HS65_LH_AO22X9 U9039 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][13] ), .B(n9187), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][13] ), .D(
        n9194), .Z(n6401) );
  HS65_LH_NOR4ABX2 U9040 ( .A(n6404), .B(n6403), .C(n6402), .D(n6401), .Z(
        n6415) );
  HS65_LH_AO22X9 U9041 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][13] ), .B(n9249), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][13] ), .D(
        n9185), .Z(n6408) );
  HS65_LH_NAND4ABX3 U9042 ( .A(n6408), .B(n6407), .C(n6406), .D(n6405), .Z(
        n6414) );
  HS65_LH_NAND4ABX3 U9043 ( .A(n6412), .B(n6411), .C(n6410), .D(n6409), .Z(
        n6413) );
  HS65_LH_AO22X9 U9045 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][4] ), .B(n9473), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][4] ), .D(
        n9474), .Z(n6417) );
  HS65_LH_NOR4ABX2 U9046 ( .A(n6420), .B(n6419), .C(n6418), .D(n6417), .Z(
        n6436) );
  HS65_LH_AOI22X1 U9047 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][4] ), .B(n8950), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][4] ), .D(
        n8855), .Z(n6424) );
  HS65_LH_AO22X9 U9048 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][4] ), .B(n9187), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][4] ), .D(
        n9194), .Z(n6421) );
  HS65_LH_NOR4ABX2 U9049 ( .A(n6424), .B(n6423), .C(n6422), .D(n6421), .Z(
        n6435) );
  HS65_LH_NAND4ABX3 U9051 ( .A(n6428), .B(n6427), .C(n6426), .D(n6425), .Z(
        n6434) );
  HS65_LH_NAND4ABX3 U9052 ( .A(n6432), .B(n6431), .C(n6430), .D(n6429), .Z(
        n6433) );
  HS65_LH_AO22X9 U9054 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][3] ), .B(n9473), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][3] ), .D(
        n9474), .Z(n6437) );
  HS65_LH_NOR4ABX2 U9055 ( .A(n6440), .B(n6439), .C(n6438), .D(n6437), .Z(
        n6456) );
  HS65_LH_AO22X9 U9056 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][3] ), .B(n9469), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][3] ), .D(
        n9475), .Z(n6442) );
  HS65_LH_NOR4ABX2 U9057 ( .A(n6444), .B(n6443), .C(n6442), .D(n6441), .Z(
        n6455) );
  HS65_LH_AO22X9 U9058 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][3] ), .B(n8940), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][3] ), .D(
        n9185), .Z(n6448) );
  HS65_LH_NAND4ABX3 U9059 ( .A(n6448), .B(n6447), .C(n6446), .D(n6445), .Z(
        n6454) );
  HS65_LH_AO22X9 U9061 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][3] ), .B(n9160), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][3] ), .D(n9164), .Z(n6451) );
  HS65_LH_NAND4ABX3 U9062 ( .A(n6452), .B(n6451), .C(n6450), .D(n6449), .Z(
        n6453) );
  HS65_LH_NOR4ABX2 U9065 ( .A(n6461), .B(n6460), .C(n6459), .D(n6458), .Z(
        n6477) );
  HS65_LH_AO22X9 U9066 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][7] ), .B(n9469), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][7] ), .D(
        n8853), .Z(n6463) );
  HS65_LH_NOR4ABX2 U9067 ( .A(n6465), .B(n6464), .C(n6463), .D(n6462), .Z(
        n6476) );
  HS65_LH_AO22X9 U9068 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][7] ), .B(n8940), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][7] ), .D(
        n8949), .Z(n6469) );
  HS65_LH_AO22X9 U9069 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][7] ), .B(n8939), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][7] ), .D(
        n9186), .Z(n6468) );
  HS65_LH_NAND4ABX3 U9070 ( .A(n6469), .B(n6468), .C(n6467), .D(n6466), .Z(
        n6475) );
  HS65_LH_NAND4ABX3 U9072 ( .A(n6473), .B(n6472), .C(n6471), .D(n6470), .Z(
        n6474) );
  HS65_LH_AOI22X1 U9073 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][11] ), .B(n8860), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][11] ), .D(
        n9192), .Z(n6503) );
  HS65_LH_AO22X9 U9074 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][11] ), .B(n9472), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][11] ), .D(
        n8857), .Z(n6501) );
  HS65_LH_AO22X9 U9075 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][11] ), .B(n9473), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][11] ), .D(
        n9474), .Z(n6500) );
  HS65_LH_NOR4ABX2 U9076 ( .A(n6503), .B(n6502), .C(n6501), .D(n6500), .Z(
        n6519) );
  HS65_LH_NOR4ABX2 U9077 ( .A(n6507), .B(n6506), .C(n6505), .D(n6504), .Z(
        n6518) );
  HS65_LH_AO22X9 U9078 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][11] ), .B(n8940), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][11] ), .D(
        n8949), .Z(n6511) );
  HS65_LH_AO22X9 U9079 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][11] ), .B(n8939), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][11] ), .D(
        n9186), .Z(n6510) );
  HS65_LH_NAND4ABX3 U9080 ( .A(n6511), .B(n6510), .C(n6509), .D(n6508), .Z(
        n6517) );
  HS65_LH_AO22X9 U9081 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][11] ), .B(n9470), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][11] ), .D(
        n9267), .Z(n6514) );
  HS65_LH_NAND4ABX3 U9082 ( .A(n6515), .B(n6514), .C(n6513), .D(n6512), .Z(
        n6516) );
  HS65_LH_AOI22X1 U9083 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][28] ), .B(n8860), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][28] ), .D(
        n9157), .Z(n6523) );
  HS65_LH_NOR4ABX2 U9085 ( .A(n6523), .B(n6522), .C(n6521), .D(n6520), .Z(
        n6542) );
  HS65_LH_AOI22X1 U9086 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][28] ), .B(n8950), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][28] ), .D(
        n8855), .Z(n6527) );
  HS65_LH_AO22X4 U9087 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][28] ), .B(n9187), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][28] ), .D(
        n9194), .Z(n6524) );
  HS65_LH_NOR4ABX2 U9088 ( .A(n6527), .B(n6526), .C(n6525), .D(n6524), .Z(
        n6541) );
  HS65_LH_BFX9 U9089 ( .A(n6529), .Z(n6916) );
  HS65_LH_AO22X9 U9090 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][28] ), .B(n9249), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][28] ), .D(
        n9185), .Z(n6534) );
  HS65_LH_NAND4ABX3 U9091 ( .A(n6534), .B(n6533), .C(n6532), .D(n6531), .Z(
        n6540) );
  HS65_LH_AO22X4 U9092 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][28] ), .B(n9470), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][28] ), .D(
        n9164), .Z(n6537) );
  HS65_LH_NAND4ABX3 U9093 ( .A(n6538), .B(n6537), .C(n6536), .D(n6535), .Z(
        n6539) );
  HS65_LH_AOI22X1 U9094 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][22] ), .B(n8860), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][22] ), .D(
        n9157), .Z(n6546) );
  HS65_LH_AO22X9 U9095 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][22] ), .B(n8858), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][22] ), .D(
        n9468), .Z(n6544) );
  HS65_LH_NOR4ABX2 U9096 ( .A(n6546), .B(n6545), .C(n6544), .D(n6543), .Z(
        n6562) );
  HS65_LH_AOI22X1 U9097 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][22] ), .B(n8950), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][22] ), .D(
        n8855), .Z(n6550) );
  HS65_LH_AO22X4 U9098 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][22] ), .B(n9187), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][22] ), .D(
        n9194), .Z(n6547) );
  HS65_LH_NOR4ABX2 U9099 ( .A(n6550), .B(n6549), .C(n6548), .D(n6547), .Z(
        n6561) );
  HS65_LH_AO22X9 U9100 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][22] ), .B(n9249), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][22] ), .D(
        n9185), .Z(n6554) );
  HS65_LH_NAND4ABX3 U9101 ( .A(n6554), .B(n6553), .C(n6552), .D(n6551), .Z(
        n6560) );
  HS65_LH_NAND4ABX3 U9102 ( .A(n6558), .B(n6557), .C(n6556), .D(n6555), .Z(
        n6559) );
  HS65_LH_AOI22X1 U9103 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][30] ), .B(n8860), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][30] ), .D(
        n9157), .Z(n6566) );
  HS65_LH_AO22X9 U9104 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][30] ), .B(n8858), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][30] ), .D(
        n9468), .Z(n6564) );
  HS65_LH_NOR4ABX2 U9105 ( .A(n6566), .B(n6565), .C(n6564), .D(n6563), .Z(
        n6582) );
  HS65_LH_AO22X4 U9106 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][30] ), .B(n9187), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][30] ), .D(
        n9194), .Z(n6567) );
  HS65_LH_NOR4ABX2 U9107 ( .A(n6570), .B(n6569), .C(n6568), .D(n6567), .Z(
        n6581) );
  HS65_LH_NAND4ABX3 U9109 ( .A(n6574), .B(n6573), .C(n6572), .D(n6571), .Z(
        n6580) );
  HS65_LH_NAND4ABX3 U9110 ( .A(n6578), .B(n6577), .C(n6576), .D(n6575), .Z(
        n6579) );
  HS65_LH_AOI22X1 U9111 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][20] ), .B(n8860), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][20] ), .D(
        n9157), .Z(n6586) );
  HS65_LH_NOR4ABX2 U9113 ( .A(n6586), .B(n6585), .C(n6584), .D(n6583), .Z(
        n6602) );
  HS65_LH_AOI22X1 U9114 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][20] ), .B(n8950), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][20] ), .D(
        n8855), .Z(n6590) );
  HS65_LH_AO22X4 U9115 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][20] ), .B(n9187), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][20] ), .D(
        n9194), .Z(n6587) );
  HS65_LH_NOR4ABX2 U9116 ( .A(n6590), .B(n6589), .C(n6588), .D(n6587), .Z(
        n6601) );
  HS65_LH_AO22X9 U9117 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][20] ), .B(n9249), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][20] ), .D(
        n9185), .Z(n6594) );
  HS65_LH_NAND4ABX3 U9119 ( .A(n6594), .B(n6593), .C(n6592), .D(n6591), .Z(
        n6600) );
  HS65_LH_NAND4ABX3 U9120 ( .A(n6598), .B(n6597), .C(n6596), .D(n6595), .Z(
        n6599) );
  HS65_LH_AOI22X1 U9121 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][31] ), .B(n8860), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][31] ), .D(
        n9157), .Z(n6606) );
  HS65_LH_NOR4ABX2 U9123 ( .A(n6606), .B(n6605), .C(n6604), .D(n6603), .Z(
        n6622) );
  HS65_LH_AOI22X1 U9124 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][31] ), .B(n8950), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][31] ), .D(
        n8855), .Z(n6610) );
  HS65_LH_AOI22X1 U9125 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][31] ), .B(n9162), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][31] ), .D(
        n8854), .Z(n6609) );
  HS65_LH_AO22X4 U9126 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][31] ), .B(n9187), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][31] ), .D(
        n9194), .Z(n6607) );
  HS65_LH_NOR4ABX2 U9127 ( .A(n6610), .B(n6609), .C(n6608), .D(n6607), .Z(
        n6621) );
  HS65_LH_AO22X9 U9128 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][31] ), .B(n9249), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][31] ), .D(
        n9185), .Z(n6614) );
  HS65_LH_NAND4ABX3 U9129 ( .A(n6614), .B(n6613), .C(n6612), .D(n6611), .Z(
        n6620) );
  HS65_LH_NAND4ABX3 U9130 ( .A(n6618), .B(n6617), .C(n6616), .D(n6615), .Z(
        n6619) );
  HS65_LH_AOI22X1 U9131 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][5] ), .B(n8860), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][5] ), .D(
        n9157), .Z(n6626) );
  HS65_LH_AO22X9 U9132 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][5] ), .B(n8858), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][5] ), .D(
        n9468), .Z(n6624) );
  HS65_LH_NOR4ABX2 U9133 ( .A(n6626), .B(n6625), .C(n6624), .D(n6623), .Z(
        n6643) );
  HS65_LH_AO22X4 U9134 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][5] ), .B(n9187), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][5] ), .D(
        n9194), .Z(n6627) );
  HS65_LH_NOR4ABX2 U9135 ( .A(n6630), .B(n6629), .C(n6628), .D(n6627), .Z(
        n6642) );
  HS65_LH_AO22X9 U9136 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][5] ), .B(n9249), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][5] ), .D(
        n9185), .Z(n6634) );
  HS65_LH_NAND4ABX3 U9137 ( .A(n6634), .B(n6633), .C(n6632), .D(n6631), .Z(
        n6641) );
  HS65_LH_NAND4ABX3 U9138 ( .A(n6639), .B(n6638), .C(n6637), .D(n6636), .Z(
        n6640) );
  HS65_LH_AOI22X1 U9139 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][8] ), .B(n8860), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][8] ), .D(
        n9192), .Z(n6647) );
  HS65_LH_NOR4ABX2 U9142 ( .A(n6647), .B(n6646), .C(n6645), .D(n6644), .Z(
        n6663) );
  HS65_LH_NOR4ABX2 U9143 ( .A(n6651), .B(n6650), .C(n6649), .D(n6648), .Z(
        n6662) );
  HS65_LH_NAND4ABX3 U9145 ( .A(n6655), .B(n6654), .C(n6653), .D(n6652), .Z(
        n6661) );
  HS65_LH_NAND4ABX3 U9147 ( .A(n6659), .B(n6658), .C(n6657), .D(n6656), .Z(
        n6660) );
  HS65_LH_AOI22X1 U9148 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][18] ), .B(n8860), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][18] ), .D(
        n9192), .Z(n6667) );
  HS65_LH_NOR4ABX2 U9151 ( .A(n6667), .B(n6666), .C(n6665), .D(n6664), .Z(
        n6683) );
  HS65_LH_NOR4ABX2 U9152 ( .A(n6671), .B(n6670), .C(n6669), .D(n6668), .Z(
        n6682) );
  HS65_LH_AO22X9 U9153 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][18] ), .B(n8939), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][18] ), .D(
        n9186), .Z(n6674) );
  HS65_LH_NAND4ABX3 U9154 ( .A(n6675), .B(n6674), .C(n6673), .D(n6672), .Z(
        n6681) );
  HS65_LH_AO22X9 U9155 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][18] ), .B(n9470), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][18] ), .D(
        n9267), .Z(n6678) );
  HS65_LH_NAND4ABX3 U9156 ( .A(n6679), .B(n6678), .C(n6677), .D(n6676), .Z(
        n6680) );
  HS65_LH_AOI22X1 U9157 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][12] ), .B(n8860), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][12] ), .D(
        n9192), .Z(n6687) );
  HS65_LH_AO22X9 U9158 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][12] ), .B(n9472), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][12] ), .D(
        n9468), .Z(n6685) );
  HS65_LH_AO22X9 U9159 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][12] ), .B(n9473), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][12] ), .D(
        n9474), .Z(n6684) );
  HS65_LH_NOR4ABX2 U9160 ( .A(n6687), .B(n6686), .C(n6685), .D(n6684), .Z(
        n6703) );
  HS65_LH_NOR4ABX2 U9161 ( .A(n6691), .B(n6690), .C(n6689), .D(n6688), .Z(
        n6702) );
  HS65_LH_AO22X9 U9162 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][12] ), .B(n8939), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][12] ), .D(
        n9186), .Z(n6694) );
  HS65_LH_NAND4ABX3 U9163 ( .A(n6695), .B(n6694), .C(n6693), .D(n6692), .Z(
        n6701) );
  HS65_LH_NAND4ABX3 U9165 ( .A(n6699), .B(n6698), .C(n6697), .D(n6696), .Z(
        n6700) );
  HS65_LH_AOI22X1 U9166 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][10] ), .B(n8860), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][10] ), .D(
        n9192), .Z(n6707) );
  HS65_LH_AO22X9 U9167 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][10] ), .B(n9472), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][10] ), .D(
        n9468), .Z(n6705) );
  HS65_LH_AO22X9 U9168 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][10] ), .B(n9473), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][10] ), .D(
        n9474), .Z(n6704) );
  HS65_LH_NOR4ABX2 U9169 ( .A(n6707), .B(n6706), .C(n6705), .D(n6704), .Z(
        n6723) );
  HS65_LH_NOR4ABX2 U9170 ( .A(n6711), .B(n6710), .C(n6709), .D(n6708), .Z(
        n6722) );
  HS65_LH_AO22X9 U9171 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][10] ), .B(n8939), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][10] ), .D(
        n9186), .Z(n6714) );
  HS65_LH_NAND4ABX3 U9172 ( .A(n6715), .B(n6714), .C(n6713), .D(n6712), .Z(
        n6721) );
  HS65_LH_NAND4ABX3 U9174 ( .A(n6719), .B(n6718), .C(n6717), .D(n6716), .Z(
        n6720) );
  HS65_LH_AOI22X1 U9175 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][6] ), .B(n8860), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][6] ), .D(
        n9192), .Z(n6731) );
  HS65_LH_AO22X9 U9176 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][6] ), .B(n9472), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][6] ), .D(
        n9468), .Z(n6729) );
  HS65_LH_AO22X9 U9177 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][6] ), .B(n9473), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][6] ), .D(
        n9474), .Z(n6728) );
  HS65_LH_NOR4ABX2 U9178 ( .A(n6731), .B(n6730), .C(n6729), .D(n6728), .Z(
        n6747) );
  HS65_LH_NOR4ABX2 U9179 ( .A(n6735), .B(n6734), .C(n6733), .D(n6732), .Z(
        n6746) );
  HS65_LH_AO22X9 U9180 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][6] ), .B(n8939), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][6] ), .D(
        n9186), .Z(n6738) );
  HS65_LH_NAND4ABX3 U9181 ( .A(n6739), .B(n6738), .C(n6737), .D(n6736), .Z(
        n6745) );
  HS65_LH_NAND4ABX3 U9183 ( .A(n6743), .B(n6742), .C(n6741), .D(n6740), .Z(
        n6744) );
  HS65_LH_NOR4ABX2 U9184 ( .A(n6764), .B(n6763), .C(n6762), .D(n6761), .Z(
        n6780) );
  HS65_LH_AO22X4 U9185 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][19] ), .B(n9364), 
        .C(n9253), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][19] ), .Z(n6766)
         );
  HS65_LH_NOR4ABX2 U9186 ( .A(n6768), .B(n6767), .C(n6766), .D(n6765), .Z(
        n6779) );
  HS65_LH_NAND4ABX3 U9187 ( .A(n6772), .B(n6771), .C(n6770), .D(n6769), .Z(
        n6778) );
  HS65_LH_NAND4ABX3 U9188 ( .A(n6776), .B(n6775), .C(n6774), .D(n6773), .Z(
        n6777) );
  HS65_LH_NOR4ABX2 U9189 ( .A(n6780), .B(n6779), .C(n6778), .D(n6777), .Z(
        n8067) );
  HS65_LH_NOR4ABX2 U9190 ( .A(n6784), .B(n6783), .C(n6782), .D(n6781), .Z(
        n6800) );
  HS65_LH_NOR4ABX2 U9191 ( .A(n6788), .B(n6787), .C(n6786), .D(n6785), .Z(
        n6799) );
  HS65_LH_NAND4ABX3 U9193 ( .A(n6792), .B(n6791), .C(n6790), .D(n6789), .Z(
        n6798) );
  HS65_LH_AO22X9 U9194 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][26] ), .B(n9363), 
        .C(n9257), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][26] ), .Z(n6796)
         );
  HS65_LH_NAND4ABX3 U9195 ( .A(n6796), .B(n6795), .C(n6794), .D(n6793), .Z(
        n6797) );
  HS65_LH_NOR4ABX2 U9196 ( .A(n6800), .B(n6799), .C(n6798), .D(n6797), .Z(
        n8248) );
  HS65_LH_NOR4ABX2 U9197 ( .A(n6804), .B(n6803), .C(n6802), .D(n6801), .Z(
        n6820) );
  HS65_LH_NOR4ABX2 U9198 ( .A(n6808), .B(n6807), .C(n6806), .D(n6805), .Z(
        n6819) );
  HS65_LH_AO22X9 U9199 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][11] ), .B(n9261), 
        .C(n9263), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][11] ), .Z(n6812)
         );
  HS65_LH_NAND4ABX3 U9200 ( .A(n6812), .B(n6811), .C(n6810), .D(n6809), .Z(
        n6818) );
  HS65_LH_AO22X9 U9201 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][11] ), .B(n9363), 
        .C(n9257), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][11] ), .Z(n6816)
         );
  HS65_LH_NAND4ABX3 U9202 ( .A(n6816), .B(n6815), .C(n6814), .D(n6813), .Z(
        n6817) );
  HS65_LH_NOR4ABX2 U9203 ( .A(n6820), .B(n6819), .C(n6818), .D(n6817), .Z(
        n8212) );
  HS65_LH_NOR4ABX2 U9204 ( .A(n6824), .B(n6823), .C(n6822), .D(n6821), .Z(
        n6840) );
  HS65_LH_NOR4ABX2 U9205 ( .A(n6828), .B(n6827), .C(n6826), .D(n6825), .Z(
        n6839) );
  HS65_LH_AO22X9 U9206 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][6] ), .B(n9261), 
        .C(n9263), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][6] ), .Z(n6832) );
  HS65_LH_NAND4ABX3 U9208 ( .A(n6832), .B(n6831), .C(n6830), .D(n6829), .Z(
        n6838) );
  HS65_LH_AO22X9 U9209 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][6] ), .B(n9363), 
        .C(n9257), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][6] ), .Z(n6836) );
  HS65_LH_NAND4ABX3 U9210 ( .A(n6836), .B(n6835), .C(n6834), .D(n6833), .Z(
        n6837) );
  HS65_LH_NOR4ABX2 U9211 ( .A(n6840), .B(n6839), .C(n6838), .D(n6837), .Z(
        n8244) );
  HS65_LH_NOR4ABX2 U9212 ( .A(n6844), .B(n6843), .C(n6842), .D(n6841), .Z(
        n6860) );
  HS65_LH_NOR4ABX2 U9213 ( .A(n6848), .B(n6847), .C(n6846), .D(n6845), .Z(
        n6859) );
  HS65_LH_AO22X9 U9214 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][8] ), .B(n9261), 
        .C(n9263), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][8] ), .Z(n6852) );
  HS65_LH_NAND4ABX3 U9216 ( .A(n6852), .B(n6851), .C(n6850), .D(n6849), .Z(
        n6858) );
  HS65_LH_AO22X9 U9217 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][8] ), .B(n9363), 
        .C(n9257), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][8] ), .Z(n6856) );
  HS65_LH_NAND4ABX3 U9218 ( .A(n6856), .B(n6855), .C(n6854), .D(n6853), .Z(
        n6857) );
  HS65_LH_NOR4ABX2 U9219 ( .A(n6860), .B(n6859), .C(n6858), .D(n6857), .Z(
        n8227) );
  HS65_LH_AO22X9 U9220 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][14] ), .B(n8858), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][14] ), .D(
        n9468), .Z(n6863) );
  HS65_LH_NOR4ABX2 U9221 ( .A(n6865), .B(n6864), .C(n6863), .D(n6862), .Z(
        n6881) );
  HS65_LH_AO22X9 U9222 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][14] ), .B(n9154), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][14] ), .D(
        n9194), .Z(n6866) );
  HS65_LH_NOR4ABX2 U9223 ( .A(n6869), .B(n6868), .C(n6867), .D(n6866), .Z(
        n6880) );
  HS65_LH_AO22X4 U9224 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][14] ), .B(n8940), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][14] ), .D(
        n8949), .Z(n6873) );
  HS65_LH_AO22X9 U9225 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][14] ), .B(n8939), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][14] ), .D(
        n9186), .Z(n6872) );
  HS65_LH_NAND4ABX3 U9226 ( .A(n6873), .B(n6872), .C(n6871), .D(n6870), .Z(
        n6879) );
  HS65_LH_NAND4ABX3 U9228 ( .A(n6877), .B(n6876), .C(n6875), .D(n6874), .Z(
        n6878) );
  HS65_LH_NOR4ABX2 U9229 ( .A(n6881), .B(n6880), .C(n6879), .D(n6878), .Z(
        n8254) );
  HS65_LH_AO22X9 U9230 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][15] ), .B(n8858), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][15] ), .D(
        n9468), .Z(n6883) );
  HS65_LH_NOR4ABX2 U9231 ( .A(n6885), .B(n6884), .C(n6883), .D(n6882), .Z(
        n6903) );
  HS65_LH_AOI22X1 U9232 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][15] ), .B(n9162), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][15] ), .D(
        n8854), .Z(n6888) );
  HS65_LH_AO22X4 U9233 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][15] ), .B(n9187), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][15] ), .D(
        n9194), .Z(n6886) );
  HS65_LH_NOR4ABX2 U9234 ( .A(n6889), .B(n6888), .C(n6887), .D(n6886), .Z(
        n6902) );
  HS65_LH_AO22X9 U9235 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][15] ), .B(n9249), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][15] ), .D(
        n9185), .Z(n6894) );
  HS65_LH_AO22X9 U9236 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][15] ), .B(n9251), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][15] ), .D(
        n9186), .Z(n6893) );
  HS65_LH_NAND4ABX3 U9237 ( .A(n6894), .B(n6893), .C(n6892), .D(n6891), .Z(
        n6901) );
  HS65_LH_NAND4ABX3 U9239 ( .A(n6899), .B(n6898), .C(n6897), .D(n6896), .Z(
        n6900) );
  HS65_LH_NOR4ABX2 U9240 ( .A(n6903), .B(n6902), .C(n6901), .D(n6900), .Z(
        n8303) );
  HS65_LH_AO22X9 U9241 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][29] ), .B(n8858), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][29] ), .D(
        n9468), .Z(n6905) );
  HS65_LH_NOR4ABX2 U9242 ( .A(n6907), .B(n6906), .C(n6905), .D(n6904), .Z(
        n6930) );
  HS65_LH_AOI22X1 U9243 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][29] ), .B(n9162), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][29] ), .D(
        n8854), .Z(n6914) );
  HS65_LH_AO22X4 U9244 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][29] ), .B(n9187), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][29] ), .D(
        n9194), .Z(n6912) );
  HS65_LH_NOR4ABX2 U9245 ( .A(n6915), .B(n6914), .C(n6913), .D(n6912), .Z(
        n6929) );
  HS65_LH_AO22X9 U9246 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][29] ), .B(n9249), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][29] ), .D(
        n9185), .Z(n6922) );
  HS65_LH_NAND4ABX3 U9248 ( .A(n6922), .B(n6921), .C(n6920), .D(n6919), .Z(
        n6928) );
  HS65_LH_NAND4ABX3 U9250 ( .A(n6926), .B(n6925), .C(n6924), .D(n6923), .Z(
        n6927) );
  HS65_LH_NOR4ABX2 U9251 ( .A(n6930), .B(n6929), .C(n6928), .D(n6927), .Z(
        n8319) );
  HS65_LH_AO22X9 U9252 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][26] ), .B(n8858), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][26] ), .D(
        n9468), .Z(n6932) );
  HS65_LH_NOR4ABX2 U9253 ( .A(n6934), .B(n6933), .C(n6932), .D(n6931), .Z(
        n6951) );
  HS65_LH_NOR4ABX2 U9254 ( .A(n6938), .B(n6937), .C(n6936), .D(n6935), .Z(
        n6950) );
  HS65_LH_AO22X9 U9255 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][26] ), .B(n8940), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][26] ), .D(
        n8949), .Z(n6942) );
  HS65_LH_AO22X9 U9256 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][26] ), .B(n8939), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][26] ), .D(
        n9186), .Z(n6941) );
  HS65_LH_NAND4ABX3 U9257 ( .A(n6942), .B(n6941), .C(n6940), .D(n6939), .Z(
        n6949) );
  HS65_LH_NAND4ABX3 U9259 ( .A(n6947), .B(n6946), .C(n6945), .D(n6944), .Z(
        n6948) );
  HS65_LH_NOR4ABX2 U9260 ( .A(n6951), .B(n6950), .C(n6949), .D(n6948), .Z(
        n8251) );
  HS65_LH_AO22X9 U9261 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][25] ), .B(n8858), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][25] ), .D(
        n9468), .Z(n6953) );
  HS65_LH_NOR4ABX2 U9262 ( .A(n6955), .B(n6954), .C(n6953), .D(n6952), .Z(
        n6971) );
  HS65_LH_NOR4ABX2 U9263 ( .A(n6959), .B(n6958), .C(n6957), .D(n6956), .Z(
        n6970) );
  HS65_LH_AO22X9 U9264 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][25] ), .B(n8939), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][25] ), .D(
        n9186), .Z(n6962) );
  HS65_LH_NAND4ABX3 U9265 ( .A(n6963), .B(n6962), .C(n6961), .D(n6960), .Z(
        n6969) );
  HS65_LH_AO22X9 U9266 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][25] ), .B(n9470), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][25] ), .D(
        n9164), .Z(n6966) );
  HS65_LH_NAND4ABX3 U9267 ( .A(n6967), .B(n6966), .C(n6965), .D(n6964), .Z(
        n6968) );
  HS65_LH_NOR4ABX2 U9268 ( .A(n6971), .B(n6970), .C(n6969), .D(n6968), .Z(
        n8256) );
  HS65_LH_AO22X9 U9269 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][9] ), .B(n8858), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][9] ), .D(
        n9468), .Z(n6979) );
  HS65_LH_NOR4ABX2 U9270 ( .A(n6981), .B(n6980), .C(n6979), .D(n6978), .Z(
        n7011) );
  HS65_LH_NOR4ABX2 U9271 ( .A(n6990), .B(n6989), .C(n6988), .D(n6987), .Z(
        n7010) );
  HS65_LH_NAND4ABX3 U9273 ( .A(n6997), .B(n6996), .C(n6995), .D(n6994), .Z(
        n7009) );
  HS65_LH_AO22X9 U9274 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][9] ), .B(n9470), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][9] ), .D(n9164), .Z(n7006) );
  HS65_LH_NAND4ABX3 U9275 ( .A(n7007), .B(n7006), .C(n7005), .D(n7004), .Z(
        n7008) );
  HS65_LH_NOR4ABX2 U9276 ( .A(n7011), .B(n7010), .C(n7009), .D(n7008), .Z(
        n8261) );
  HS65_LH_NAND3X2 U9277 ( .A(n9334), .B(n9209), .C(n9172), .Z(n8009) );
  HS65_LH_NOR2AX3 U9278 ( .A(n7015), .B(n7014), .Z(n7217) );
  HS65_LH_NAND2X2 U9279 ( .A(n8847), .B(n9173), .Z(n8011) );
  HS65_LH_NOR4ABX2 U9280 ( .A(n7019), .B(n7018), .C(n7017), .D(n7016), .Z(
        n7035) );
  HS65_LH_AO22X9 U9281 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][13] ), .B(n9364), 
        .C(n9253), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][13] ), .Z(n7021)
         );
  HS65_LH_NOR4ABX2 U9282 ( .A(n7023), .B(n7022), .C(n7021), .D(n7020), .Z(
        n7034) );
  HS65_LH_NAND4ABX3 U9283 ( .A(n7027), .B(n7026), .C(n7025), .D(n7024), .Z(
        n7033) );
  HS65_LH_NAND4ABX3 U9284 ( .A(n7031), .B(n7030), .C(n7029), .D(n7028), .Z(
        n7032) );
  HS65_LH_NOR4ABX2 U9285 ( .A(n7035), .B(n7034), .C(n7033), .D(n7032), .Z(
        n8153) );
  HS65_LH_NOR4ABX2 U9286 ( .A(n7039), .B(n7038), .C(n7037), .D(n7036), .Z(
        n7055) );
  HS65_LH_NOR4ABX2 U9288 ( .A(n7043), .B(n7042), .C(n7041), .D(n7040), .Z(
        n7054) );
  HS65_LH_NAND4ABX3 U9289 ( .A(n7047), .B(n7046), .C(n7045), .D(n7044), .Z(
        n7053) );
  HS65_LH_AOI22X1 U9290 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][10] ), .B(n9113), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][10] ), .D(
        n9166), .Z(n7048) );
  HS65_LH_NAND4ABX3 U9291 ( .A(n7051), .B(n7050), .C(n7049), .D(n7048), .Z(
        n7052) );
  HS65_LH_NOR4ABX2 U9292 ( .A(n7055), .B(n7054), .C(n7053), .D(n7052), .Z(
        n8062) );
  HS65_LH_NOR4ABX2 U9293 ( .A(n7059), .B(n7058), .C(n7057), .D(n7056), .Z(
        n7075) );
  HS65_LH_NOR4ABX2 U9294 ( .A(n7063), .B(n7062), .C(n7061), .D(n7060), .Z(
        n7074) );
  HS65_LH_AO22X9 U9295 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][9] ), .B(n9261), 
        .C(n9263), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][9] ), .Z(n7067) );
  HS65_LH_NAND4ABX3 U9296 ( .A(n7067), .B(n7066), .C(n7065), .D(n7064), .Z(
        n7073) );
  HS65_LH_NAND4ABX3 U9298 ( .A(n7071), .B(n7070), .C(n7069), .D(n7068), .Z(
        n7072) );
  HS65_LH_NOR4ABX2 U9299 ( .A(n7075), .B(n7074), .C(n7073), .D(n7072), .Z(
        n8257) );
  HS65_LH_NOR4ABX2 U9300 ( .A(n7079), .B(n7078), .C(n7077), .D(n7076), .Z(
        n7095) );
  HS65_LH_NOR4ABX2 U9301 ( .A(n7083), .B(n7082), .C(n7081), .D(n7080), .Z(
        n7094) );
  HS65_LH_AO22X9 U9302 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][5] ), .B(n9261), 
        .C(n9263), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][5] ), .Z(n7087) );
  HS65_LH_NAND4ABX3 U9303 ( .A(n7087), .B(n7086), .C(n7085), .D(n7084), .Z(
        n7093) );
  HS65_LH_AO22X9 U9304 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][5] ), .B(n9363), 
        .C(n9257), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][5] ), .Z(n7091) );
  HS65_LH_NAND4ABX3 U9305 ( .A(n7091), .B(n7090), .C(n7089), .D(n7088), .Z(
        n7092) );
  HS65_LH_NOR4ABX2 U9306 ( .A(n7095), .B(n7094), .C(n7093), .D(n7092), .Z(
        n8262) );
  HS65_LH_NOR4ABX2 U9307 ( .A(n7099), .B(n7098), .C(n7097), .D(n7096), .Z(
        n7115) );
  HS65_LH_NOR4ABX2 U9309 ( .A(n7103), .B(n7102), .C(n7101), .D(n7100), .Z(
        n7114) );
  HS65_LH_NAND4ABX3 U9311 ( .A(n7107), .B(n7106), .C(n7105), .D(n7104), .Z(
        n7113) );
  HS65_LH_NAND4ABX3 U9312 ( .A(n7111), .B(n7110), .C(n7109), .D(n7108), .Z(
        n7112) );
  HS65_LH_NOR4ABX2 U9313 ( .A(n7115), .B(n7114), .C(n7113), .D(n7112), .Z(
        n8274) );
  HS65_LH_NOR4ABX2 U9314 ( .A(n7119), .B(n7118), .C(n7117), .D(n7116), .Z(
        n7135) );
  HS65_LH_NOR4ABX2 U9315 ( .A(n7123), .B(n7122), .C(n7121), .D(n7120), .Z(
        n7134) );
  HS65_LH_NAND4ABX3 U9317 ( .A(n7127), .B(n7126), .C(n7125), .D(n7124), .Z(
        n7133) );
  HS65_LH_AO22X9 U9318 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][23] ), .B(n9363), 
        .C(n9257), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][23] ), .Z(n7131)
         );
  HS65_LH_NAND4ABX3 U9319 ( .A(n7131), .B(n7130), .C(n7129), .D(n7128), .Z(
        n7132) );
  HS65_LH_NOR4ABX2 U9320 ( .A(n7135), .B(n7134), .C(n7133), .D(n7132), .Z(
        n8208) );
  HS65_LH_NOR4ABX2 U9321 ( .A(n7139), .B(n7138), .C(n7137), .D(n7136), .Z(
        n7155) );
  HS65_LH_NOR4ABX2 U9322 ( .A(n7143), .B(n7142), .C(n7141), .D(n7140), .Z(
        n7154) );
  HS65_LH_NAND4ABX3 U9324 ( .A(n7147), .B(n7146), .C(n7145), .D(n7144), .Z(
        n7153) );
  HS65_LH_NAND4ABX3 U9325 ( .A(n7151), .B(n7150), .C(n7149), .D(n7148), .Z(
        n7152) );
  HS65_LH_NOR4ABX2 U9326 ( .A(n7155), .B(n7154), .C(n7153), .D(n7152), .Z(
        n8236) );
  HS65_LH_NOR4ABX2 U9327 ( .A(n7159), .B(n7158), .C(n7157), .D(n7156), .Z(
        n7175) );
  HS65_LH_NOR4ABX2 U9328 ( .A(n7163), .B(n7162), .C(n7161), .D(n7160), .Z(
        n7174) );
  HS65_LH_AO22X9 U9329 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][27] ), .B(n9261), 
        .C(n9263), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][27] ), .Z(n7167)
         );
  HS65_LH_NAND4ABX3 U9330 ( .A(n7167), .B(n7166), .C(n7165), .D(n7164), .Z(
        n7173) );
  HS65_LH_AO22X9 U9331 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][27] ), .B(n9363), 
        .C(n9257), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][27] ), .Z(n7171)
         );
  HS65_LH_NAND4ABX3 U9332 ( .A(n7171), .B(n7170), .C(n7169), .D(n7168), .Z(
        n7172) );
  HS65_LH_NOR4ABX2 U9333 ( .A(n7175), .B(n7174), .C(n7173), .D(n7172), .Z(
        n8204) );
  HS65_LH_NOR4ABX2 U9334 ( .A(n7179), .B(n7178), .C(n7177), .D(n7176), .Z(
        n7195) );
  HS65_LH_AO22X9 U9335 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][22] ), .B(n9364), 
        .C(n9068), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][22] ), .Z(n7181)
         );
  HS65_LH_NOR4ABX2 U9336 ( .A(n7183), .B(n7182), .C(n7181), .D(n7180), .Z(
        n7194) );
  HS65_LH_NAND4ABX3 U9338 ( .A(n7187), .B(n7186), .C(n7185), .D(n7184), .Z(
        n7193) );
  HS65_LH_NAND4ABX3 U9339 ( .A(n7191), .B(n7190), .C(n7189), .D(n7188), .Z(
        n7192) );
  HS65_LH_NOR4ABX2 U9340 ( .A(n7195), .B(n7194), .C(n7193), .D(n7192), .Z(
        n8272) );
  HS65_LH_NAND2X2 U9341 ( .A(n8847), .B(n9335), .Z(n8008) );
  HS65_LH_NOR4ABX2 U9342 ( .A(n7221), .B(n7220), .C(n7219), .D(n7218), .Z(
        n7237) );
  HS65_LH_AO22X9 U9343 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][18] ), .B(n9364), 
        .C(n9253), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][18] ), .Z(n7223)
         );
  HS65_LH_NOR4ABX2 U9344 ( .A(n7225), .B(n7224), .C(n7223), .D(n7222), .Z(
        n7236) );
  HS65_LH_NAND4ABX3 U9345 ( .A(n7229), .B(n7228), .C(n7227), .D(n7226), .Z(
        n7235) );
  HS65_LH_AOI22X1 U9346 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][18] ), .B(n9113), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][18] ), .D(
        n9166), .Z(n7230) );
  HS65_LH_NAND4ABX3 U9347 ( .A(n7233), .B(n7232), .C(n7231), .D(n7230), .Z(
        n7234) );
  HS65_LH_NOR4ABX2 U9348 ( .A(n7237), .B(n7236), .C(n7235), .D(n7234), .Z(
        n8061) );
  HS65_LH_NOR4ABX2 U9349 ( .A(n7241), .B(n7240), .C(n7239), .D(n7238), .Z(
        n7257) );
  HS65_LH_AO22X9 U9350 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][1] ), .B(n9364), 
        .C(n9253), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][1] ), .Z(n7243)
         );
  HS65_LH_NOR4ABX2 U9351 ( .A(n7245), .B(n7244), .C(n7243), .D(n7242), .Z(
        n7256) );
  HS65_LH_NAND4ABX3 U9352 ( .A(n7249), .B(n7248), .C(n7247), .D(n7246), .Z(
        n7255) );
  HS65_LH_AOI22X1 U9353 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][1] ), .B(n9113), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][1] ), .D(n9166), .Z(n7250) );
  HS65_LH_NAND4ABX3 U9354 ( .A(n7253), .B(n7252), .C(n7251), .D(n7250), .Z(
        n7254) );
  HS65_LH_NOR4ABX2 U9355 ( .A(n7257), .B(n7256), .C(n7255), .D(n7254), .Z(
        n8052) );
  HS65_LH_NOR4ABX2 U9356 ( .A(n7261), .B(n7260), .C(n7259), .D(n7258), .Z(
        n7277) );
  HS65_LH_NOR4ABX2 U9357 ( .A(n7265), .B(n7264), .C(n7263), .D(n7262), .Z(
        n7276) );
  HS65_LH_NAND4ABX3 U9358 ( .A(n7269), .B(n7268), .C(n7267), .D(n7266), .Z(
        n7275) );
  HS65_LH_AO22X4 U9359 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][15] ), .B(n9152), 
        .C(n9257), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][15] ), .Z(n7273)
         );
  HS65_LH_NAND4ABX3 U9360 ( .A(n7273), .B(n7272), .C(n7271), .D(n7270), .Z(
        n7274) );
  HS65_LH_NOR4ABX2 U9361 ( .A(n7277), .B(n7276), .C(n7275), .D(n7274), .Z(
        n8276) );
  HS65_LH_NOR4ABX2 U9362 ( .A(n7284), .B(n7283), .C(n7282), .D(n7281), .Z(
        n7301) );
  HS65_LH_NOR4ABX2 U9363 ( .A(n7288), .B(n7287), .C(n7286), .D(n7285), .Z(
        n7300) );
  HS65_LH_NAND4ABX3 U9365 ( .A(n7292), .B(n7291), .C(n7290), .D(n7289), .Z(
        n7299) );
  HS65_LH_AO22X4 U9366 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][0] ), .B(n9152), 
        .C(n9097), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][0] ), .Z(n7297) );
  HS65_LH_AO22X4 U9367 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][0] ), .B(n9070), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][0] ), .D(
        n9064), .Z(n7296) );
  HS65_LH_NAND4ABX3 U9368 ( .A(n7297), .B(n7296), .C(n7295), .D(n7294), .Z(
        n7298) );
  HS65_LH_NOR4ABX2 U9369 ( .A(n7301), .B(n7300), .C(n7299), .D(n7298), .Z(
        n8367) );
  HS65_LH_CNIVX3 U9370 ( .A(n8028), .Z(n8006) );
  HS65_LH_CNIVX3 U9371 ( .A(n8029), .Z(n8003) );
  HS65_LH_NAND2X2 U9373 ( .A(n7310), .B(n7309), .Z(n8013) );
  HS65_LH_NOR2X2 U9375 ( .A(\u_DataPath/cw_to_ex_i [0]), .B(n7315), .Z(
        \u_DataPath/u_execute/EXALU/N810 ) );
  HS65_LH_NAND2X2 U9376 ( .A(n7316), .B(n5148), .Z(n7319) );
  HS65_LH_NOR2X2 U9377 ( .A(n7316), .B(n5148), .Z(n7318) );
  HS65_LH_MUX21I1X3 U9378 ( .D0(n7319), .D1(n7318), .S0(n7317), .Z(n7326) );
  HS65_LH_NAND2X2 U9379 ( .A(n7320), .B(n5148), .Z(n7323) );
  HS65_LH_NOR2X2 U9380 ( .A(n7320), .B(n5148), .Z(n7322) );
  HS65_LH_MUX21I1X3 U9381 ( .D0(n7323), .D1(n7322), .S0(n7321), .Z(n7324) );
  HS65_LH_AOI22X1 U9382 ( .A(n7327), .B(n7326), .C(n7325), .D(n7324), .Z(n7328) );
  HS65_LH_NOR2X2 U9383 ( .A(\u_DataPath/cw_to_ex_i [0]), .B(n7328), .Z(
        \u_DataPath/u_execute/EXALU/N811 ) );
  HS65_LH_CNIVX3 U9384 ( .A(n7990), .Z(n7350) );
  HS65_LH_NOR2X2 U9385 ( .A(n8790), .B(n8791), .Z(n7348) );
  HS65_LH_NOR2X2 U9386 ( .A(\u_DataPath/immediate_ext_dec_i [3]), .B(
        \u_DataPath/immediate_ext_dec_i [6]), .Z(n7347) );
  HS65_LH_NOR3X1 U9387 ( .A(n8792), .B(n8817), .C(n8793), .Z(n7346) );
  HS65_LH_CNIVX3 U9395 ( .A(n7360), .Z(n7361) );
  HS65_LH_IVX9 U9396 ( .A(addr_to_iram_21), .Z(n7469) );
  HS65_LH_NOR2X6 U9397 ( .A(n7469), .B(n7381), .Z(n7365) );
  HS65_LH_CNIVX3 U9398 ( .A(n8020), .Z(n7395) );
  HS65_LH_AOI21X2 U9399 ( .A(opcode_i[0]), .B(n7395), .C(n7394), .Z(n7396) );
  HS65_LH_NAND2X2 U9400 ( .A(opcode_i[1]), .B(opcode_i[2]), .Z(n7399) );
  HS65_LH_CBI4I1X3 U9401 ( .A(opcode_i[0]), .B(n7404), .C(n7403), .D(n7411), 
        .Z(n7951) );
  HS65_LH_MUXI21X2 U9402 ( .D0(opcode_i[1]), .D1(opcode_i[2]), .S0(opcode_i[0]), .Z(n7607) );
  HS65_LH_NOR3X1 U9403 ( .A(n8802), .B(n8806), .C(n9422), .Z(n7987) );
  HS65_LH_IVX9 U9404 ( .A(n7422), .Z(n7624) );
  HS65_LH_IVX9 U9405 ( .A(n7428), .Z(n7437) );
  HS65_LH_CNIVX3 U9407 ( .A(n7431), .Z(n7432) );
  HS65_LH_NOR4ABX2 U9408 ( .A(n7479), .B(n7478), .C(n7477), .D(n7476), .Z(
        n7495) );
  HS65_LH_AO22X9 U9409 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][25] ), .B(n9364), 
        .C(n9253), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][25] ), .Z(n7481)
         );
  HS65_LH_NOR4ABX2 U9410 ( .A(n7483), .B(n7482), .C(n7481), .D(n7480), .Z(
        n7494) );
  HS65_LH_NAND4ABX3 U9411 ( .A(n7487), .B(n7486), .C(n7485), .D(n7484), .Z(
        n7493) );
  HS65_LH_AOI22X1 U9412 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][25] ), .B(n9113), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][25] ), .D(
        n9166), .Z(n7488) );
  HS65_LH_NAND4ABX3 U9413 ( .A(n7491), .B(n7490), .C(n7489), .D(n7488), .Z(
        n7492) );
  HS65_LH_NOR4ABX2 U9414 ( .A(n7495), .B(n7494), .C(n7493), .D(n7492), .Z(
        n8058) );
  HS65_LH_NOR4ABX2 U9415 ( .A(n7499), .B(n7498), .C(n7497), .D(n7496), .Z(
        n7526) );
  HS65_LH_NOR4ABX2 U9416 ( .A(n7507), .B(n7506), .C(n7505), .D(n7504), .Z(
        n7525) );
  HS65_LH_NAND4ABX3 U9417 ( .A(n7514), .B(n7513), .C(n7512), .D(n7511), .Z(
        n7524) );
  HS65_LH_NAND4ABX3 U9418 ( .A(n7522), .B(n7521), .C(n7520), .D(n7519), .Z(
        n7523) );
  HS65_LH_NOR4ABX2 U9419 ( .A(n7526), .B(n7525), .C(n7524), .D(n7523), .Z(
        n8039) );
  HS65_LH_AO22X9 U9421 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][30] ), .B(n9096), 
        .C(n9198), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][30] ), .Z(n7527)
         );
  HS65_LH_NOR4ABX2 U9422 ( .A(n7530), .B(n7529), .C(n7528), .D(n7527), .Z(
        n7546) );
  HS65_LH_NOR4ABX2 U9423 ( .A(n7534), .B(n7533), .C(n7532), .D(n7531), .Z(
        n7545) );
  HS65_LH_NAND4ABX3 U9424 ( .A(n7538), .B(n7537), .C(n7536), .D(n7535), .Z(
        n7544) );
  HS65_LH_NAND4ABX3 U9425 ( .A(n7542), .B(n7541), .C(n7540), .D(n7539), .Z(
        n7543) );
  HS65_LH_NOR4ABX2 U9426 ( .A(n7546), .B(n7545), .C(n7544), .D(n7543), .Z(
        n8271) );
  HS65_LH_AO22X9 U9427 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][29] ), .B(n9098), 
        .C(n9200), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][29] ), .Z(n7548)
         );
  HS65_LH_NOR4ABX2 U9428 ( .A(n7550), .B(n7549), .C(n7548), .D(n7547), .Z(
        n7568) );
  HS65_LH_NOR4ABX2 U9430 ( .A(n7554), .B(n7553), .C(n7552), .D(n7551), .Z(
        n7567) );
  HS65_LH_NAND4ABX3 U9431 ( .A(n7559), .B(n7558), .C(n7557), .D(n7556), .Z(
        n7566) );
  HS65_LH_NAND4ABX3 U9432 ( .A(n7564), .B(n7563), .C(n7562), .D(n7561), .Z(
        n7565) );
  HS65_LH_NOR4ABX2 U9433 ( .A(n7568), .B(n7567), .C(n7566), .D(n7565), .Z(
        n8269) );
  HS65_LH_AO22X9 U9434 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][28] ), .B(n9208), 
        .C(n9100), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][28] ), .Z(n7574)
         );
  HS65_LH_AO22X9 U9435 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][28] ), .B(n9096), 
        .C(n9158), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][28] ), .Z(n7573)
         );
  HS65_LH_NOR4ABX2 U9436 ( .A(n7576), .B(n7575), .C(n7574), .D(n7573), .Z(
        n7603) );
  HS65_LH_AO22X9 U9437 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][28] ), .B(n9261), 
        .C(n9263), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][28] ), .Z(n7582)
         );
  HS65_LH_NOR4ABX2 U9438 ( .A(n7584), .B(n7583), .C(n7582), .D(n7581), .Z(
        n7602) );
  HS65_LH_AOI22X1 U9440 ( .A(n9161), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][28] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][28] ), .D(n9095), 
        .Z(n7590) );
  HS65_LH_NAND4ABX3 U9441 ( .A(n7592), .B(n7591), .C(n7590), .D(n7589), .Z(
        n7601) );
  HS65_LH_NAND4ABX3 U9442 ( .A(n7599), .B(n7598), .C(n7597), .D(n7596), .Z(
        n7600) );
  HS65_LH_NOR4ABX2 U9443 ( .A(n7603), .B(n7602), .C(n7601), .D(n7600), .Z(
        n8268) );
  HS65_LH_CNIVX3 U9444 ( .A(\u_DataPath/immediate_ext_dec_i [4]), .Z(n7604) );
  HS65_LH_NAND4ABX3 U9445 ( .A(n8801), .B(n8806), .C(n8817), .D(n9179), .Z(
        n7968) );
  HS65_LH_CNIVX3 U9446 ( .A(n7607), .Z(n7610) );
  HS65_LH_AOI21X2 U9447 ( .A(n7611), .B(n7610), .C(n7609), .Z(n7612) );
  HS65_LH_AOI21X2 U9448 ( .A(n7615), .B(n7614), .C(n8321), .Z(n7993) );
  HS65_LHS_XOR2X3 U9449 ( .A(n9293), .B(n7633), .Z(
        \u_DataPath/u_execute/link_value_i [27]) );
  HS65_LHS_XOR2X3 U9450 ( .A(n9458), .B(n7635), .Z(
        \u_DataPath/u_execute/link_value_i [25]) );
  HS65_LL_OAI21X12 U9452 ( .A(n8726), .B(n8014), .C(n1885), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N125 ) );
  HS65_LL_OAI21X12 U9453 ( .A(n3532), .B(n8014), .C(n1885), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N128 ) );
  HS65_LL_OAI21X12 U9454 ( .A(n7644), .B(n8014), .C(n1885), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N129 ) );
  HS65_LL_AOI22X1 U9455 ( .A(n8313), .B(n9429), .C(n7695), .D(
        \u_DataPath/u_execute/link_value_i [24]), .Z(n7662) );
  HS65_LL_NOR4ABX2 U9456 ( .A(n9052), .B(n7949), .C(n8798), .D(n8802), .Z(
        n7996) );
  HS65_LL_AO222X9 U9457 ( .A(n8352), .B(n8315), .C(n7695), .D(
        \u_DataPath/u_execute/link_value_i [16]), .E(n9137), .F(n8313), .Z(
        \u_DataPath/dataOut_exe_i [16]) );
  HS65_LH_AO222X4 U9458 ( .A(n7706), .B(n8961), .C(n7691), .D(n8614), .E(n8876), .F(n7685), .Z(addr_to_iram_24) );
  HS65_LH_AO222X4 U9459 ( .A(n7706), .B(n9017), .C(n7690), .D(n8617), .E(n8840), .F(n7685), .Z(addr_to_iram_20) );
  HS65_LH_AO222X4 U9460 ( .A(n7706), .B(n8962), .C(n7690), .D(n9377), .E(n8836), .F(n7685), .Z(addr_to_iram_18) );
  HS65_LH_AND2X4 U9461 ( .A(n1885), .B(n8967), .Z(
        \u_DataPath/pc4_to_idexreg_i [29]) );
  HS65_LH_NAND3X2 U9462 ( .A(n1885), .B(n8563), .C(n9445), .Z(n8280) );
  HS65_LH_AND2X4 U9463 ( .A(n1885), .B(\u_DataPath/toPC2_i [24]), .Z(
        \u_DataPath/branch_target_i [24]) );
  HS65_LH_NOR4ABX2 U9464 ( .A(n8441), .B(n8386), .C(n8385), .D(n8384), .Z(
        \u_DataPath/mem_writedata_out_i [5]) );
  HS65_LH_NOR4ABX2 U9465 ( .A(n8441), .B(n8416), .C(n8415), .D(n8414), .Z(
        \u_DataPath/mem_writedata_out_i [14]) );
  HS65_LH_NOR4ABX2 U9466 ( .A(n8441), .B(n8428), .C(n8427), .D(n8426), .Z(
        \u_DataPath/mem_writedata_out_i [18]) );
  HS65_LH_NOR4ABX2 U9467 ( .A(n8441), .B(n8440), .C(n8439), .D(n8438), .Z(
        \u_DataPath/mem_writedata_out_i [22]) );
  HS65_LH_NOR4ABX2 U9468 ( .A(n8441), .B(n8431), .C(n8430), .D(n8429), .Z(
        \u_DataPath/mem_writedata_out_i [19]) );
  HS65_LH_NOR4ABX2 U9469 ( .A(n8441), .B(n8422), .C(n8421), .D(n8420), .Z(
        \u_DataPath/mem_writedata_out_i [16]) );
  HS65_LH_NAND2X7 U9470 ( .A(n8728), .B(n8186), .Z(n8317) );
  HS65_LH_AND2X4 U9471 ( .A(n1885), .B(\u_DataPath/toPC2_i [15]), .Z(
        \u_DataPath/branch_target_i [15]) );
  HS65_LH_NOR3AX4 U9472 ( .A(n8752), .B(rst), .C(n9445), .Z(n8313) );
  HS65_LH_NOR4ABX2 U9473 ( .A(n8441), .B(n8392), .C(n8391), .D(n8390), .Z(
        \u_DataPath/mem_writedata_out_i [7]) );
  HS65_LH_NOR4ABX2 U9474 ( .A(n8441), .B(n8419), .C(n8418), .D(n8417), .Z(
        \u_DataPath/mem_writedata_out_i [15]) );
  HS65_LH_NOR4ABX2 U9475 ( .A(n8413), .B(n8412), .C(rst), .D(n8411), .Z(
        \u_DataPath/mem_writedata_out_i [13]) );
  HS65_LH_NOR4ABX2 U9476 ( .A(n8425), .B(n8424), .C(n8423), .D(rst), .Z(
        \u_DataPath/mem_writedata_out_i [17]) );
  HS65_LH_NOR4ABX2 U9477 ( .A(n8395), .B(n8394), .C(n8393), .D(rst), .Z(
        \u_DataPath/mem_writedata_out_i [8]) );
  HS65_LH_NOR4ABX2 U9478 ( .A(n8402), .B(n8401), .C(n8400), .D(rst), .Z(
        \u_DataPath/mem_writedata_out_i [10]) );
  HS65_LH_NOR4ABX2 U9479 ( .A(n8380), .B(n8379), .C(n7670), .D(rst), .Z(
        \u_DataPath/mem_writedata_out_i [3]) );
  HS65_LH_NOR4ABX2 U9480 ( .A(n8441), .B(n8434), .C(n8433), .D(n8432), .Z(
        \u_DataPath/mem_writedata_out_i [20]) );
  HS65_LH_NOR4ABX2 U9481 ( .A(n8441), .B(n8437), .C(n8436), .D(n8435), .Z(
        \u_DataPath/mem_writedata_out_i [21]) );
  HS65_LH_AND2X4 U9482 ( .A(n1885), .B(\u_DataPath/toPC2_i [22]), .Z(
        \u_DataPath/branch_target_i [22]) );
  HS65_LH_AND2X4 U9483 ( .A(n1885), .B(\u_DataPath/toPC2_i [19]), .Z(
        \u_DataPath/branch_target_i [19]) );
  HS65_LH_AND2X4 U9484 ( .A(n1885), .B(\u_DataPath/toPC2_i [18]), .Z(
        \u_DataPath/branch_target_i [18]) );
  HS65_LH_AND2X4 U9485 ( .A(n1885), .B(\u_DataPath/toPC2_i [17]), .Z(
        \u_DataPath/branch_target_i [17]) );
  HS65_LH_AND2X4 U9486 ( .A(n1885), .B(\u_DataPath/toPC2_i [20]), .Z(
        \u_DataPath/branch_target_i [20]) );
  HS65_LH_AND2X4 U9487 ( .A(n1885), .B(n9019), .Z(
        \u_DataPath/pc4_to_idexreg_i [16]) );
  HS65_LH_NOR3AX2 U9488 ( .A(n8994), .B(n9063), .C(n8071), .Z(
        \u_DataPath/cw_exmem_i [9]) );
  HS65_LH_NOR4ABX2 U9489 ( .A(n8799), .B(n8817), .C(n7973), .D(n8363), .Z(
        n7997) );
  HS65_LH_NAND3X2 U9490 ( .A(n8007), .B(n9058), .C(n9061), .Z(n8014) );
  HS65_LH_NOR2X2 U9491 ( .A(n9066), .B(rst), .Z(n8007) );
  HS65_LH_BFX4 U9492 ( .A(n8502), .Z(n7923) );
  HS65_LH_BFX4 U9493 ( .A(n8475), .Z(n7756) );
  HS65_LH_BFX4 U9494 ( .A(n8503), .Z(n7927) );
  HS65_LH_BFX4 U9495 ( .A(n8503), .Z(n7926) );
  HS65_LH_BFX4 U9496 ( .A(n8502), .Z(n7925) );
  HS65_LH_BFX4 U9497 ( .A(n8475), .Z(n7757) );
  HS65_LH_BFX4 U9498 ( .A(n8475), .Z(n7758) );
  HS65_LH_CNIVX3 U9499 ( .A(n8226), .Z(n8475) );
  HS65_LH_BFX4 U9500 ( .A(n8501), .Z(n7922) );
  HS65_LH_BFX4 U9501 ( .A(n8503), .Z(n7928) );
  HS65_LH_CNIVX3 U9502 ( .A(n8282), .Z(n8503) );
  HS65_LH_BFX4 U9503 ( .A(n8502), .Z(n7924) );
  HS65_LH_CNIVX3 U9504 ( .A(n8298), .Z(n8502) );
  HS65_LH_BFX4 U9505 ( .A(n8501), .Z(n7920) );
  HS65_LH_BFX4 U9506 ( .A(n8501), .Z(n7921) );
  HS65_LH_CNIVX3 U9507 ( .A(n8055), .Z(n8501) );
  HS65_LH_AND2X4 U9508 ( .A(n1885), .B(n8871), .Z(
        \u_DataPath/branch_target_i [1]) );
  HS65_LH_AND2X4 U9509 ( .A(n1885), .B(n9387), .Z(
        \u_DataPath/pc4_to_idexreg_i [2]) );
  HS65_LH_NOR4ABX2 U9510 ( .A(n8441), .B(n8374), .C(n8373), .D(n8372), .Z(
        \u_DataPath/mem_writedata_out_i [1]) );
  HS65_LH_AND2X4 U9511 ( .A(n1885), .B(\u_DataPath/toPC2_i [2]), .Z(
        \u_DataPath/branch_target_i [2]) );
  HS65_LH_NOR4ABX2 U9512 ( .A(n8383), .B(n8382), .C(n8381), .D(rst), .Z(
        \u_DataPath/mem_writedata_out_i [4]) );
  HS65_LH_NOR4ABX2 U9513 ( .A(n8405), .B(n8404), .C(n8403), .D(rst), .Z(
        \u_DataPath/mem_writedata_out_i [11]) );
  HS65_LH_NOR4ABX2 U9514 ( .A(n8371), .B(n8370), .C(n8369), .D(rst), .Z(
        \u_DataPath/mem_writedata_out_i [0]) );
  HS65_LH_NOR4ABX2 U9515 ( .A(n8389), .B(n8388), .C(n8387), .D(rst), .Z(
        \u_DataPath/mem_writedata_out_i [6]) );
  HS65_LH_AO222X4 U9516 ( .A(n7707), .B(n8997), .C(n7689), .D(n8616), .E(n9365), .F(n7687), .Z(addr_to_iram_1) );
  HS65_LH_AND2X4 U9517 ( .A(n1885), .B(\u_DataPath/toPC2_i [5]), .Z(
        \u_DataPath/branch_target_i [5]) );
  HS65_LH_AND2X4 U9518 ( .A(n1885), .B(n9099), .Z(
        \u_DataPath/pc4_to_idexreg_i [6]) );
  HS65_LH_AND2X4 U9519 ( .A(n1885), .B(\u_DataPath/toPC2_i [6]), .Z(
        \u_DataPath/branch_target_i [6]) );
  HS65_LH_AND2X4 U9520 ( .A(n1885), .B(\u_DataPath/toPC2_i [8]), .Z(
        \u_DataPath/branch_target_i [8]) );
  HS65_LH_AND2X4 U9521 ( .A(n1885), .B(n9015), .Z(
        \u_DataPath/pc4_to_idexreg_i [12]) );
  HS65_LH_AND2X4 U9522 ( .A(n1885), .B(n8955), .Z(
        \u_DataPath/pc4_to_idexreg_i [25]) );
  HS65_LH_AND2X4 U9523 ( .A(n1885), .B(\u_DataPath/toPC2_i [13]), .Z(
        \u_DataPath/branch_target_i [13]) );
  HS65_LH_AND2X4 U9524 ( .A(n1885), .B(n9078), .Z(
        \u_DataPath/pc4_to_idexreg_i [18]) );
  HS65_LH_AND2X4 U9525 ( .A(n1885), .B(\u_DataPath/toPC2_i [11]), .Z(
        \u_DataPath/branch_target_i [11]) );
  HS65_LH_AND2X4 U9526 ( .A(n1885), .B(\u_DataPath/toPC2_i [12]), .Z(
        \u_DataPath/branch_target_i [12]) );
  HS65_LH_OAI12X6 U9527 ( .A(n8846), .B(n8012), .C(n1885), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N139 ) );
  HS65_LH_OAI12X6 U9528 ( .A(n8011), .B(n8012), .C(n1885), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N138 ) );
  HS65_LH_OAI12X6 U9529 ( .A(n8008), .B(n8012), .C(n1885), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N134 ) );
  HS65_LH_OAI12X6 U9530 ( .A(n8008), .B(n8014), .C(n1885), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N126 ) );
  HS65_LH_OAI12X6 U9531 ( .A(n8004), .B(n8008), .C(n1885), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N150 ) );
  HS65_LH_OAI12X6 U9532 ( .A(n8846), .B(n8014), .C(n1885), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N131 ) );
  HS65_LH_OAI12X6 U9533 ( .A(n8011), .B(n8014), .C(n1885), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N130 ) );
  HS65_LH_OAI12X6 U9534 ( .A(n8011), .B(n8004), .C(n1885), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N154 ) );
  HS65_LH_OAI12X6 U9535 ( .A(n8011), .B(n8005), .C(n1885), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N146 ) );
  HS65_LH_OAI12X6 U9536 ( .A(n8005), .B(n8846), .C(n1885), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N147 ) );
  HS65_LH_NAND3X5 U9537 ( .A(n9184), .B(n9233), .C(n8007), .Z(n8012) );
  HS65_LH_OAI12X6 U9538 ( .A(n8005), .B(n8008), .C(n1885), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N142 ) );
  HS65_LH_NAND3X5 U9539 ( .A(n9270), .B(n9183), .C(n8007), .Z(n8005) );
  HS65_LH_CNIVX3 U9540 ( .A(n7742), .Z(n7748) );
  HS65_LH_CNIVX3 U9541 ( .A(n7906), .Z(n7911) );
  HS65_LH_CNIVX3 U9542 ( .A(n7836), .Z(n7841) );
  HS65_LH_CNIVX3 U9543 ( .A(n7766), .Z(n7771) );
  HS65_LH_CNIVX3 U9544 ( .A(n7878), .Z(n7883) );
  HS65_LH_CNIVX3 U9545 ( .A(n7885), .Z(n7890) );
  HS65_LH_CNIVX3 U9546 ( .A(n7787), .Z(n7792) );
  HS65_LH_CNIVX3 U9547 ( .A(n7815), .Z(n7820) );
  HS65_LH_CNIVX3 U9548 ( .A(n7871), .Z(n7876) );
  HS65_LH_CNIVX3 U9549 ( .A(n7749), .Z(n7754) );
  HS65_LH_CNIVX3 U9550 ( .A(n7801), .Z(n7806) );
  HS65_LH_CNIVX3 U9551 ( .A(n7794), .Z(n7799) );
  HS65_LH_CNIVX3 U9552 ( .A(n7822), .Z(n7828) );
  HS65_LH_CNIVX3 U9553 ( .A(n7735), .Z(n7741) );
  HS65_LH_CNIVX3 U9554 ( .A(n7857), .Z(n7863) );
  HS65_LH_CNIVX3 U9555 ( .A(n7864), .Z(n7870) );
  HS65_LH_CNIVX3 U9556 ( .A(n7780), .Z(n7786) );
  HS65_LH_CNIVX3 U9557 ( .A(n7892), .Z(n7898) );
  HS65_LH_CNIVX3 U9558 ( .A(n7728), .Z(n7734) );
  HS65_LH_CNIVX3 U9559 ( .A(n7850), .Z(n7856) );
  HS65_LH_CNIVX3 U9560 ( .A(n7843), .Z(n7849) );
  HS65_LH_CNIVX3 U9561 ( .A(n7759), .Z(n7765) );
  HS65_LH_CNIVX3 U9562 ( .A(n7773), .Z(n7779) );
  HS65_LH_CNIVX3 U9563 ( .A(n7899), .Z(n7905) );
  HS65_LH_CNIVX3 U9564 ( .A(n7906), .Z(n7912) );
  HS65_LH_CNIVX3 U9565 ( .A(n7836), .Z(n7842) );
  HS65_LH_CNIVX3 U9566 ( .A(n7766), .Z(n7772) );
  HS65_LH_CNIVX3 U9567 ( .A(n7878), .Z(n7884) );
  HS65_LH_CNIVX3 U9568 ( .A(n7885), .Z(n7891) );
  HS65_LH_CNIVX3 U9569 ( .A(n7787), .Z(n7793) );
  HS65_LH_CNIVX3 U9570 ( .A(n7815), .Z(n7821) );
  HS65_LH_CNIVX3 U9571 ( .A(n7871), .Z(n7877) );
  HS65_LH_CNIVX3 U9572 ( .A(n7749), .Z(n7755) );
  HS65_LH_CNIVX3 U9573 ( .A(n7899), .Z(n7904) );
  HS65_LH_CNIVX3 U9574 ( .A(n7801), .Z(n7807) );
  HS65_LH_CNIVX3 U9575 ( .A(n7794), .Z(n7800) );
  HS65_LH_CNIVX3 U9576 ( .A(n7913), .Z(n7918) );
  HS65_LH_CNIVX3 U9577 ( .A(n7913), .Z(n7919) );
  HS65_LH_CNIVX3 U9578 ( .A(n7721), .Z(n7726) );
  HS65_LH_CNIVX3 U9579 ( .A(n7721), .Z(n7727) );
  HS65_LH_CNIVX3 U9580 ( .A(n7829), .Z(n7835) );
  HS65_LH_CNIVX3 U9581 ( .A(n7773), .Z(n7778) );
  HS65_LH_CNIVX3 U9582 ( .A(n7759), .Z(n7764) );
  HS65_LH_CNIVX3 U9583 ( .A(n7808), .Z(n7814) );
  HS65_LH_CNIVX3 U9584 ( .A(n7882), .Z(n7881) );
  HS65_LH_CNIVX3 U9585 ( .A(n7843), .Z(n7848) );
  HS65_LH_CNIVX3 U9586 ( .A(n7850), .Z(n7855) );
  HS65_LH_CNIVX3 U9587 ( .A(n7791), .Z(n7790) );
  HS65_LH_CNIVX3 U9588 ( .A(n7854), .Z(n7853) );
  HS65_LH_CNIVX3 U9589 ( .A(n7728), .Z(n7733) );
  HS65_LH_CNIVX3 U9590 ( .A(n7875), .Z(n7874) );
  HS65_LH_CNIVX3 U9591 ( .A(n7732), .Z(n7731) );
  HS65_LH_CNIVX3 U9592 ( .A(n7753), .Z(n7752) );
  HS65_LH_CNIVX3 U9593 ( .A(n7892), .Z(n7897) );
  HS65_LH_CNIVX3 U9594 ( .A(n7798), .Z(n7797) );
  HS65_LH_CNIVX3 U9595 ( .A(n7896), .Z(n7895) );
  HS65_LH_CNIVX3 U9596 ( .A(n7780), .Z(n7785) );
  HS65_LH_CNIVX3 U9597 ( .A(n7784), .Z(n7783) );
  HS65_LH_CNIVX3 U9598 ( .A(n7808), .Z(n7813) );
  HS65_LH_CNIVX3 U9599 ( .A(n7864), .Z(n7869) );
  HS65_LH_CNIVX3 U9600 ( .A(n7861), .Z(n7860) );
  HS65_LH_CNIVX3 U9601 ( .A(n7829), .Z(n7834) );
  HS65_LH_CNIVX3 U9602 ( .A(n7857), .Z(n7862) );
  HS65_LH_CNIVX3 U9603 ( .A(n7903), .Z(n7902) );
  HS65_LH_CNIVX3 U9604 ( .A(n7822), .Z(n7827) );
  HS65_LH_CNIVX3 U9605 ( .A(n7735), .Z(n7740) );
  HS65_LH_CNIVX3 U9606 ( .A(n7742), .Z(n7747) );
  HS65_LH_CNIVX3 U9607 ( .A(n8042), .Z(\u_DataPath/u_execute/psw_status_i [1])
         );
  HS65_LH_CNIVX3 U9610 ( .A(n8154), .Z(\u_DataPath/cw_memwb_i [1]) );
  HS65_LH_CNIVX3 U9611 ( .A(n8366), .Z(\u_DataPath/reg_write_i ) );
  HS65_LL_NAND2X2 U9612 ( .A(n7945), .B(n8513), .Z(n7946) );
  HS65_LH_IVX9 U9613 ( .A(n8071), .Z(n8023) );
  HS65_LH_NOR2X6 U9614 ( .A(n8802), .B(n7962), .Z(n7991) );
  HS65_LH_IVX9 U9615 ( .A(n7949), .Z(n7962) );
  HS65_LH_NOR2AX3 U9616 ( .A(n9351), .B(rst), .Z(n8184) );
  HS65_LH_CNIVX3 U9618 ( .A(n7748), .Z(n7743) );
  HS65_LH_CNIVX3 U9619 ( .A(n7911), .Z(n7908) );
  HS65_LH_CNIVX3 U9620 ( .A(n7841), .Z(n7838) );
  HS65_LH_CNIVX3 U9621 ( .A(n7771), .Z(n7768) );
  HS65_LH_CNIVX3 U9622 ( .A(n7883), .Z(n7880) );
  HS65_LH_CNIVX3 U9623 ( .A(n7890), .Z(n7887) );
  HS65_LH_CNIVX3 U9624 ( .A(n7792), .Z(n7789) );
  HS65_LH_CNIVX3 U9625 ( .A(n7820), .Z(n7817) );
  HS65_LH_CNIVX3 U9626 ( .A(n7876), .Z(n7873) );
  HS65_LH_CNIVX3 U9627 ( .A(n7754), .Z(n7751) );
  HS65_LH_CNIVX3 U9628 ( .A(n7806), .Z(n7803) );
  HS65_LH_CNIVX3 U9629 ( .A(n7799), .Z(n7796) );
  HS65_LH_CNIVX3 U9630 ( .A(n7828), .Z(n7823) );
  HS65_LH_CNIVX3 U9631 ( .A(n7741), .Z(n7736) );
  HS65_LH_CNIVX3 U9632 ( .A(n7863), .Z(n7858) );
  HS65_LH_CNIVX3 U9633 ( .A(n7870), .Z(n7865) );
  HS65_LH_CNIVX3 U9634 ( .A(n7786), .Z(n7781) );
  HS65_LH_CNIVX3 U9635 ( .A(n7898), .Z(n7893) );
  HS65_LH_CNIVX3 U9636 ( .A(n7734), .Z(n7729) );
  HS65_LH_CNIVX3 U9637 ( .A(n7856), .Z(n7851) );
  HS65_LH_CNIVX3 U9638 ( .A(n7849), .Z(n7844) );
  HS65_LH_CNIVX3 U9639 ( .A(n7765), .Z(n7760) );
  HS65_LH_CNIVX3 U9640 ( .A(n7779), .Z(n7774) );
  HS65_LH_CNIVX3 U9641 ( .A(n7905), .Z(n7900) );
  HS65_LH_CNIVX3 U9642 ( .A(n7912), .Z(n7907) );
  HS65_LH_CNIVX3 U9643 ( .A(n7842), .Z(n7837) );
  HS65_LH_CNIVX3 U9644 ( .A(n7772), .Z(n7767) );
  HS65_LH_CNIVX3 U9645 ( .A(n7884), .Z(n7879) );
  HS65_LH_CNIVX3 U9646 ( .A(n7891), .Z(n7886) );
  HS65_LH_CNIVX3 U9647 ( .A(n7793), .Z(n7788) );
  HS65_LH_CNIVX3 U9648 ( .A(n7821), .Z(n7816) );
  HS65_LH_CNIVX3 U9649 ( .A(n7877), .Z(n7872) );
  HS65_LH_CNIVX3 U9650 ( .A(n7755), .Z(n7750) );
  HS65_LH_CNIVX3 U9651 ( .A(n7904), .Z(n7901) );
  HS65_LH_CNIVX3 U9652 ( .A(n7807), .Z(n7802) );
  HS65_LH_CNIVX3 U9653 ( .A(n7800), .Z(n7795) );
  HS65_LH_CNIVX3 U9654 ( .A(n7918), .Z(n7915) );
  HS65_LH_CNIVX3 U9655 ( .A(n7919), .Z(n7914) );
  HS65_LH_CNIVX3 U9656 ( .A(n7726), .Z(n7723) );
  HS65_LH_CNIVX3 U9657 ( .A(n7727), .Z(n7722) );
  HS65_LH_CNIVX3 U9658 ( .A(n7910), .Z(n7909) );
  HS65_LH_CNIVX3 U9659 ( .A(n7835), .Z(n7830) );
  HS65_LH_CNIVX3 U9660 ( .A(n7868), .Z(n7867) );
  HS65_LH_CNIVX3 U9661 ( .A(n7778), .Z(n7775) );
  HS65_LH_CNIVX3 U9662 ( .A(n7777), .Z(n7776) );
  HS65_LH_CNIVX3 U9663 ( .A(n7764), .Z(n7761) );
  HS65_LH_CNIVX3 U9664 ( .A(n7763), .Z(n7762) );
  HS65_LH_CNIVX3 U9665 ( .A(n7840), .Z(n7839) );
  HS65_LH_CNIVX3 U9666 ( .A(n7814), .Z(n7809) );
  HS65_LH_CNIVX3 U9667 ( .A(n7770), .Z(n7769) );
  HS65_LH_CNIVX3 U9668 ( .A(n7848), .Z(n7845) );
  HS65_LH_CNIVX3 U9669 ( .A(n7889), .Z(n7888) );
  HS65_LH_CNIVX3 U9670 ( .A(n7847), .Z(n7846) );
  HS65_LH_CNIVX3 U9671 ( .A(n7855), .Z(n7852) );
  HS65_LH_CNIVX3 U9672 ( .A(n7819), .Z(n7818) );
  HS65_LH_CNIVX3 U9673 ( .A(n7733), .Z(n7730) );
  HS65_LH_CNIVX3 U9674 ( .A(n7805), .Z(n7804) );
  HS65_LH_CNIVX3 U9675 ( .A(n7897), .Z(n7894) );
  HS65_LH_CNIVX3 U9676 ( .A(n7785), .Z(n7782) );
  HS65_LH_CNIVX3 U9677 ( .A(n7725), .Z(n7724) );
  HS65_LH_CNIVX3 U9678 ( .A(n7813), .Z(n7810) );
  HS65_LH_CNIVX3 U9679 ( .A(n7869), .Z(n7866) );
  HS65_LH_CNIVX3 U9680 ( .A(n7812), .Z(n7811) );
  HS65_LH_CNIVX3 U9681 ( .A(n7834), .Z(n7831) );
  HS65_LH_CNIVX3 U9682 ( .A(n7862), .Z(n7859) );
  HS65_LH_CNIVX3 U9683 ( .A(n7833), .Z(n7832) );
  HS65_LH_CNIVX3 U9684 ( .A(n7827), .Z(n7824) );
  HS65_LH_CNIVX3 U9685 ( .A(n7826), .Z(n7825) );
  HS65_LH_CNIVX3 U9686 ( .A(n7739), .Z(n7738) );
  HS65_LH_CNIVX3 U9687 ( .A(n7740), .Z(n7737) );
  HS65_LH_CNIVX3 U9688 ( .A(n7746), .Z(n7745) );
  HS65_LH_CNIVX3 U9689 ( .A(n7747), .Z(n7744) );
  HS65_LH_CNIVX3 U9690 ( .A(n7917), .Z(n7916) );
  HS65_LH_NOR2AX3 U9691 ( .A(n8587), .B(rst), .Z(\u_DataPath/cw_tomem_i [3])
         );
  HS65_LH_NOR2AX3 U9692 ( .A(n9385), .B(rst), .Z(\u_DataPath/rs_ex_i [0]) );
  HS65_LH_NOR2AX3 U9693 ( .A(n8805), .B(rst), .Z(\u_DataPath/rs_ex_i [1]) );
  HS65_LH_NOR2AX3 U9694 ( .A(n8797), .B(rst), .Z(\u_DataPath/idex_rt_i [0]) );
  HS65_LH_NOR2AX3 U9695 ( .A(n8813), .B(rst), .Z(\u_DataPath/idex_rt_i [1]) );
  HS65_LH_NOR2X6 U9696 ( .A(n9167), .B(rst), .Z(n8515) );
  HS65_LH_NOR2AX3 U9697 ( .A(n8802), .B(rst), .Z(n8467) );
  HS65_LH_NOR2AX3 U9698 ( .A(iram_data[27]), .B(n7702), .Z(opcode_i[1]) );
  HS65_LH_NOR2AX3 U9699 ( .A(iram_data[2]), .B(n7703), .Z(
        \u_DataPath/immediate_ext_dec_i [2]) );
  HS65_LH_NOR2AX3 U9700 ( .A(iram_data[11]), .B(n7703), .Z(
        \u_DataPath/immediate_ext_dec_i [11]) );
  HS65_LH_NOR2AX3 U9701 ( .A(iram_data[6]), .B(n7703), .Z(
        \u_DataPath/immediate_ext_dec_i [6]) );
  HS65_LH_NOR2AX3 U9702 ( .A(iram_data[21]), .B(n7702), .Z(
        \u_DataPath/u_ifidreg/N57 ) );
  HS65_LH_NOR2AX3 U9703 ( .A(iram_data[17]), .B(n7702), .Z(
        \u_DataPath/jaddr_i [17]) );
  HS65_LH_NOR2AX3 U9704 ( .A(iram_data[18]), .B(n7702), .Z(
        \u_DataPath/jaddr_i [18]) );
  HS65_LH_NOR2AX3 U9705 ( .A(iram_data[20]), .B(n7702), .Z(
        \u_DataPath/jaddr_i [20]) );
  HS65_LH_NOR2AX3 U9706 ( .A(iram_data[24]), .B(n7702), .Z(
        \u_DataPath/jaddr_i [24]) );
  HS65_LH_NOR2AX3 U9707 ( .A(iram_data[13]), .B(n7703), .Z(
        \u_DataPath/immediate_ext_dec_i [13]) );
  HS65_LH_NOR2AX3 U9708 ( .A(iram_data[23]), .B(n7702), .Z(
        \u_DataPath/u_ifidreg/N59 ) );
  HS65_LH_NOR2AX3 U9709 ( .A(iram_data[14]), .B(n7703), .Z(
        \u_DataPath/immediate_ext_dec_i [14]) );
  HS65_LH_NOR2AX3 U9710 ( .A(iram_data[29]), .B(n7702), .Z(opcode_i[3]) );
  HS65_LH_NOR2AX3 U9711 ( .A(iram_data[5]), .B(n7703), .Z(
        \u_DataPath/immediate_ext_dec_i [5]) );
  HS65_LH_NOR2AX3 U9712 ( .A(iram_data[22]), .B(n7702), .Z(
        \u_DataPath/jaddr_i [22]) );
  HS65_LH_NOR2AX3 U9713 ( .A(iram_data[25]), .B(n7702), .Z(
        \u_DataPath/u_ifidreg/N61 ) );
  HS65_LH_NOR2AX3 U9714 ( .A(iram_data[15]), .B(n7703), .Z(
        \u_DataPath/immediate_ext_dec_i [15]) );
  HS65_LH_NOR2AX3 U9715 ( .A(iram_data[12]), .B(n7703), .Z(
        \u_DataPath/immediate_ext_dec_i [12]) );
  HS65_LH_NOR2AX3 U9716 ( .A(iram_data[4]), .B(n7703), .Z(
        \u_DataPath/immediate_ext_dec_i [4]) );
  HS65_LH_NOR2AX3 U9717 ( .A(iram_data[19]), .B(n7702), .Z(
        \u_DataPath/jaddr_i [19]) );
  HS65_LH_NOR2AX3 U9718 ( .A(iram_data[3]), .B(n7703), .Z(
        \u_DataPath/immediate_ext_dec_i [3]) );
  HS65_LH_NOR2AX3 U9719 ( .A(iram_data[0]), .B(n7703), .Z(
        \u_DataPath/immediate_ext_dec_i [0]) );
  HS65_LH_NOR2AX3 U9720 ( .A(iram_data[1]), .B(n7703), .Z(
        \u_DataPath/immediate_ext_dec_i [1]) );
  HS65_LH_NOR2AX3 U9721 ( .A(iram_data[16]), .B(n7702), .Z(
        \u_DataPath/jaddr_i [16]) );
  HS65_LH_NAND2X14 U9722 ( .A(n1885), .B(n8037), .Z(n8071) );
  HS65_LH_NAND2AX4 U9723 ( .A(n7714), .B(n9327), .Z(n8079) );
  HS65_LH_NAND2AX4 U9724 ( .A(n7714), .B(n8843), .Z(n8080) );
  HS65_LH_NAND2AX4 U9725 ( .A(n7714), .B(n9447), .Z(n8082) );
  HS65_LH_NAND2AX4 U9726 ( .A(n7713), .B(n8783), .Z(n8092) );
  HS65_LH_NAND2AX4 U9727 ( .A(n7714), .B(n8782), .Z(n8083) );
  HS65_LH_NAND2AX4 U9728 ( .A(n7713), .B(n9454), .Z(n8085) );
  HS65_LH_NAND2AX4 U9729 ( .A(n7713), .B(n8826), .Z(n8086) );
  HS65_LH_NAND2AX4 U9730 ( .A(n7713), .B(n9372), .Z(n8088) );
  HS65_LH_NAND2AX4 U9731 ( .A(n7713), .B(n8784), .Z(n8089) );
  HS65_LH_NAND2AX4 U9732 ( .A(n7713), .B(n9371), .Z(n8091) );
  HS65_LH_NAND2AX4 U9733 ( .A(n7713), .B(n9370), .Z(n8094) );
  HS65_LH_NAND2AX4 U9734 ( .A(n7713), .B(n9369), .Z(n8096) );
  HS65_LH_NAND2AX4 U9735 ( .A(n7713), .B(n8824), .Z(n8097) );
  HS65_LH_NAND2AX4 U9736 ( .A(n7713), .B(n9405), .Z(n8099) );
  HS65_LH_NAND2AX4 U9737 ( .A(n7713), .B(n8835), .Z(n8100) );
  HS65_LH_NAND2AX4 U9738 ( .A(n7713), .B(n9451), .Z(n8102) );
  HS65_LH_NAND2AX4 U9739 ( .A(n7713), .B(n9279), .Z(n8104) );
  HS65_LH_NAND2AX4 U9740 ( .A(n7713), .B(n9368), .Z(n8106) );
  HS65_LH_NAND2AX4 U9741 ( .A(n7713), .B(n8827), .Z(n8107) );
  HS65_LH_NAND2AX4 U9742 ( .A(n7713), .B(n8786), .Z(n8108) );
  HS65_LH_NAND2AX4 U9743 ( .A(n7713), .B(n9440), .Z(n8110) );
  HS65_LH_NAND2AX4 U9744 ( .A(n7713), .B(n8785), .Z(n8111) );
  HS65_LH_NAND2AX4 U9745 ( .A(n7713), .B(n9442), .Z(n8113) );
  HS65_LH_NAND2AX4 U9746 ( .A(n7714), .B(n8732), .Z(n8048) );
  HS65_LH_NAND2AX4 U9747 ( .A(n7713), .B(\u_DataPath/cw_exmem_i [10]), .Z(
        n8365) );
  HS65_LH_NAND2AX4 U9748 ( .A(n7714), .B(n9083), .Z(n8034) );
  HS65_LH_NAND2AX4 U9749 ( .A(n7714), .B(n9082), .Z(n8032) );
  HS65_LH_NAND2AX4 U9750 ( .A(n7714), .B(n9141), .Z(n8033) );
  HS65_LH_NOR2AX3 U9751 ( .A(\u_DataPath/dataOut_exe_i [31]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [31]) );
  HS65_LH_NOR2AX3 U9752 ( .A(n8553), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [16]) );
  HS65_LH_NOR2AX3 U9753 ( .A(n8747), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [2]) );
  HS65_LH_NOR2AX3 U9754 ( .A(n9330), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [11]) );
  HS65_LH_NOR2AX3 U9755 ( .A(\u_DataPath/dataOut_exe_i [4]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [4]) );
  HS65_LH_NOR2AX3 U9756 ( .A(\u_DataPath/dataOut_exe_i [3]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [3]) );
  HS65_LH_NOR2AX3 U9757 ( .A(\u_DataPath/dataOut_exe_i [25]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [25]) );
  HS65_LH_NOR2AX3 U9758 ( .A(\u_DataPath/dataOut_exe_i [22]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [22]) );
  HS65_LH_NOR2AX3 U9759 ( .A(\u_DataPath/dataOut_exe_i [18]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [18]) );
  HS65_LH_NOR2AX3 U9760 ( .A(\u_DataPath/dataOut_exe_i [21]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [21]) );
  HS65_LH_NOR2AX3 U9761 ( .A(\u_DataPath/dataOut_exe_i [15]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [15]) );
  HS65_LH_NOR2AX3 U9762 ( .A(\u_DataPath/dataOut_exe_i [20]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [20]) );
  HS65_LH_NOR2AX3 U9763 ( .A(\u_DataPath/dataOut_exe_i [30]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [30]) );
  HS65_LH_NOR2AX3 U9764 ( .A(n9541), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [5]) );
  HS65_LH_NOR2AX3 U9765 ( .A(\u_DataPath/dataOut_exe_i [19]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [19]) );
  HS65_LH_NOR2AX3 U9766 ( .A(n9125), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [24]) );
  HS65_LH_NOR2AX3 U9767 ( .A(\u_DataPath/dataOut_exe_i [28]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [28]) );
  HS65_LH_NOR2AX3 U9768 ( .A(\u_DataPath/dataOut_exe_i [14]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [14]) );
  HS65_LH_NOR2AX3 U9769 ( .A(\u_DataPath/dataOut_exe_i [12]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [12]) );
  HS65_LH_NOR2AX3 U9770 ( .A(\u_DataPath/dataOut_exe_i [27]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [27]) );
  HS65_LH_NOR2AX3 U9771 ( .A(\u_DataPath/dataOut_exe_i [13]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [13]) );
  HS65_LH_NOR2AX3 U9772 ( .A(n8748), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [10]) );
  HS65_LH_NOR2AX3 U9773 ( .A(\u_DataPath/dataOut_exe_i [6]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [6]) );
  HS65_LH_NOR2AX3 U9774 ( .A(\u_DataPath/dataOut_exe_i [17]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [17]) );
  HS65_LH_NOR2AX3 U9775 ( .A(n8734), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [9]) );
  HS65_LH_NOR2AX3 U9776 ( .A(\u_DataPath/dataOut_exe_i [23]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [23]) );
  HS65_LH_NOR2AX3 U9777 ( .A(\u_DataPath/dataOut_exe_i [29]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [29]) );
  HS65_LH_NOR2AX3 U9778 ( .A(\u_DataPath/dataOut_exe_i [26]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [26]) );
  HS65_LH_NOR2AX3 U9779 ( .A(n8764), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [8]) );
  HS65_LH_AO22X4 U9780 ( .A(n8461), .B(n9144), .C(n8463), .D(n8454), .Z(
        \u_DataPath/u_execute/psw_status_i [0]) );
  HS65_LH_NOR2AX3 U9781 ( .A(iram_data[9]), .B(n7704), .Z(
        \u_DataPath/immediate_ext_dec_i [9]) );
  HS65_LH_NOR2AX3 U9782 ( .A(iram_data[10]), .B(n7704), .Z(
        \u_DataPath/immediate_ext_dec_i [10]) );
  HS65_LH_NOR2AX3 U9783 ( .A(iram_data[7]), .B(n7704), .Z(
        \u_DataPath/immediate_ext_dec_i [7]) );
  HS65_LH_NOR2AX3 U9784 ( .A(iram_data[8]), .B(n7704), .Z(
        \u_DataPath/immediate_ext_dec_i [8]) );
  HS65_LH_NOR2AX3 U9785 ( .A(iram_data[31]), .B(n7704), .Z(opcode_i[5]) );
  HS65_LH_NOR3AX2 U9786 ( .A(n8443), .B(rst), .C(n8442), .Z(
        \u_DataPath/mem_writedata_out_i [23]) );
  HS65_LH_AO222X4 U9787 ( .A(n7707), .B(n9387), .C(n7689), .D(n8591), .E(n8832), .F(n7687), .Z(addr_to_iram_0) );
  HS65_LH_AO222X4 U9788 ( .A(n7707), .B(n8547), .C(n7689), .D(n8589), .E(n9395), .F(n7687), .Z(\u_DataPath/pc_4_i [0]) );
  HS65_LH_AO222X4 U9789 ( .A(n7707), .B(n8546), .C(n7689), .D(n8590), .E(n8834), .F(n7687), .Z(\u_DataPath/pc_4_i [1]) );
  HS65_LH_AND2X4 U9790 ( .A(n1885), .B(n9140), .Z(
        \u_DataPath/pc4_to_idexreg_i [5]) );
  HS65_LH_AO222X4 U9791 ( .A(n7707), .B(n8936), .C(n7689), .D(n8604), .E(n9404), .F(n7686), .Z(addr_to_iram_2) );
  HS65_LH_AND2X4 U9792 ( .A(n8441), .B(n8459), .Z(
        \u_DataPath/u_decode_unit/hdu_0/current_state [0]) );
  HS65_LH_BFX4 U9793 ( .A(n8181), .Z(n7683) );
  HS65_LH_AO222X4 U9794 ( .A(n7707), .B(n9140), .C(n7689), .D(
        \u_DataPath/jump_address_i [5]), .E(n8831), .F(n7686), .Z(
        addr_to_iram_3) );
  HS65_LH_AO222X4 U9795 ( .A(n7707), .B(n9099), .C(n7689), .D(
        \u_DataPath/jump_address_i [6]), .E(n8829), .F(n7686), .Z(
        addr_to_iram_4) );
  HS65_LH_AND2X4 U9796 ( .A(n1885), .B(n8957), .Z(
        \u_DataPath/pc4_to_idexreg_i [11]) );
  HS65_LH_AND2X4 U9797 ( .A(n1885), .B(n8956), .Z(
        \u_DataPath/pc4_to_idexreg_i [9]) );
  HS65_LH_OAI222X2 U9798 ( .A(n8224), .B(n8223), .C(n8222), .D(n8221), .E(
        n8302), .F(n8220), .Z(\u_DataPath/from_mem_data_out_i [7]) );
  HS65_LH_AO222X4 U9799 ( .A(n7707), .B(n8953), .C(n7689), .D(n8607), .E(n9321), .F(n7686), .Z(addr_to_iram_5) );
  HS65_LH_AO222X4 U9800 ( .A(n7707), .B(n9074), .C(n7689), .D(n8615), .E(n9449), .F(n7686), .Z(addr_to_iram_8) );
  HS65_LH_AO222X4 U9801 ( .A(n7707), .B(n9014), .C(n7689), .D(
        \u_DataPath/jump_address_i [8]), .E(n8828), .F(n7686), .Z(
        addr_to_iram_6) );
  HS65_LH_AO222X4 U9802 ( .A(n7707), .B(n9015), .C(n7690), .D(
        \u_DataPath/jump_address_i [12]), .E(n8822), .F(n7686), .Z(
        addr_to_iram_10) );
  HS65_LH_AO222X4 U9803 ( .A(n7706), .B(n8955), .C(n7691), .D(n9376), .E(n9325), .F(n7685), .Z(addr_to_iram_23) );
  HS65_LH_AO222X4 U9804 ( .A(n7707), .B(n8957), .C(n7689), .D(n9378), .E(n8823), .F(n7686), .Z(addr_to_iram_9) );
  HS65_LH_AO222X4 U9805 ( .A(n7707), .B(n8956), .C(n7689), .D(n8611), .E(n9322), .F(n7686), .Z(addr_to_iram_7) );
  HS65_LH_AO222X4 U9806 ( .A(n7706), .B(n9078), .C(n7690), .D(
        \u_DataPath/jump_address_i [18]), .E(n8838), .F(n7685), .Z(
        addr_to_iram_16) );
  HS65_LH_AO222X4 U9807 ( .A(n7706), .B(n9145), .C(n7690), .D(n8612), .E(n9324), .F(n7686), .Z(addr_to_iram_12) );
  HS65_LH_AO222X4 U9808 ( .A(n7706), .B(n8958), .C(n7690), .D(n9326), .E(n8841), .F(n7686), .Z(addr_to_iram_13) );
  HS65_LH_AO222X4 U9809 ( .A(n7707), .B(n8959), .C(n7690), .D(n9375), .E(n8825), .F(n7686), .Z(addr_to_iram_11) );
  HS65_LH_AND2X4 U9810 ( .A(n1885), .B(n8883), .Z(
        \u_DataPath/pc4_to_idexreg_i [23]) );
  HS65_LH_AND2X4 U9811 ( .A(n1885), .B(n8965), .Z(
        \u_DataPath/pc4_to_idexreg_i [21]) );
  HS65_LH_AO222X4 U9812 ( .A(n7706), .B(n9016), .C(n7691), .D(n8609), .E(n8842), .F(n7685), .Z(addr_to_iram_22) );
  HS65_LH_AO222X4 U9813 ( .A(n7706), .B(n8960), .C(n7690), .D(n8608), .E(n8839), .F(n7685), .Z(addr_to_iram_17) );
  HS65_LH_AND2X4 U9814 ( .A(n1885), .B(n8964), .Z(
        \u_DataPath/pc4_to_idexreg_i [27]) );
  HS65_LH_AND2X4 U9816 ( .A(n9348), .B(n7695), .Z(n8266) );
  HS65_LH_BFX213 U9817 ( .A(n8364), .Z(n7710) );
  HS65_LH_BFX213 U9818 ( .A(n8364), .Z(n7711) );
  HS65_LH_BFX213 U9819 ( .A(n8364), .Z(n7712) );
  HS65_LH_BFX213 U9820 ( .A(n8364), .Z(n7713) );
  HS65_LH_BFX213 U9821 ( .A(n8364), .Z(n7714) );
  HS65_LH_BFX213 U9822 ( .A(n8364), .Z(n7715) );
  HS65_LH_CNIVX27 U9823 ( .A(rst), .Z(n8441) );
  HS65_LH_CNIVX27 U9824 ( .A(n1885), .Z(n8364) );
  HS65_LL_DFPQX4 clk_r_REG515_S1 ( .D(n2785), .CP(clk), .Q(n9463) );
  HS65_LL_DFPQX4 clk_r_REG531_S2 ( .D(n5836), .CP(clk), .Q(n9461) );
  HS65_LL_DFPQX4 clk_r_REG207_S2 ( .D(n5757), .CP(clk), .Q(n9460) );
  HS65_LL_DFPQX4 clk_r_REG137_S2 ( .D(n3034), .CP(clk), .Q(n9459) );
  HS65_LL_DFPQX4 clk_r_REG593_S2 ( .D(n7636), .CP(clk), .Q(n9458) );
  HS65_LL_DFPQX4 clk_r_REG639_S6 ( .D(n3444), .CP(clk), .Q(n9456) );
  HS65_LL_DFPQX4 clk_r_REG213_S3 ( .D(\u_DataPath/jump_address_i [29]), .CP(
        clk), .Q(n9453) );
  HS65_LL_DFPQX4 clk_r_REG182_S1 ( .D(\u_DataPath/branch_target_i [27]), .CP(
        clk), .Q(n9450) );
  HS65_LL_DFPQX4 clk_r_REG32_S2 ( .D(\u_DataPath/dataOut_exe_i [7]), .CP(clk), 
        .Q(n9448) );
  HS65_LL_DFPQX4 clk_r_REG682_S1 ( .D(\u_DataPath/cw_to_ex_i [15]), .CP(clk), 
        .Q(n9445) );
  HS65_LL_DFPQX4 clk_r_REG713_S1 ( .D(\u_DataPath/cw_exmem_i [0]), .CP(clk), 
        .Q(n9443) );
  HS65_LL_DFPQX4 clk_r_REG633_S6 ( .D(n8458), .CP(clk), .Q(n9438) );
  HS65_LL_DFPQX4 clk_r_REG47_S2 ( .D(n5828), .CP(clk), .Q(n9437) );
  HS65_LL_DFPQX4 clk_r_REG928_S6 ( .D(n9427), .CP(clk), .Q(n9426) );
  HS65_LL_DFPQX4 clk_r_REG642_S7 ( .D(n3148), .CP(clk), .Q(n9425) );
  HS65_LL_DFPQX4 clk_r_REG533_S2 ( .D(n5680), .CP(clk), .Q(n9424) );
  HS65_LL_DFPQX4 clk_r_REG543_S2 ( .D(n5597), .CP(clk), .Q(n9423) );
  HS65_LL_DFPQX4 clk_r_REG361_S2 ( .D(n5604), .CP(clk), .Q(n9417) );
  HS65_LL_DFPQX4 clk_r_REG336_S2 ( .D(n7424), .CP(clk), .Q(n9416) );
  HS65_LL_DFPQX4 clk_r_REG644_S7 ( .D(n3235), .CP(clk), .Q(n9415) );
  HS65_LL_DFPQX4 clk_r_REG470_S2 ( .D(n5906), .CP(clk), .Q(n9413) );
  HS65_LL_DFPQX4 clk_r_REG560_S3 ( .D(n2958), .CP(clk), .Q(n9412) );
  HS65_LL_DFPQX4 clk_r_REG222_S2 ( .D(n7308), .CP(clk), .Q(n9411) );
  HS65_LL_DFPQX4 clk_r_REG517_S3 ( .D(n3016), .CP(clk), .Q(n9409) );
  HS65_LL_DFPQX4 clk_r_REG536_S2 ( .D(n7642), .CP(clk), .Q(n9408) );
  HS65_LL_DFPQX4 clk_r_REG400_S3 ( .D(n3129), .CP(clk), .Q(n9407) );
  HS65_LL_DFPQX4 clk_r_REG110_S3 ( .D(\u_DataPath/jump_address_i [31]), .CP(
        clk), .Q(n9406) );
  HS65_LL_DFPQX4 clk_r_REG466_S1 ( .D(\u_DataPath/branch_target_i [4]), .CP(
        clk), .Q(n9404) );
  HS65_LL_DFPQX4 clk_r_REG294_S2 ( .D(n7639), .CP(clk), .Q(n9403) );
  HS65_LL_DFPQX4 clk_r_REG5_S2 ( .D(n2931), .CP(clk), .Q(n9402) );
  HS65_LL_DFPQX4 clk_r_REG397_S1 ( .D(n3029), .CP(clk), .Q(n9401) );
  HS65_LL_DFPQX4 clk_r_REG99_S1 ( .D(n3007), .CP(clk), .Q(n9398) );
  HS65_LL_DFPQX4 clk_r_REG290_S2 ( .D(n5635), .CP(clk), .Q(n9397) );
  HS65_LL_DFPQX4 clk_r_REG354_S2 ( .D(n5577), .CP(clk), .Q(n9394) );
  HS65_LL_DFPQX4 clk_r_REG351_S2 ( .D(n5576), .CP(clk), .Q(n9393) );
  HS65_LL_DFPQX4 clk_r_REG377_S2 ( .D(n5596), .CP(clk), .Q(n9392) );
  HS65_LL_DFPQX4 clk_r_REG345_S2 ( .D(n5870), .CP(clk), .Q(n9391) );
  HS65_LL_DFPQX4 clk_r_REG532_S2 ( .D(n5882), .CP(clk), .Q(n9388) );
  HS65_LL_DFPQX4 clk_r_REG480_S4 ( .D(\u_DataPath/pc_4_i [2]), .CP(net3007), 
        .Q(n9387) );
  HS65_LL_DFPQX4 clk_r_REG358_S2 ( .D(n5606), .CP(clk), .Q(n9386) );
  HS65_LL_DFPQX4 clk_r_REG295_S2 ( .D(n7426), .CP(clk), .Q(n9383) );
  HS65_LL_DFPQX4 clk_r_REG299_S2 ( .D(n3027), .CP(clk), .Q(n9382) );
  HS65_LL_DFPQX4 clk_r_REG489_S2 ( .D(\u_DataPath/u_execute/link_value_i [2]), 
        .CP(clk), .Q(n9381) );
  HS65_LL_DFPQX4 clk_r_REG349_S2 ( .D(n7438), .CP(clk), .Q(n9380) );
  HS65_LL_DFPQX4 clk_r_REG165_S3 ( .D(\u_DataPath/jump_address_i [21]), .CP(
        clk), .Q(n9379) );
  HS65_LL_DFPQX4 clk_r_REG368_S3 ( .D(\u_DataPath/jump_address_i [11]), .CP(
        clk), .Q(n9378) );
  HS65_LL_DFPQX4 clk_r_REG234_S4 ( .D(\u_DataPath/jump_address_i [25]), .CP(
        clk), .Q(n9376) );
  HS65_LL_DFPQX4 clk_r_REG40_S3 ( .D(\u_DataPath/jump_address_i [13]), .CP(clk), .Q(n9375) );
  HS65_LL_DFPQX4 clk_r_REG630_S5 ( .D(n8024), .CP(clk), .Q(n9374) );
  HS65_LL_DFPQX4 clk_r_REG652_S1 ( .D(n8025), .CP(clk), .Q(n9373) );
  HS65_LL_DFPQX4 clk_r_REG693_S1 ( .D(n8363), .CP(clk), .Q(n9367) );
  HS65_LL_DFPQX4 clk_r_REG610_S1 ( .D(n2904), .CP(clk), .Q(n9366) );
  HS65_LL_DFPQX4 clk_r_REG608_S1 ( .D(n2960), .CP(clk), .Q(n9362) );
  HS65_LL_DFPQX4 clk_r_REG325_S2 ( .D(n5779), .CP(clk), .Q(n9347) );
  HS65_LL_DFPQX4 clk_r_REG363_S2 ( .D(n5814), .CP(clk), .Q(n9342) );
  HS65_LL_DFPQX4 clk_r_REG541_S2 ( .D(n5684), .CP(clk), .Q(n9341) );
  HS65_LL_DFPQX4 clk_r_REG413_S3 ( .D(n3096), .CP(clk), .Q(n9340) );
  HS65_LL_DFPQX4 clk_r_REG884_S1 ( .D(n2893), .CP(clk), .Q(n9339) );
  HS65_LL_DFPQX4 clk_r_REG617_S5 ( .D(n3981), .CP(clk), .Q(n9338) );
  HS65_LL_DFPQX4 clk_r_REG393_S2 ( .D(n7436), .CP(clk), .Q(n9337) );
  HS65_LL_DFPQX4 clk_r_REG362_S2 ( .D(n7630), .CP(clk), .Q(n9333) );
  HS65_LL_DFPQX4 clk_r_REG512_S3 ( .D(n8409), .CP(clk), .Q(n9332) );
  HS65_LL_DFPQX4 clk_r_REG410_S3 ( .D(n3145), .CP(clk), .Q(n9331) );
  HS65_LL_DFPQX4 clk_r_REG96_S2 ( .D(\u_DataPath/dataOut_exe_i [11]), .CP(clk), 
        .Q(n9330) );
  HS65_LL_DFPQX4 clk_r_REG128_S5 ( .D(n8196), .CP(clk), .Q(n9329) );
  HS65_LL_DFPQX4 clk_r_REG226_S3 ( .D(\u_DataPath/jump_address_i [27]), .CP(
        clk), .Q(n9328) );
  HS65_LL_DFPQX4 clk_r_REG14_S1 ( .D(\u_DataPath/branch_target_i [25]), .CP(
        clk), .Q(n9325) );
  HS65_LL_DFPQX4 clk_r_REG347_S1 ( .D(\u_DataPath/branch_target_i [14]), .CP(
        clk), .Q(n9324) );
  HS65_LL_DFPQX4 clk_r_REG243_S1 ( .D(\u_DataPath/branch_target_i [23]), .CP(
        clk), .Q(n9323) );
  HS65_LL_DFPQX4 clk_r_REG307_S1 ( .D(\u_DataPath/branch_target_i [9]), .CP(
        clk), .Q(n9322) );
  HS65_LL_DFPQX4 clk_r_REG433_S1 ( .D(\u_DataPath/branch_target_i [7]), .CP(
        clk), .Q(n9321) );
  HS65_LL_DFPQX4 clk_r_REG159_S1 ( .D(\u_DataPath/branch_target_i [21]), .CP(
        clk), .Q(n9320) );
  HS65_LL_DFPQX4 clk_r_REG332_S1 ( .D(\u_DataPath/branch_target_i [16]), .CP(
        clk), .Q(n9319) );
  HS65_LL_DFPQX4 clk_r_REG382_S2 ( .D(n5804), .CP(clk), .Q(n9312) );
  HS65_LL_DFPQX4 clk_r_REG227_S2 ( .D(n5554), .CP(clk), .Q(n9309) );
  HS65_LL_DFPQX4 clk_r_REG589_S2 ( .D(n5553), .CP(clk), .Q(n9308) );
  HS65_LL_DFPQX4 clk_r_REG258_S2 ( .D(n5750), .CP(clk), .Q(n9307) );
  HS65_LL_DFPQX4 clk_r_REG525_S2 ( .D(n5753), .CP(clk), .Q(n9306) );
  HS65_LL_DFPQX4 clk_r_REG245_S2 ( .D(n5552), .CP(clk), .Q(n9305) );
  HS65_LL_DFPQX4 clk_r_REG215_S2 ( .D(n5555), .CP(clk), .Q(n9304) );
  HS65_LL_DFPQX4 clk_r_REG220_S2 ( .D(n5756), .CP(clk), .Q(n9301) );
  HS65_LL_DFPQX4 clk_r_REG262_S2 ( .D(n5548), .CP(clk), .Q(n9300) );
  HS65_LL_DFPQX4 clk_r_REG587_S2 ( .D(n5755), .CP(clk), .Q(n9299) );
  HS65_LL_DFPQX4 clk_r_REG255_S2 ( .D(n5551), .CP(clk), .Q(n9298) );
  HS65_LL_DFPQX4 clk_r_REG233_S2 ( .D(n5754), .CP(clk), .Q(n9297) );
  HS65_LL_DFPQX4 clk_r_REG291_S2 ( .D(n5547), .CP(clk), .Q(n9296) );
  HS65_LL_DFPQX4 clk_r_REG399_S3 ( .D(n3026), .CP(clk), .Q(n9291) );
  HS65_LL_DFPQX4 clk_r_REG263_S2 ( .D(n7442), .CP(clk), .Q(n9290) );
  HS65_LL_DFPQX4 clk_r_REG74_S1 ( .D(n2942), .CP(clk), .Q(n9289) );
  HS65_LL_DFPQX4 clk_r_REG580_S3 ( .D(n3112), .CP(clk), .Q(n9288) );
  HS65_LL_DFPQX4 clk_r_REG100_S3 ( .D(n3010), .CP(clk), .Q(n9287) );
  HS65_LL_DFPQX4 clk_r_REG645_S5 ( .D(n8035), .CP(clk), .Q(n9285) );
  HS65_LL_DFPQX4 clk_r_REG472_S1 ( .D(n2986), .CP(clk), .Q(n9284) );
  HS65_LL_DFPQX4 clk_r_REG78_S3 ( .D(n3066), .CP(clk), .Q(n9283) );
  HS65_LL_DFPQX4 clk_r_REG116_S1 ( .D(\u_DataPath/branch_target_i [31]), .CP(
        clk), .Q(n9281) );
  HS65_LL_DFPQX4 clk_r_REG196_S1 ( .D(\u_DataPath/branch_target_i [29]), .CP(
        clk), .Q(n9280) );
  HS65_LL_DFPQX4 clk_r_REG355_S2 ( .D(n5780), .CP(clk), .Q(n9277) );
  HS65_LL_DFPQX4 clk_r_REG344_S2 ( .D(n5781), .CP(clk), .Q(n9276) );
  HS65_LL_DFPQX4 clk_r_REG538_S2 ( .D(n5805), .CP(clk), .Q(n9275) );
  HS65_LL_DFPQX4 clk_r_REG450_S2 ( .D(n5855), .CP(clk), .Q(n9273) );
  HS65_LL_DFPQX4 clk_r_REG348_S2 ( .D(n5578), .CP(clk), .Q(n9272) );
  HS65_LL_DFPQX4 clk_r_REG357_S2 ( .D(n5812), .CP(clk), .Q(n9271) );
  HS65_LL_DFPQX4 clk_r_REG712_S1 ( .D(n8358), .CP(clk), .Q(n9269) );
  HS65_LL_DFPQX4 clk_r_REG33_S2 ( .D(n8455), .CP(clk), .Q(n9268) );
  HS65_LL_DFPQX4 clk_r_REG677_S6 ( .D(n7694), .CP(clk), .Q(n9252) );
  HS65_LL_DFPQX4 clk_r_REG635_S6 ( .D(n3553), .CP(clk), .Q(n9241) );
  HS65_LL_DFPQX4 clk_r_REG310_S2 ( .D(n5595), .CP(clk), .Q(n9239) );
  HS65_LL_DFPQX4 clk_r_REG553_S2 ( .D(n5711), .CP(clk), .Q(n9238) );
  HS65_LL_DFPQX4 clk_r_REG540_S2 ( .D(n5886), .CP(clk), .Q(n9235) );
  HS65_LL_DFPQX4 clk_r_REG53_S2 ( .D(n7306), .CP(clk), .Q(n9234) );
  HS65_LL_DFPQX4 clk_r_REG285_S2 ( .D(n7640), .CP(clk), .Q(n9232) );
  HS65_LL_DFPQX4 clk_r_REG330_S2 ( .D(n7430), .CP(clk), .Q(n9231) );
  HS65_LL_DFPQX4 clk_r_REG492_S1 ( .D(n8378), .CP(clk), .Q(n9229) );
  HS65_LL_DFPQX4 clk_r_REG707_S1 ( .D(n7941), .CP(clk), .Q(n9228) );
  HS65_LL_DFPQX4 clk_r_REG268_S2 ( .D(n7444), .CP(clk), .Q(n9224) );
  HS65_LL_DFPQX4 clk_r_REG171_S2 ( .D(n6759), .CP(clk), .Q(n9223) );
  HS65_LL_DFPQX4 clk_r_REG574_S5 ( .D(n2956), .CP(clk), .Q(n9222) );
  HS65_LL_DFPQX4 clk_r_REG698_S1 ( .D(n8026), .CP(clk), .Q(n9220) );
  HS65_LL_DFPQX4 clk_r_REG705_S1 ( .D(n7937), .CP(clk), .Q(n9219) );
  HS65_LL_DFPQX4 clk_r_REG701_S1 ( .D(n7940), .CP(clk), .Q(n9218) );
  HS65_LL_DFPQX4 clk_r_REG366_S2 ( .D(n7626), .CP(clk), .Q(n9217) );
  HS65_LL_DFPQX4 clk_r_REG539_S2 ( .D(n7427), .CP(clk), .Q(n9216) );
  HS65_LL_DFPQX4 clk_r_REG431_S2 ( .D(n7419), .CP(clk), .Q(n9214) );
  HS65_LL_DFPQX4 clk_r_REG320_S2 ( .D(n7434), .CP(clk), .Q(n9213) );
  HS65_LL_DFPQX4 clk_r_REG305_S2 ( .D(n7623), .CP(clk), .Q(n9212) );
  HS65_LL_DFPQX4 clk_r_REG674_S7 ( .D(n3527), .CP(clk), .Q(n9210) );
  HS65_LL_DFPQX4 clk_r_REG667_S7 ( .D(n7012), .CP(clk), .Q(n9209) );
  HS65_LL_DFPQX4 clk_r_REG383_S2 ( .D(n7624), .CP(clk), .Q(n9181) );
  HS65_LL_DFPQX4 clk_r_REG373_S2 ( .D(n7432), .CP(clk), .Q(n9180) );
  HS65_LL_DFPQX4 clk_r_REG650_S1 ( .D(n8023), .CP(clk), .Q(n9174) );
  HS65_LL_DFPQX4 clk_r_REG714_S1 ( .D(n2803), .CP(clk), .Q(n9171) );
  HS65_LL_DFPQX4 clk_r_REG603_S6 ( .D(n2912), .CP(clk), .Q(n9151) );
  HS65_LL_DFPQX4 clk_r_REG297_S2 ( .D(n5795), .CP(clk), .Q(n9150) );
  HS65_LL_DFPQX4 clk_r_REG588_S2 ( .D(n5562), .CP(clk), .Q(n9149) );
  HS65_LL_DFPQX4 clk_r_REG436_S2 ( .D(n7621), .CP(clk), .Q(n9148) );
  HS65_LL_DFPQX4 clk_r_REG449_S2 ( .D(n5698), .CP(clk), .Q(n9147) );
  HS65_LL_DFPQX4 clk_r_REG7_S3 ( .D(n8131), .CP(clk), .Q(n9146) );
  HS65_LL_DFPQX4 clk_r_REG341_S5 ( .D(\u_DataPath/pc_4_i [14]), .CP(net3007), 
        .Q(n9145) );
  HS65_LL_DFPQX4 clk_r_REG637_S1 ( .D(n8267), .CP(clk), .Q(n9144) );
  HS65_LL_DFPQX4 clk_r_REG716_S1 ( .D(\u_DataPath/cw_exmem_i [6]), .CP(clk), 
        .Q(n9141) );
  HS65_LL_DFPQX4 clk_r_REG453_S4 ( .D(\u_DataPath/pc_4_i [5]), .CP(net3007), 
        .Q(n9140) );
  HS65_LL_DFPQX4 clk_r_REG340_S2 ( .D(n5747), .CP(clk), .Q(n9139) );
  HS65_LL_DFPQX4 clk_r_REG467_S2 ( .D(\u_DataPath/u_execute/link_value_i [4]), 
        .CP(clk), .Q(n9138) );
  HS65_LL_DFPQX4 clk_r_REG202_S2 ( .D(n5556), .CP(clk), .Q(n9136) );
  HS65_LL_DFPQX4 clk_r_REG205_S2 ( .D(n5869), .CP(clk), .Q(n9133) );
  HS65_LL_DFPQX4 clk_r_REG209_S2 ( .D(n5866), .CP(clk), .Q(n9132) );
  HS65_LL_DFPQX4 clk_r_REG251_S2 ( .D(n5839), .CP(clk), .Q(n9131) );
  HS65_LL_DFPQX4 clk_r_REG394_S2 ( .D(n5691), .CP(clk), .Q(n9130) );
  HS65_LL_DFPQX4 clk_r_REG448_S2 ( .D(n5903), .CP(clk), .Q(n9129) );
  HS65_LL_DFPQX4 clk_r_REG592_S2 ( .D(n5784), .CP(clk), .Q(n9128) );
  HS65_LL_DFPQX4 clk_r_REG237_S2 ( .D(n5581), .CP(clk), .Q(n9127) );
  HS65_LL_DFPQX4 clk_r_REG127_S4 ( .D(\u_DataPath/dataOut_exe_i [24]), .CP(clk), .Q(n9125) );
  HS65_LL_DFPQX4 clk_r_REG582_S1 ( .D(\u_DataPath/mem_writedata_out_i [26]), 
        .CP(clk), .Q(n9122) );
  HS65_LL_DFPQX4 clk_r_REG497_S1 ( .D(\u_DataPath/mem_writedata_out_i [30]), 
        .CP(clk), .Q(n9120) );
  HS65_LL_DFPQX4 clk_r_REG578_S1 ( .D(\u_DataPath/mem_writedata_out_i [28]), 
        .CP(clk), .Q(n9119) );
  HS65_LL_DFPQX4 clk_r_REG632_S6 ( .D(n3566), .CP(clk), .Q(n9115) );
  HS65_LL_DFPQX4 clk_r_REG658_S7 ( .D(n2887), .CP(clk), .Q(n9114) );
  HS65_LL_DFPQX4 clk_r_REG460_S2 ( .D(n5648), .CP(clk), .Q(n9109) );
  HS65_LL_DFPQX4 clk_r_REG195_S2 ( .D(n5675), .CP(clk), .Q(n9108) );
  HS65_LL_DFPQX4 clk_r_REG292_S2 ( .D(n5877), .CP(clk), .Q(n9107) );
  HS65_LL_DFPQX4 clk_r_REG20_S3 ( .D(\u_DataPath/u_execute/link_value_i [26]), 
        .CP(clk), .Q(n9105) );
  HS65_LL_DFPQX4 clk_r_REG649_S1 ( .D(
        \u_DataPath/u_decode_unit/hdu_0/current_state [1]), .CP(clk), .Q(n9104) );
  HS65_LL_DFPQX4 clk_r_REG660_S7 ( .D(n2988), .CP(clk), .Q(n9103) );
  HS65_LL_DFPQX4 clk_r_REG439_S4 ( .D(\u_DataPath/pc_4_i [6]), .CP(net3007), 
        .Q(n9099) );
  HS65_LL_DFPQX4 clk_r_REG606_S1 ( .D(n2888), .CP(clk), .Q(n9094) );
  HS65_LL_DFPQX4 clk_r_REG432_S2 ( .D(n5702), .CP(clk), .Q(n9088) );
  HS65_LL_DFPQX4 clk_r_REG293_S2 ( .D(n5626), .CP(clk), .Q(n9087) );
  HS65_LL_DFPQX4 clk_r_REG488_S2 ( .D(n5710), .CP(clk), .Q(n9086) );
  HS65_LL_DFPQX4 clk_r_REG485_S2 ( .D(n5712), .CP(clk), .Q(n9085) );
  HS65_LL_DFPQX4 clk_r_REG277_S2 ( .D(n7440), .CP(clk), .Q(n9084) );
  HS65_LL_DFPQX4 clk_r_REG629_S5 ( .D(\u_DataPath/u_idexreg/N15 ), .CP(clk), 
        .Q(n9083) );
  HS65_LL_DFPQX4 clk_r_REG651_S1 ( .D(\u_DataPath/u_idexreg/N16 ), .CP(clk), 
        .Q(n9082) );
  HS65_LL_DFPQX4 clk_r_REG575_S2 ( .D(n8305), .CP(clk), .Q(n9081) );
  HS65_LL_DFPQX4 clk_r_REG681_S1 ( .D(n8513), .CP(clk), .Q(n9080) );
  HS65_LL_DFPQX4 clk_r_REG54_S3 ( .D(\u_DataPath/u_execute/link_value_i [22]), 
        .CP(clk), .Q(n9079) );
  HS65_LL_DFPQX4 clk_r_REG280_S2 ( .D(\u_DataPath/pc_4_i [18]), .CP(net3007), 
        .Q(n9078) );
  HS65_LL_DFPQX4 clk_r_REG468_S3 ( .D(n8304), .CP(clk), .Q(n9077) );
  HS65_LL_DFPQX4 clk_r_REG264_S2 ( .D(n7631), .CP(clk), .Q(n9075) );
  HS65_LL_DFPQX4 clk_r_REG36_S4 ( .D(\u_DataPath/pc_4_i [10]), .CP(net3007), 
        .Q(n9074) );
  HS65_LL_DFPQX4 clk_r_REG605_S1 ( .D(n8041), .CP(clk), .Q(n9066) );
  HS65_LL_DFPQX4 clk_r_REG478_S2 ( .D(n5534), .CP(clk), .Q(n9060) );
  HS65_LL_DFPQX4 clk_r_REG442_S2 ( .D(n5649), .CP(clk), .Q(n9057) );
  HS65_LL_DFPQX4 clk_r_REG375_S2 ( .D(n5574), .CP(clk), .Q(n9056) );
  HS65_LL_DFPQX4 clk_r_REG435_S2 ( .D(n5538), .CP(clk), .Q(n9055) );
  HS65_LL_DFPQX4 clk_r_REG274_S2 ( .D(n5826), .CP(clk), .Q(n9050) );
  HS65_LL_DFPQX4 clk_r_REG376_S2 ( .D(n5777), .CP(clk), .Q(n9049) );
  HS65_LL_DFPQX4 clk_r_REG479_S2 ( .D(n5735), .CP(clk), .Q(n9048) );
  HS65_LL_DFPQX4 clk_r_REG335_S2 ( .D(n5783), .CP(clk), .Q(n9047) );
  HS65_LL_DFPQX4 clk_r_REG648_S6 ( .D(n7215), .CP(clk), .Q(n9043) );
  HS65_LL_DFPQX4 clk_r_REG356_S2 ( .D(n7423), .CP(clk), .Q(n9042) );
  HS65_LL_DFPQX4 clk_r_REG115_S2 ( .D(n5671), .CP(clk), .Q(n9041) );
  HS65_LL_DFPQX4 clk_r_REG164_S2 ( .D(n5822), .CP(clk), .Q(n9039) );
  HS65_LL_DFPQX4 clk_r_REG221_S2 ( .D(n5559), .CP(clk), .Q(n9037) );
  HS65_LL_DFPQX4 clk_r_REG236_S2 ( .D(n5930), .CP(clk), .Q(n9035) );
  HS65_LL_DFPQX4 clk_r_REG208_S2 ( .D(n5667), .CP(clk), .Q(n9034) );
  HS65_LL_DFPQX4 clk_r_REG246_S2 ( .D(n5841), .CP(clk), .Q(n9033) );
  HS65_LL_DFPQX4 clk_r_REG526_S2 ( .D(n5640), .CP(clk), .Q(n9032) );
  HS65_LL_DFPQX4 clk_r_REG590_S2 ( .D(n5786), .CP(clk), .Q(n9031) );
  HS65_LL_DFPQX4 clk_r_REG252_S2 ( .D(n5715), .CP(clk), .Q(n9030) );
  HS65_LL_DFPQX4 clk_r_REG228_S2 ( .D(n5767), .CP(clk), .Q(n9029) );
  HS65_LL_DFPQX4 clk_r_REG214_S2 ( .D(n5762), .CP(clk), .Q(n9028) );
  HS65_LL_DFPQX4 clk_r_REG276_S2 ( .D(n5631), .CP(clk), .Q(n9027) );
  HS65_LL_DFPQX4 clk_r_REG585_S2 ( .D(n5564), .CP(clk), .Q(n9026) );
  HS65_LL_DFPQX4 clk_r_REG172_S2 ( .D(n5583), .CP(clk), .Q(n9025) );
  HS65_LL_DFPQX4 clk_r_REG261_S2 ( .D(n5825), .CP(clk), .Q(n9024) );
  HS65_LL_DFPQX4 clk_r_REG203_S1 ( .D(\u_DataPath/branch_target_i [30]), .CP(
        clk), .Q(n9022) );
  HS65_LL_DFPQX4 clk_r_REG690_S1 ( .D(n7974), .CP(clk), .Q(n9021) );
  HS65_LL_DFPQX4 clk_r_REG43_S4 ( .D(\u_DataPath/pc_4_i [16]), .CP(net3007), 
        .Q(n9019) );
  HS65_LL_DFPQX4 clk_r_REG609_S1 ( .D(n3214), .CP(clk), .Q(n9018) );
  HS65_LL_DFPQX4 clk_r_REG50_S4 ( .D(\u_DataPath/pc_4_i [22]), .CP(net3007), 
        .Q(n9017) );
  HS65_LL_DFPQX4 clk_r_REG168_S4 ( .D(\u_DataPath/pc_4_i [24]), .CP(net3007), 
        .Q(n9016) );
  HS65_LL_DFPQX4 clk_r_REG313_S4 ( .D(\u_DataPath/pc_4_i [12]), .CP(net3007), 
        .Q(n9015) );
  HS65_LL_DFPQX4 clk_r_REG384_S4 ( .D(\u_DataPath/pc_4_i [8]), .CP(net3007), 
        .Q(n9014) );
  HS65_LL_DFPQX4 clk_r_REG447_S2 ( .D(n7418), .CP(clk), .Q(n9013) );
  HS65_LL_DFPQX4 clk_r_REG473_S2 ( .D(n5917), .CP(clk), .Q(n9011) );
  HS65_LL_DFPQX4 clk_r_REG591_S2 ( .D(n5788), .CP(clk), .Q(n9008) );
  HS65_LL_DFPQX4 clk_r_REG380_S2 ( .D(n5897), .CP(clk), .Q(n9007) );
  HS65_LL_DFPQX4 clk_r_REG483_S2 ( .D(n5860), .CP(clk), .Q(n9004) );
  HS65_LL_DFPQX4 clk_r_REG337_S2 ( .D(n5544), .CP(clk), .Q(n9003) );
  HS65_LL_DFPQX4 clk_r_REG225_S2 ( .D(n5769), .CP(clk), .Q(n9002) );
  HS65_LL_DFPQX4 clk_r_REG173_S2 ( .D(n5585), .CP(clk), .Q(n9001) );
  HS65_LL_DFPQX4 clk_r_REG247_S2 ( .D(n5843), .CP(clk), .Q(n8999) );
  HS65_LL_DFPQX4 clk_r_REG339_S2 ( .D(n5745), .CP(clk), .Q(n8998) );
  HS65_LL_DFPQX4 clk_r_REG89_S4 ( .D(\u_DataPath/pc_4_i [3]), .CP(net3007), 
        .Q(n8997) );
  HS65_LL_DFPQX4 clk_r_REG586_S2 ( .D(n5566), .CP(clk), .Q(n8995) );
  HS65_LL_DFPQX4 clk_r_REG13_S2 ( .D(n5730), .CP(clk), .Q(n8993) );
  HS65_LL_DFPQX4 clk_r_REG181_S2 ( .D(n5722), .CP(clk), .Q(n8992) );
  HS65_LL_DFPQX4 clk_r_REG117_S2 ( .D(n5759), .CP(clk), .Q(n8991) );
  HS65_LL_DFPQX4 clk_r_REG456_S2 ( .D(n5849), .CP(clk), .Q(n8988) );
  HS65_LL_DFPQX4 clk_r_REG524_S2 ( .D(n5925), .CP(clk), .Q(n8987) );
  HS65_LL_DFPQX4 clk_r_REG484_S2 ( .D(n5913), .CP(clk), .Q(n8985) );
  HS65_LL_DFPQX4 clk_r_REG211_S2 ( .D(n5760), .CP(clk), .Q(n8984) );
  HS65_LL_DFPQX4 clk_r_REG217_S2 ( .D(n5926), .CP(clk), .Q(n8983) );
  HS65_LL_DFPQX4 clk_r_REG224_S2 ( .D(n5765), .CP(clk), .Q(n8982) );
  HS65_LL_DFPQX4 clk_r_REG583_S2 ( .D(n5918), .CP(clk), .Q(n8981) );
  HS65_LL_DFPQX4 clk_r_REG187_S2 ( .D(n5557), .CP(clk), .Q(n8979) );
  HS65_LL_DFPQX4 clk_r_REG201_S2 ( .D(n5669), .CP(clk), .Q(n8978) );
  HS65_LL_DFPQX4 clk_r_REG392_S2 ( .D(n5893), .CP(clk), .Q(n8977) );
  HS65_LL_DFPQX4 clk_r_REG163_S2 ( .D(n5817), .CP(clk), .Q(n8976) );
  HS65_LL_DFPQX4 clk_r_REG259_S2 ( .D(n5823), .CP(clk), .Q(n8975) );
  HS65_LL_DFPQX4 clk_r_REG444_S2 ( .D(n5901), .CP(clk), .Q(n8974) );
  HS65_LL_DFPQX4 clk_r_REG12_S2 ( .D(n5727), .CP(clk), .Q(n8973) );
  HS65_LL_DFPQX4 clk_r_REG389_S2 ( .D(n5692), .CP(clk), .Q(n8972) );
  HS65_LL_DFPQX4 clk_r_REG23_S2 ( .D(n8340), .CP(clk), .Q(n8970) );
  HS65_LL_DFPQX4 clk_r_REG191_S4 ( .D(\u_DataPath/pc_4_i [29]), .CP(net3007), 
        .Q(n8967) );
  HS65_LL_DFPQX4 clk_r_REG146_S3 ( .D(\u_DataPath/pc_4_i [17]), .CP(net3007), 
        .Q(n8966) );
  HS65_LL_DFPQX4 clk_r_REG161_S2 ( .D(\u_DataPath/pc_4_i [21]), .CP(net3007), 
        .Q(n8965) );
  HS65_LL_DFPQX4 clk_r_REG178_S4 ( .D(\u_DataPath/pc_4_i [27]), .CP(net3007), 
        .Q(n8964) );
  HS65_LL_DFPQX4 clk_r_REG624_S5 ( .D(n8468), .CP(clk), .Q(n8963) );
  HS65_LL_DFPQX4 clk_r_REG16_S4 ( .D(\u_DataPath/pc_4_i [26]), .CP(net3007), 
        .Q(n8961) );
  HS65_LL_DFPQX4 clk_r_REG266_S2 ( .D(\u_DataPath/pc_4_i [19]), .CP(net3007), 
        .Q(n8960) );
  HS65_LL_DFPQX4 clk_r_REG318_S4 ( .D(\u_DataPath/pc_4_i [13]), .CP(net3007), 
        .Q(n8959) );
  HS65_LL_DFPQX4 clk_r_REG328_S5 ( .D(\u_DataPath/pc_4_i [15]), .CP(net3007), 
        .Q(n8958) );
  HS65_LL_DFPQX4 clk_r_REG364_S4 ( .D(\u_DataPath/pc_4_i [11]), .CP(net3007), 
        .Q(n8957) );
  HS65_LL_DFPQX4 clk_r_REG303_S4 ( .D(\u_DataPath/pc_4_i [9]), .CP(net3007), 
        .Q(n8956) );
  HS65_LL_DFPQX4 clk_r_REG429_S4 ( .D(\u_DataPath/pc_4_i [7]), .CP(net3007), 
        .Q(n8953) );
  HS65_LL_DFPQX4 clk_r_REG446_S2 ( .D(\u_DataPath/u_execute/link_value_i [6]), 
        .CP(clk), .Q(n8952) );
  HS65_LL_DFPQX4 clk_r_REG669_S7 ( .D(n2889), .CP(clk), .Q(n8945) );
  HS65_LL_DFPQX4 clk_r_REG475_S2 ( .D(n5714), .CP(clk), .Q(n8944) );
  HS65_LL_DFPQX4 clk_r_REG91_S2 ( .D(\u_DataPath/u_execute/link_value_i [3]), 
        .CP(clk), .Q(n8943) );
  HS65_LL_DFPQX4 clk_r_REG676_S7 ( .D(n2910), .CP(clk), .Q(n8941) );
  HS65_LL_DFPQX4 clk_r_REG421_S4 ( .D(\u_DataPath/pc_4_i [4]), .CP(net3007), 
        .Q(n8936) );
  HS65_LL_DFPQX4 clk_r_REG643_S7 ( .D(n2952), .CP(clk), .Q(n8935) );
  HS65_LL_DFPQX4 clk_r_REG346_S2 ( .D(n5679), .CP(clk), .Q(n8932) );
  HS65_LL_DFPQX4 clk_r_REG188_S2 ( .D(n5561), .CP(clk), .Q(n8931) );
  HS65_LL_DFPQX4 clk_r_REG359_S2 ( .D(n5588), .CP(clk), .Q(n8930) );
  HS65_LL_DFPQX4 clk_r_REG352_S2 ( .D(n5608), .CP(clk), .Q(n8929) );
  HS65_LL_DFPQX4 clk_r_REG370_S2 ( .D(n5599), .CP(clk), .Q(n8928) );
  HS65_LL_DFPQX4 clk_r_REG542_S2 ( .D(n5687), .CP(clk), .Q(n8926) );
  HS65_LL_DFPQX4 clk_r_REG697_S1 ( .D(n2911), .CP(clk), .Q(n8925) );
  HS65_LL_DFPQX4 clk_r_REG306_S2 ( .D(n5694), .CP(clk), .Q(n8924) );
  HS65_LL_DFPQX4 clk_r_REG390_S2 ( .D(n5644), .CP(clk), .Q(n8923) );
  HS65_LL_DFPQX4 clk_r_REG527_S2 ( .D(n5642), .CP(clk), .Q(n8922) );
  HS65_LL_DFPQX4 clk_r_REG457_S2 ( .D(n5656), .CP(clk), .Q(n8921) );
  HS65_LL_DFPQX4 clk_r_REG465_S2 ( .D(n5706), .CP(clk), .Q(n8920) );
  HS65_LL_DFPQX4 clk_r_REG149_S2 ( .D(n5622), .CP(clk), .Q(n8919) );
  HS65_LL_DFPQX4 clk_r_REG534_S2 ( .D(n5683), .CP(clk), .Q(n8918) );
  HS65_LL_DFPQX4 clk_r_REG455_S2 ( .D(n5857), .CP(clk), .Q(n8916) );
  HS65_LL_DFPQX4 clk_r_REG212_S2 ( .D(n5764), .CP(clk), .Q(n8915) );
  HS65_LL_DFPQX4 clk_r_REG321_S2 ( .D(n5816), .CP(clk), .Q(n8914) );
  HS65_LL_DFPQX4 clk_r_REG437_S2 ( .D(n5905), .CP(clk), .Q(n8913) );
  HS65_LL_DFPQX4 clk_r_REG438_S2 ( .D(n5739), .CP(clk), .Q(n8911) );
  HS65_LL_DFPQX4 clk_r_REG537_S2 ( .D(n5889), .CP(clk), .Q(n8910) );
  HS65_LL_DFPQX4 clk_r_REG367_S2 ( .D(n5807), .CP(clk), .Q(n8909) );
  HS65_LL_DFPQX4 clk_r_REG343_S2 ( .D(n5873), .CP(clk), .Q(n8908) );
  HS65_LL_DFPQX4 clk_r_REG445_S2 ( .D(n5850), .CP(clk), .Q(n8907) );
  HS65_LL_DFPQX4 clk_r_REG283_S2 ( .D(n5796), .CP(clk), .Q(n8905) );
  HS65_LL_DFPQX4 clk_r_REG148_S2 ( .D(n5838), .CP(clk), .Q(n8904) );
  HS65_LL_DFPQX4 clk_r_REG260_S2 ( .D(n5831), .CP(clk), .Q(n8903) );
  HS65_LL_DFPQX4 clk_r_REG388_S2 ( .D(n5845), .CP(clk), .Q(n8902) );
  HS65_LL_DFPQX4 clk_r_REG704_S1 ( .D(n2913), .CP(clk), .Q(n8899) );
  HS65_LL_DFPQX4 clk_r_REG253_S2 ( .D(n5718), .CP(clk), .Q(n8896) );
  HS65_LL_DFPQX4 clk_r_REG157_S2 ( .D(n5615), .CP(clk), .Q(n8895) );
  HS65_LL_DFPQX4 clk_r_REG288_S2 ( .D(n5628), .CP(clk), .Q(n8894) );
  HS65_LL_DFPQX4 clk_r_REG180_S2 ( .D(n5719), .CP(clk), .Q(n8892) );
  HS65_LL_DFPQX4 clk_r_REG287_S2 ( .D(n5623), .CP(clk), .Q(n8891) );
  HS65_LL_DFPQX4 clk_r_REG156_S2 ( .D(n5609), .CP(clk), .Q(n8890) );
  HS65_LL_DFPQX4 clk_r_REG241_S2 ( .D(n5723), .CP(clk), .Q(n8889) );
  HS65_LL_DFPQX4 clk_r_REG387_S2 ( .D(n5895), .CP(clk), .Q(n8888) );
  HS65_LL_DFPQX4 clk_r_REG482_S2 ( .D(n5915), .CP(clk), .Q(n8887) );
  HS65_LL_DFPQX4 clk_r_REG282_S2 ( .D(n5879), .CP(clk), .Q(n8886) );
  HS65_LL_DFPQX4 clk_r_REG239_S4 ( .D(\u_DataPath/pc_4_i [23]), .CP(net3007), 
        .Q(n8883) );
  HS65_LL_DFPQX4 clk_r_REG231_S2 ( .D(n5933), .CP(clk), .Q(n8881) );
  HS65_LL_DFPQX4 clk_r_REG584_S2 ( .D(n5921), .CP(clk), .Q(n8880) );
  HS65_LL_DFPQX4 clk_r_REG189_S1 ( .D(\u_DataPath/branch_target_i [28]), .CP(
        clk), .Q(n8877) );
  HS65_LL_DFPQX4 clk_r_REG83_S1 ( .D(n2863), .CP(clk), .Q(n8875) );
  HS65_LL_DFPQX4 clk_r_REG95_S2 ( .D(n8323), .CP(clk), .Q(n8873) );
  HS65_LL_DFPQX4 clk_r_REG550_S2 ( .D(\u_DataPath/toPC2_i [1]), .CP(clk), .Q(
        n8871) );
  HS65_LL_DFPQX4 clk_r_REG569_S2 ( .D(\u_DataPath/u_execute/resAdd1_i [0]), 
        .CP(clk), .Q(n8870) );
  HS65_LL_DFPQX4 clk_r_REG554_S2 ( .D(\u_DataPath/u_execute/resAdd1_i [1]), 
        .CP(clk), .Q(n8869) );
  HS65_LL_DFPQX4 clk_r_REG673_S7 ( .D(n7217), .CP(clk), .Q(n8847) );
  HS65_LL_DFPQX4 clk_r_REG662_S7 ( .D(n8013), .CP(clk), .Q(n8846) );
  HS65_LL_DFPQX4 clk_r_REG238_S3 ( .D(\u_DataPath/u_execute/link_value_i [25]), 
        .CP(clk), .Q(n8844) );
  HS65_LL_DFPQX4 clk_r_REG174_S1 ( .D(\u_DataPath/branch_target_i [24]), .CP(
        clk), .Q(n8842) );
  HS65_LL_DFPQX4 clk_r_REG334_S1 ( .D(\u_DataPath/branch_target_i [15]), .CP(
        clk), .Q(n8841) );
  HS65_LL_DFPQX4 clk_r_REG254_S1 ( .D(\u_DataPath/branch_target_i [22]), .CP(
        clk), .Q(n8840) );
  HS65_LL_DFPQX4 clk_r_REG152_S1 ( .D(\u_DataPath/branch_target_i [19]), .CP(
        clk), .Q(n8839) );
  HS65_LL_DFPQX4 clk_r_REG278_S1 ( .D(\u_DataPath/branch_target_i [18]), .CP(
        clk), .Q(n8838) );
  HS65_LL_DFPQX4 clk_r_REG150_S1 ( .D(\u_DataPath/branch_target_i [17]), .CP(
        clk), .Q(n8837) );
  HS65_LL_DFPQX4 clk_r_REG458_S1 ( .D(\u_DataPath/branch_target_i [5]), .CP(
        clk), .Q(n8831) );
  HS65_LL_DFPQX4 clk_r_REG391_S1 ( .D(\u_DataPath/branch_target_i [8]), .CP(
        clk), .Q(n8828) );
  HS65_LL_DFPQX4 clk_r_REG353_S1 ( .D(\u_DataPath/branch_target_i [13]), .CP(
        clk), .Q(n8825) );
  HS65_LL_DFPQX4 clk_r_REG371_S1 ( .D(\u_DataPath/branch_target_i [11]), .CP(
        clk), .Q(n8823) );
  HS65_LL_DFPQX4 clk_r_REG360_S1 ( .D(\u_DataPath/branch_target_i [12]), .CP(
        clk), .Q(n8822) );
  HS65_LL_DFPQX4 clk_r_REG688_S1 ( .D(n7991), .CP(clk), .Q(n8821) );
  HS65_LL_DFPQX4 clk_r_REG797_S1 ( .D(\u_DataPath/idex_rt_i [0]), .CP(clk), 
        .Q(n8820) );
  HS65_LL_DFPQX4 clk_r_REG647_S6 ( .D(
        \u_DataPath/u_decode_unit/hdu_0/current_state [0]), .CP(clk), .Q(n8787) );
  HS65_LL_DFPQX4 clk_r_REG556_S3 ( .D(n8266), .CP(clk), .Q(n8781) );
  HS65_LL_DFPQX4 clk_r_REG131_S2 ( .D(n8324), .CP(clk), .Q(n8780) );
  HS65_LL_DFPQX4 clk_r_REG140_S3 ( .D(n8332), .CP(clk), .Q(n8779) );
  HS65_LL_DFPQX4 clk_r_REG646_S5 ( .D(n7211), .CP(clk), .Q(n8778) );
  HS65_LL_DFPQX4 clk_r_REG39_S2 ( .D(n5776), .CP(clk), .Q(n8777) );
  HS65_LL_DFPQX4 clk_r_REG426_S2 ( .D(n5738), .CP(clk), .Q(n8776) );
  HS65_LL_DFPQX4 clk_r_REG474_S2 ( .D(n5734), .CP(clk), .Q(n8773) );
  HS65_LL_DFPQX4 clk_r_REG595_S5 ( .D(n7999), .CP(clk), .Q(n8772) );
  HS65_LL_DFPQX4 clk_r_REG4_S2 ( .D(n8066), .CP(clk), .Q(n8771) );
  HS65_LL_DFPQX4 clk_r_REG577_S2 ( .D(n8308), .CP(clk), .Q(n8770) );
  HS65_LL_DFPQX4 clk_r_REG514_S1 ( .D(n8160), .CP(clk), .Q(n8769) );
  HS65_LL_DFPQX4 clk_r_REG3_S1 ( .D(n7666), .CP(clk), .Q(n8768) );
  HS65_LL_DFPQX4 clk_r_REG105_S3 ( .D(n8337), .CP(clk), .Q(n8765) );
  HS65_LL_DFPQX4 clk_r_REG298_S2 ( .D(\u_DataPath/dataOut_exe_i [8]), .CP(clk), 
        .Q(n8764) );
  HS65_LL_DFPQX4 clk_r_REG73_S2 ( .D(n8341), .CP(clk), .Q(n8763) );
  HS65_LL_DFPQX4 clk_r_REG107_S1 ( .D(\u_DataPath/mem_writedata_out_i [31]), 
        .CP(clk), .Q(n8762) );
  HS65_LL_DFPQX4 clk_r_REG521_S4 ( .D(\u_DataPath/mem_writedata_out_i [25]), 
        .CP(clk), .Q(n8761) );
  HS65_LL_DFPQX4 clk_r_REG607_S1 ( .D(n2885), .CP(clk), .Q(n8760) );
  HS65_LL_DFPQX4 clk_r_REG46_S2 ( .D(n5827), .CP(clk), .Q(n8759) );
  HS65_LL_DFPQX4 clk_r_REG654_S5 ( .D(n8155), .CP(clk), .Q(n8758) );
  HS65_LL_DFPQX4 clk_r_REG124_S2 ( .D(n8331), .CP(clk), .Q(n8755) );
  HS65_LL_DFPQX4 clk_r_REG82_S2 ( .D(n8328), .CP(clk), .Q(n8754) );
  HS65_LL_DFPQX4 clk_r_REG132_S4 ( .D(n8355), .CP(clk), .Q(n8753) );
  HS65_LL_DFPQX4 clk_r_REG710_S1 ( .D(\u_DataPath/cw_to_ex_i [17]), .CP(clk), 
        .Q(n8752) );
  HS65_LL_DFPQX4 clk_r_REG24_S1 ( .D(n7653), .CP(clk), .Q(n8751) );
  HS65_LL_DFPQX4 clk_r_REG119_S3 ( .D(n8329), .CP(clk), .Q(n8749) );
  HS65_LL_DFPQX4 clk_r_REG64_S3 ( .D(\u_DataPath/dataOut_exe_i [10]), .CP(clk), 
        .Q(n8748) );
  HS65_LL_DFPQX4 clk_r_REG86_S2 ( .D(\u_DataPath/dataOut_exe_i [2]), .CP(clk), 
        .Q(n8747) );
  HS65_LL_DFPQX4 clk_r_REG102_S4 ( .D(n8335), .CP(clk), .Q(n8746) );
  HS65_LL_DFPQX4 clk_r_REG22_S2 ( .D(n8334), .CP(clk), .Q(n8745) );
  HS65_LL_DFPQX4 clk_r_REG79_S4 ( .D(n8336), .CP(clk), .Q(n8744) );
  HS65_LL_DFPQX4 clk_r_REG622_S5 ( .D(n7952), .CP(clk), .Q(n8743) );
  HS65_LL_DFPQX4 clk_r_REG680_S1 ( .D(n7975), .CP(clk), .Q(n8742) );
  HS65_LL_DFPQX4 clk_r_REG631_S6 ( .D(n8163), .CP(clk), .Q(n8740) );
  HS65_LL_DFPQX4 clk_r_REG552_S2 ( .D(n5658), .CP(clk), .Q(n8736) );
  HS65_LL_DFPQX4 clk_r_REG29_S3 ( .D(n8343), .CP(clk), .Q(n8735) );
  HS65_LL_DFPQX4 clk_r_REG136_S2 ( .D(\u_DataPath/dataOut_exe_i [9]), .CP(clk), 
        .Q(n8734) );
  HS65_LL_DFPQX4 clk_r_REG561_S2 ( .D(\u_DataPath/from_mem_data_out_i [30]), 
        .CP(clk), .Q(n8733) );
  HS65_LL_DFPQX4 clk_r_REG689_S1 ( .D(n7989), .CP(clk), .Q(n8731) );
  HS65_LL_DFPQX4 clk_r_REG616_S5 ( .D(n8526), .CP(clk), .Q(n8730) );
  HS65_LL_DFPQX4 clk_r_REG686_S1 ( .D(n7998), .CP(clk), .Q(n8729) );
  HS65_LL_DFPQX4 clk_r_REG636_S1 ( .D(n3561), .CP(clk), .Q(n8728) );
  HS65_LL_DFPQX4 clk_r_REG1_S1 ( .D(n3562), .CP(clk), .Q(n8727) );
  HS65_LL_DFPQX4 clk_r_REG663_S7 ( .D(n3531), .CP(clk), .Q(n8726) );
  HS65_LL_DFPQX4 clk_r_REG98_S1 ( .D(n8213), .CP(clk), .Q(n8724) );
  HS65_LL_DFPQX4 clk_r_REG477_S2 ( .D(n5533), .CP(clk), .Q(n8722) );
  HS65_LL_DFPQX4 clk_r_REG659_S7 ( .D(n3530), .CP(clk), .Q(n8720) );
  HS65_LL_DFPQX4 clk_r_REG55_S1 ( .D(n8273), .CP(clk), .Q(n8719) );
  HS65_LL_DFPQX4 clk_r_REG129_S1 ( .D(n8144), .CP(clk), .Q(n8717) );
  HS65_LL_DFPQX4 clk_r_REG331_S2 ( .D(n5543), .CP(clk), .Q(n8716) );
  HS65_LL_DFPQX4 clk_r_REG45_S2 ( .D(n5794), .CP(clk), .Q(n8715) );
  HS65_LL_DFPQX4 clk_r_REG309_S2 ( .D(n5594), .CP(clk), .Q(n8714) );
  HS65_LL_DFPQX4 clk_r_REG555_S2 ( .D(n5859), .CP(clk), .Q(n8713) );
  HS65_LL_DFPQX4 clk_r_REG425_S2 ( .D(n5848), .CP(clk), .Q(n8712) );
  HS65_LL_DFPQX4 clk_r_REG151_S2 ( .D(n5625), .CP(clk), .Q(n8711) );
  HS65_LL_DFPQX4 clk_r_REG459_S2 ( .D(n5647), .CP(clk), .Q(n8710) );
  HS65_LL_DFPQX4 clk_r_REG396_S1 ( .D(n8228), .CP(clk), .Q(n8709) );
  HS65_LL_DFPQX4 clk_r_REG322_S2 ( .D(n5744), .CP(clk), .Q(n8708) );
  HS65_LL_DFPQX4 clk_r_REG511_S2 ( .D(\u_DataPath/mem_writedata_out_i [12]), 
        .CP(clk), .Q(n8705) );
  HS65_LL_DFPQX4 clk_r_REG405_S1 ( .D(n8399), .CP(clk), .Q(n8702) );
  HS65_LL_DFPQX4 clk_r_REG72_S1 ( .D(n8277), .CP(clk), .Q(n8701) );
  HS65_LL_DFPQX4 clk_r_REG69_S1 ( .D(n8151), .CP(clk), .Q(n8700) );
  HS65_LL_DFPQX4 clk_r_REG76_S1 ( .D(n8410), .CP(clk), .Q(n8698) );
  HS65_LL_DFPQX4 clk_r_REG412_S1 ( .D(n8138), .CP(clk), .Q(n8697) );
  HS65_LL_DFPQX4 clk_r_REG120_S1 ( .D(n8205), .CP(clk), .Q(n8696) );
  HS65_LL_DFPQX4 clk_r_REG61_S1 ( .D(n8270), .CP(clk), .Q(n8695) );
  HS65_LL_DFPQX4 clk_r_REG141_S1 ( .D(n8191), .CP(clk), .Q(n8694) );
  HS65_LL_DFPQX4 clk_r_REG401_S1 ( .D(n8148), .CP(clk), .Q(n8693) );
  HS65_LL_DFPQX4 clk_r_REG80_S1 ( .D(n8209), .CP(clk), .Q(n8692) );
  HS65_LL_DFPQX4 clk_r_REG133_S1 ( .D(n8275), .CP(clk), .Q(n8691) );
  HS65_LL_DFPQX4 clk_r_REG125_S1 ( .D(n8200), .CP(clk), .Q(n8690) );
  HS65_LL_DFPQX4 clk_r_REG668_S7 ( .D(n7645), .CP(clk), .Q(n8689) );
  HS65_LL_DFPQX4 clk_r_REG684_S1 ( .D(n8313), .CP(clk), .Q(n8687) );
  HS65_LL_DFPQX4 clk_r_REG653_S5 ( .D(\u_DataPath/cw_exmem_i [9]), .CP(clk), 
        .Q(n8686) );
  HS65_LL_DFPQX4 clk_r_REG81_S1 ( .D(\u_DataPath/mem_writedata_out_i [23]), 
        .CP(clk), .Q(n8685) );
  HS65_LL_DFPQX4 clk_r_REG284_S3 ( .D(n8146), .CP(clk), .Q(n8684) );
  HS65_LL_DFPQX4 clk_r_REG520_S3 ( .D(\u_DataPath/data_read_ex_2_i [25]), .CP(
        clk), .Q(n8682) );
  HS65_LL_DFPQX4 clk_r_REG522_S2 ( .D(\u_DataPath/data_read_ex_2_i [22]), .CP(
        clk), .Q(n8681) );
  HS65_LL_DFPQX4 clk_r_REG104_S2 ( .D(\u_DataPath/data_read_ex_1_i [18]), .CP(
        clk), .Q(n8680) );
  HS65_LL_DFPQX4 clk_r_REG75_S3 ( .D(n8161), .CP(clk), .Q(n8679) );
  HS65_LL_DFPQX4 clk_r_REG71_S4 ( .D(n8299), .CP(clk), .Q(n8678) );
  HS65_LL_DFPQX4 clk_r_REG564_S5 ( .D(\u_DataPath/data_read_ex_1_i [0]), .CP(
        clk), .Q(n8677) );
  HS65_LL_DFPQX4 clk_r_REG471_S1 ( .D(\u_DataPath/data_read_ex_1_i [3]), .CP(
        clk), .Q(n8676) );
  HS65_LL_DFPQX4 clk_r_REG427_S2 ( .D(n8176), .CP(clk), .Q(n8675) );
  HS65_LL_DFPQX4 clk_r_REG493_S1 ( .D(\u_DataPath/data_read_ex_1_i [2]), .CP(
        clk), .Q(n8674) );
  HS65_LL_DFPQX4 clk_r_REG504_S1 ( .D(\u_DataPath/data_read_ex_2_i [4]), .CP(
        clk), .Q(n8673) );
  HS65_LL_DFPQX4 clk_r_REG402_S3 ( .D(\u_DataPath/data_read_ex_1_i [16]), .CP(
        clk), .Q(n8671) );
  HS65_LL_DFPQX4 clk_r_REG505_S1 ( .D(\u_DataPath/data_read_ex_1_i [4]), .CP(
        clk), .Q(n8670) );
  HS65_LL_DFPQX4 clk_r_REG559_S3 ( .D(\u_DataPath/data_read_ex_1_i [1]), .CP(
        clk), .Q(n8669) );
  HS65_LL_DFPQX4 clk_r_REG101_S3 ( .D(\u_DataPath/data_read_ex_1_i [11]), .CP(
        clk), .Q(n8668) );
  HS65_LL_DFPQX4 clk_r_REG143_S3 ( .D(\u_DataPath/data_read_ex_1_i [17]), .CP(
        clk), .Q(n8666) );
  HS65_LL_DFPQX4 clk_r_REG144_S2 ( .D(n8147), .CP(clk), .Q(n8665) );
  HS65_LL_DFPQX4 clk_r_REG84_S2 ( .D(n8246), .CP(clk), .Q(n8664) );
  HS65_LL_DFPQX4 clk_r_REG68_S2 ( .D(n8252), .CP(clk), .Q(n8663) );
  HS65_LL_DFPQX4 clk_r_REG66_S4 ( .D(n8238), .CP(clk), .Q(n8662) );
  HS65_LL_DFPQX4 clk_r_REG403_S3 ( .D(\u_DataPath/data_read_ex_2_i [16]), .CP(
        clk), .Q(n8661) );
  HS65_LL_DFPQX4 clk_r_REG414_S3 ( .D(\u_DataPath/data_read_ex_2_i [24]), .CP(
        clk), .Q(n8660) );
  HS65_LL_DFPQX4 clk_r_REG417_S2 ( .D(\u_DataPath/data_read_ex_2_i [18]), .CP(
        clk), .Q(n8659) );
  HS65_LL_DFPQX4 clk_r_REG126_S3 ( .D(\u_DataPath/data_read_ex_1_i [21]), .CP(
        clk), .Q(n8658) );
  HS65_LL_DFPQX4 clk_r_REG502_S3 ( .D(\u_DataPath/data_read_ex_1_i [13]), .CP(
        clk), .Q(n8656) );
  HS65_LL_DFPQX4 clk_r_REG301_S3 ( .D(n8174), .CP(clk), .Q(n8655) );
  HS65_LL_DFPQX4 clk_r_REG57_S2 ( .D(n8330), .CP(clk), .Q(n8654) );
  HS65_LL_DFPQX4 clk_r_REG581_S3 ( .D(\u_DataPath/data_read_ex_2_i [26]), .CP(
        clk), .Q(n8653) );
  HS65_LL_DFPQX4 clk_r_REG498_S2 ( .D(\u_DataPath/data_read_ex_2_i [30]), .CP(
        clk), .Q(n8652) );
  HS65_LL_DFPQX4 clk_r_REG500_S3 ( .D(\u_DataPath/data_read_ex_2_i [23]), .CP(
        clk), .Q(n8650) );
  HS65_LL_DFPQX4 clk_r_REG121_S3 ( .D(\u_DataPath/data_read_ex_2_i [27]), .CP(
        clk), .Q(n8649) );
  HS65_LL_DFPQX4 clk_r_REG518_S2 ( .D(\u_DataPath/data_read_ex_2_i [29]), .CP(
        clk), .Q(n8648) );
  HS65_LL_DFPQX4 clk_r_REG407_S2 ( .D(\u_DataPath/data_read_ex_2_i [9]), .CP(
        clk), .Q(n8647) );
  HS65_LL_DFPQX4 clk_r_REG545_S2 ( .D(\u_DataPath/data_read_ex_2_i [5]), .CP(
        clk), .Q(n8646) );
  HS65_LL_DFPQX4 clk_r_REG316_S3 ( .D(n8170), .CP(clk), .Q(n8645) );
  HS65_LL_DFPQX4 clk_r_REG248_S3 ( .D(n8139), .CP(clk), .Q(n8644) );
  HS65_LL_DFPQX4 clk_r_REG109_S2 ( .D(\u_DataPath/data_read_ex_1_i [31]), .CP(
        clk), .Q(n8642) );
  HS65_LL_DFPQX4 clk_r_REG579_S2 ( .D(\u_DataPath/data_read_ex_1_i [28]), .CP(
        clk), .Q(n8640) );
  HS65_LL_DFPQX4 clk_r_REG573_S5 ( .D(\u_DataPath/data_read_ex_2_i [0]), .CP(
        clk), .Q(n8639) );
  HS65_LL_DFPQX4 clk_r_REG508_S2 ( .D(\u_DataPath/data_read_ex_2_i [15]), .CP(
        clk), .Q(n8638) );
  HS65_LL_DFPQX4 clk_r_REG56_S2 ( .D(\u_DataPath/data_read_ex_1_i [22]), .CP(
        clk), .Q(n8637) );
  HS65_LL_DFPQX4 clk_r_REG495_S3 ( .D(\u_DataPath/data_read_ex_1_i [6]), .CP(
        clk), .Q(n8636) );
  HS65_LL_DFPQX4 clk_r_REG516_S3 ( .D(\u_DataPath/data_read_ex_1_i [10]), .CP(
        clk), .Q(n8635) );
  HS65_LL_DFPQX4 clk_r_REG408_S2 ( .D(\u_DataPath/data_read_ex_2_i [20]), .CP(
        clk), .Q(n8633) );
  HS65_LL_DFPQX4 clk_r_REG135_S2 ( .D(\u_DataPath/data_read_ex_1_i [20]), .CP(
        clk), .Q(n8632) );
  HS65_LL_DFPQX4 clk_r_REG406_S2 ( .D(\u_DataPath/data_read_ex_1_i [9]), .CP(
        clk), .Q(n8631) );
  HS65_LL_DFPQX4 clk_r_REG415_S3 ( .D(\u_DataPath/data_read_ex_2_i [21]), .CP(
        clk), .Q(n8630) );
  HS65_LL_DFPQX4 clk_r_REG507_S2 ( .D(\u_DataPath/data_read_ex_1_i [15]), .CP(
        clk), .Q(n8629) );
  HS65_LL_DFPQX4 clk_r_REG513_S3 ( .D(\u_DataPath/data_read_ex_1_i [12]), .CP(
        clk), .Q(n8628) );
  HS65_LL_DFPQX4 clk_r_REG59_S3 ( .D(\u_DataPath/data_read_ex_1_i [25]), .CP(
        clk), .Q(n8627) );
  HS65_LL_DFPQX4 clk_r_REG62_S2 ( .D(\u_DataPath/data_read_ex_1_i [29]), .CP(
        clk), .Q(n8625) );
  HS65_LL_DFPQX4 clk_r_REG611_S2 ( .D(\u_DataPath/data_read_ex_2_i [7]), .CP(
        clk), .Q(n8624) );
  HS65_LL_DFPQX4 clk_r_REG562_S3 ( .D(n8307), .CP(clk), .Q(n8623) );
  HS65_LL_DFPQX4 clk_r_REG692_S1 ( .D(n7969), .CP(clk), .Q(n8622) );
  HS65_LL_DFPQX4 clk_r_REG614_S5 ( .D(n7980), .CP(clk), .Q(n8621) );
  HS65_LL_DFPQX4 clk_r_REG210_S3 ( .D(n8287), .CP(clk), .Q(n8620) );
  HS65_LL_DFPQX4 clk_r_REG206_S2 ( .D(\u_DataPath/jump_address_i [30]), .CP(
        clk), .Q(n8619) );
  HS65_LL_DFPQX4 clk_r_REG166_S2 ( .D(\u_DataPath/jump_address_i [22]), .CP(
        clk), .Q(n8617) );
  HS65_LL_DFPQX4 clk_r_REG419_S4 ( .D(\u_DataPath/jump_address_i [3]), .CP(clk), .Q(n8616) );
  HS65_LL_DFPQX4 clk_r_REG379_S3 ( .D(\u_DataPath/jump_address_i [10]), .CP(
        clk), .Q(n8615) );
  HS65_LL_DFPQX4 clk_r_REG235_S2 ( .D(\u_DataPath/jump_address_i [26]), .CP(
        clk), .Q(n8614) );
  HS65_LL_DFPQX4 clk_r_REG323_S3 ( .D(\u_DataPath/jump_address_i [16]), .CP(
        clk), .Q(n8613) );
  HS65_LL_DFPQX4 clk_r_REG326_S4 ( .D(\u_DataPath/jump_address_i [14]), .CP(
        clk), .Q(n8612) );
  HS65_LL_DFPQX4 clk_r_REG409_S3 ( .D(\u_DataPath/data_read_ex_2_i [19]), .CP(
        clk), .Q(n8610) );
  HS65_LL_DFPQX4 clk_r_REG232_S3 ( .D(\u_DataPath/jump_address_i [24]), .CP(
        clk), .Q(n8609) );
  HS65_LL_DFPQX4 clk_r_REG273_S3 ( .D(\u_DataPath/jump_address_i [19]), .CP(
        clk), .Q(n8608) );
  HS65_LL_DFPQX4 clk_r_REG34_S3 ( .D(\u_DataPath/jump_address_i [7]), .CP(clk), 
        .Q(n8607) );
  HS65_LL_DFPQX4 clk_r_REG451_S3 ( .D(n8177), .CP(clk), .Q(n8606) );
  HS65_LL_DFPQX4 clk_r_REG597_S5 ( .D(n7960), .CP(clk), .Q(n8605) );
  HS65_LL_DFPQX4 clk_r_REG462_S3 ( .D(\u_DataPath/jump_address_i [4]), .CP(clk), .Q(n8604) );
  HS65_LL_DFPQX4 clk_r_REG685_S1 ( .D(n7988), .CP(clk), .Q(n8602) );
  HS65_LL_DFPQX4 clk_r_REG269_S3 ( .D(n8195), .CP(clk), .Q(n8598) );
  HS65_LL_DFPQX4 clk_r_REG250_S3 ( .D(n8210), .CP(clk), .Q(n8597) );
  HS65_LL_DFPQX4 clk_r_REG216_S3 ( .D(n7656), .CP(clk), .Q(n8596) );
  HS65_LL_DFPQX4 clk_r_REG257_S3 ( .D(n8201), .CP(clk), .Q(n8595) );
  HS65_LL_DFPQX4 clk_r_REG223_S3 ( .D(n8293), .CP(clk), .Q(n8594) );
  HS65_LL_DFPQX4 clk_r_REG296_S3 ( .D(n8192), .CP(clk), .Q(n8592) );
  HS65_LL_DFPQX4 clk_r_REG87_S3 ( .D(\u_DataPath/jump_address_i [2]), .CP(clk), 
        .Q(n8591) );
  HS65_LL_DFPQX4 clk_r_REG546_S3 ( .D(\u_DataPath/jump_address_i [1]), .CP(clk), .Q(n8590) );
  HS65_LL_DFPQX4 clk_r_REG565_S4 ( .D(\u_DataPath/jump_address_i [0]), .CP(clk), .Q(n8589) );
  HS65_LL_DFPQX4 clk_r_REG118_S3 ( .D(n8309), .CP(clk), .Q(n8588) );
  HS65_LL_DFPQX4 clk_r_REG678_S1 ( .D(\u_DataPath/cw_exmem_i [3]), .CP(clk), 
        .Q(n8587) );
  HS65_LL_DFPQX4 clk_r_REG687_S1 ( .D(n7996), .CP(clk), .Q(n8585) );
  HS65_LL_DFPQX4 clk_r_REG31_S2 ( .D(\u_DataPath/mem_writedata_out_i [5]), 
        .CP(clk), .Q(n8584) );
  HS65_LL_DFPQX4 clk_r_REG510_S4 ( .D(\u_DataPath/mem_writedata_out_i [14]), 
        .CP(clk), .Q(n8583) );
  HS65_LL_DFPQX4 clk_r_REG506_S2 ( .D(\u_DataPath/mem_writedata_out_i [15]), 
        .CP(clk), .Q(n8577) );
  HS65_LL_DFPQX4 clk_r_REG77_S1 ( .D(\u_DataPath/mem_writedata_out_i [13]), 
        .CP(clk), .Q(n8576) );
  HS65_LL_DFPQX4 clk_r_REG142_S1 ( .D(\u_DataPath/mem_writedata_out_i [17]), 
        .CP(clk), .Q(n8575) );
  HS65_LL_DFPQX4 clk_r_REG94_S1 ( .D(\u_DataPath/mem_writedata_out_i [3]), 
        .CP(clk), .Q(n8572) );
  HS65_LL_DFPQX4 clk_r_REG558_S2 ( .D(\u_DataPath/mem_writedata_out_i [1]), 
        .CP(clk), .Q(n8568) );
  HS65_LL_DFPQX4 clk_r_REG503_S1 ( .D(\u_DataPath/mem_writedata_out_i [4]), 
        .CP(clk), .Q(n8567) );
  HS65_LL_DFPQX4 clk_r_REG563_S1 ( .D(\u_DataPath/mem_writedata_out_i [0]), 
        .CP(clk), .Q(n8565) );
  HS65_LL_DFPQX4 clk_r_REG494_S1 ( .D(\u_DataPath/mem_writedata_out_i [6]), 
        .CP(clk), .Q(n8564) );
  HS65_LL_DFPQX4 clk_r_REG138_S3 ( .D(\u_DataPath/dataOut_exe_i [16]), .CP(clk), .Q(n8553) );
  HS65_LL_DFPQX4 clk_r_REG566_S4 ( .D(\u_DataPath/pc_4_i [0]), .CP(net3007), 
        .Q(n8547) );
  HS65_LL_DFPQX4 clk_r_REG547_S4 ( .D(\u_DataPath/pc_4_i [1]), .CP(net3007), 
        .Q(n8546) );
  HS65_LL_IVX27 U3584 ( .A(\u_DataPath/u_ifidreg/N61 ), .Z(n2811) );
  HS65_LL_IVX27 U3779 ( .A(\u_DataPath/u_ifidreg/N59 ), .Z(n2817) );
  HS65_LL_IVX27 U9372 ( .A(\u_DataPath/u_ifidreg/N57 ), .Z(n2815) );
  HS65_LL_IVX27 U9608 ( .A(\u_DataPath/u_memwbreg/N74 ), .Z(n7649) );
  HS65_LL_IVX27 U9609 ( .A(\u_DataPath/u_idexreg/N12 ), .Z(n2803) );
  HS65_LL_IVX27 U9825 ( .A(\u_DataPath/u_memwbreg/N70 ), .Z(n7647) );
  HS65_LL_IVX27 U9826 ( .A(\u_DataPath/u_memwbreg/N73 ), .Z(n7648) );
  HS65_LL_IVX27 U9827 ( .A(\u_DataPath/u_memwbreg/N45 ), .Z(n7675) );
  HS65_LL_IVX27 U9828 ( .A(\u_DataPath/u_memwbreg/N71 ), .Z(n7672) );
  HS65_LL_IVX27 U9829 ( .A(\u_DataPath/u_memwbreg/N72 ), .Z(n7673) );
  HS65_LL_DFPQX27 clk_r_REG655_S6 ( .D(n8310), .CP(clk), .Q(n9044) );
  HS65_LL_DFPQX35 clk_r_REG112_S4 ( .D(\u_DataPath/pc_4_i [31]), .CP(net3007), 
        .Q(n8969) );
  HS65_LH_DFPQX4 clk_r_REG675_S7 ( .D(n7643), .CP(clk), .Q(n2720) );
  HS65_LH_DFPQX4 clk_r_REG620_S5 ( .D(n8601), .CP(clk), .Q(n8600) );
  HS65_LH_DFPQX4 clk_r_REG599_S5 ( .D(n8707), .CP(clk), .Q(n8706) );
  HS65_LH_DFPQX4 clk_r_REG572_S3 ( .D(n9315), .CP(clk), .Q(n9314) );
  HS65_LH_DFPQX4 clk_r_REG424_S3 ( .D(n9073), .CP(clk), .Q(n9072) );
  HS65_LH_DFPQX4 clk_r_REG92_S3 ( .D(n8943), .CP(clk), .Q(n8942) );
  HS65_LH_DFPQX4 clk_r_REG28_S2 ( .D(n9178), .CP(clk), .Q(n9177) );
  HS65_LH_DFPQX4 clk_r_REG892_S5 ( .D(n9090), .CP(clk), .Q(n9089) );
  HS65_LH_DFPQX4 clk_r_REG906_S5 ( .D(n9311), .CP(clk), .Q(n9310) );
  HS65_LH_DFPQX4 clk_r_REG945_S6 ( .D(n9433), .CP(clk), .Q(n9432) );
  HS65_LH_DFPQX4 clk_r_REG889_S5 ( .D(n8990), .CP(clk), .Q(n8989) );
  HS65_LH_DFPQX4 clk_r_REG935_S2 ( .D(n9054), .CP(clk), .Q(n9053) );
  HS65_LH_DFPQX4 clk_r_REG899_S5 ( .D(n9052), .CP(clk), .Q(n9051) );
  HS65_LH_DFPQX4 clk_r_REG895_S5 ( .D(n8901), .CP(clk), .Q(n8900) );
  HS65_LH_DFPQX4 clk_r_REG908_S5 ( .D(n8801), .CP(clk), .Q(n8800) );
  HS65_LH_DFPQX4 clk_r_REG933_S5 ( .D(n9422), .CP(clk), .Q(n9421) );
  HS65_LH_DFPQX4 clk_r_REG683_S2 ( .D(n9445), .CP(clk), .Q(n9444) );
  HS65_LH_DFPQX4 clk_r_REG936_S5 ( .D(n8817), .CP(clk), .Q(n8816) );
  HS65_LH_DFPQX4 clk_r_REG0_S1 ( .D(n1885), .CP(clk), .Q(n9504) );
  HS65_LH_DFPQX4 clk_r_REG976_S1 ( .D(Data_out_fromRAM[0]), .CP(clk), .Q(n9476) );
  HS65_LH_DFPQX4 clk_r_REG975_S1 ( .D(Data_out_fromRAM[1]), .CP(clk), .Q(n9477) );
  HS65_LH_DFPQX4 clk_r_REG974_S1 ( .D(Data_out_fromRAM[2]), .CP(clk), .Q(n9478) );
  HS65_LH_DFPQX4 clk_r_REG973_S1 ( .D(Data_out_fromRAM[3]), .CP(clk), .Q(n9479) );
  HS65_LH_DFPQX4 clk_r_REG972_S1 ( .D(Data_out_fromRAM[4]), .CP(clk), .Q(n9480) );
  HS65_LH_DFPQX4 clk_r_REG971_S1 ( .D(Data_out_fromRAM[5]), .CP(clk), .Q(n9481) );
  HS65_LH_DFPQX4 clk_r_REG970_S1 ( .D(Data_out_fromRAM[6]), .CP(clk), .Q(n9482) );
  HS65_LH_DFPQX4 clk_r_REG962_S1 ( .D(Data_out_fromRAM[16]), .CP(clk), .Q(
        n9490) );
  HS65_LH_DFPQX4 clk_r_REG961_S1 ( .D(Data_out_fromRAM[17]), .CP(clk), .Q(
        n9491) );
  HS65_LH_DFPQX4 clk_r_REG960_S1 ( .D(Data_out_fromRAM[18]), .CP(clk), .Q(
        n9492) );
  HS65_LH_DFPQX4 clk_r_REG959_S1 ( .D(Data_out_fromRAM[19]), .CP(clk), .Q(
        n9493) );
  HS65_LH_DFPQX4 clk_r_REG958_S1 ( .D(Data_out_fromRAM[20]), .CP(clk), .Q(
        n9494) );
  HS65_LH_DFPQX4 clk_r_REG957_S1 ( .D(Data_out_fromRAM[21]), .CP(clk), .Q(
        n9495) );
  HS65_LH_DFPQX4 clk_r_REG956_S1 ( .D(Data_out_fromRAM[22]), .CP(clk), .Q(
        n9496) );
  HS65_LH_DFPQX4 clk_r_REG955_S1 ( .D(Data_out_fromRAM[24]), .CP(clk), .Q(
        n9497) );
  HS65_LH_DFPQX4 clk_r_REG954_S1 ( .D(Data_out_fromRAM[25]), .CP(clk), .Q(
        n9498) );
  HS65_LH_DFPQX4 clk_r_REG953_S1 ( .D(Data_out_fromRAM[26]), .CP(clk), .Q(
        n9499) );
  HS65_LH_DFPQX4 clk_r_REG952_S1 ( .D(Data_out_fromRAM[27]), .CP(clk), .Q(
        n9500) );
  HS65_LH_DFPQX4 clk_r_REG951_S1 ( .D(Data_out_fromRAM[28]), .CP(clk), .Q(
        n9501) );
  HS65_LH_DFPQX4 clk_r_REG950_S1 ( .D(Data_out_fromRAM[29]), .CP(clk), .Q(
        n9502) );
  HS65_LH_DFPQX4 clk_r_REG949_S1 ( .D(Data_out_fromRAM[30]), .CP(clk), .Q(
        n9503) );
  HS65_LH_DFPQX4 clk_r_REG969_S1 ( .D(Data_out_fromRAM[8]), .CP(clk), .Q(n9483) );
  HS65_LH_DFPQX4 clk_r_REG968_S1 ( .D(Data_out_fromRAM[9]), .CP(clk), .Q(n9484) );
  HS65_LH_DFPQX4 clk_r_REG967_S1 ( .D(Data_out_fromRAM[10]), .CP(clk), .Q(
        n9485) );
  HS65_LH_DFPQX4 clk_r_REG966_S1 ( .D(Data_out_fromRAM[11]), .CP(clk), .Q(
        n9486) );
  HS65_LH_DFPQX4 clk_r_REG965_S1 ( .D(Data_out_fromRAM[12]), .CP(clk), .Q(
        n9487) );
  HS65_LH_DFPQX4 clk_r_REG964_S1 ( .D(Data_out_fromRAM[13]), .CP(clk), .Q(
        n9488) );
  HS65_LH_DFPQX4 clk_r_REG963_S1 ( .D(Data_out_fromRAM[14]), .CP(clk), .Q(
        n9489) );
  HS65_LH_DFPQX4 clk_r_REG909_S5 ( .D(n7994), .CP(clk), .Q(n9400) );
  HS65_LH_DFPQX4 clk_r_REG286_S3 ( .D(\u_DataPath/u_execute/link_value_i [18]), 
        .CP(clk), .Q(n9117) );
  HS65_LH_DFPQX4 clk_r_REG551_S1 ( .D(\u_DataPath/branch_target_i [1]), .CP(
        clk), .Q(n8834) );
  HS65_LH_DFPQX4 clk_r_REG27_S1 ( .D(\u_DataPath/u_execute/psw_status_i [1]), 
        .CP(clk), .Q(n9178) );
  HS65_LH_DFPQX4 clk_r_REG571_S1 ( .D(\u_DataPath/branch_target_i [0]), .CP(
        clk), .Q(n9395) );
  HS65_LH_DFPQX4 clk_r_REG487_S1 ( .D(\u_DataPath/branch_target_i [2]), .CP(
        clk), .Q(n8832) );
  HS65_LH_DFPQX4 clk_r_REG491_S1 ( .D(n2971), .CP(clk), .Q(n9457) );
  HS65_LH_DFPQX4 clk_r_REG557_S1 ( .D(n8461), .CP(clk), .Q(n8878) );
  HS65_LH_DFPQX4 clk_r_REG641_S6 ( .D(\u_DataPath/cw_memwb_i [0]), .CP(clk), 
        .Q(n9349) );
  HS65_LH_DFPQX4 clk_r_REG934_S1 ( .D(n8465), .CP(clk), .Q(n9054) );
  HS65_LH_DFPQX4 clk_r_REG656_S6 ( .D(n8315), .CP(clk), .Q(n9278) );
  HS65_LH_DFPQX4 clk_r_REG902_S1 ( .D(n8500), .CP(clk), .Q(n9137) );
  HS65_LH_DFPQX4 clk_r_REG30_S1 ( .D(\u_DataPath/from_alu_data_out_i [5]), 
        .CP(clk), .Q(n8795) );
  HS65_LH_DFPQX4 clk_r_REG896_S1 ( .D(n8498), .CP(clk), .Q(n9135) );
  HS65_LH_DFPQX4 clk_r_REG657_S6 ( .D(\u_DataPath/cw_memwb_i [1]), .CP(clk), 
        .Q(n9176) );
  HS65_LH_DFPQX4 clk_r_REG85_S1 ( .D(\u_DataPath/from_alu_data_out_i [6]), 
        .CP(clk), .Q(n8794) );
  HS65_LH_DFPQX4 clk_r_REG907_S1 ( .D(n8466), .CP(clk), .Q(n9134) );
  HS65_LH_DFPQX4 clk_r_REG604_S1 ( .D(\u_DataPath/reg_write_i ), .CP(clk), .Q(
        n9175) );
  HS65_LH_DFPQX4 clk_r_REG93_S1 ( .D(\u_DataPath/from_alu_data_out_i [3]), 
        .CP(clk), .Q(n8796) );
  HS65_LH_DFPQX4 clk_r_REG717_S2 ( .D(\u_DataPath/cw_tomem_i [6]), .CP(clk), 
        .Q(n9350) );
  HS65_LH_DFPQX4 clk_r_REG927_S5 ( .D(n8523), .CP(clk), .Q(n9427) );
  HS65_LH_DFPQX4 clk_r_REG947_S5 ( .D(n8525), .CP(clk), .Q(n9431) );
  HS65_LH_DFPQX4 clk_r_REG801_S1 ( .D(\u_DataPath/idex_rt_i [3]), .CP(clk), 
        .Q(n9112) );
  HS65_LH_DFPQX4 clk_r_REG923_S5 ( .D(n8504), .CP(clk), .Q(n9434) );
  HS65_LH_DFPQX4 clk_r_REG715_S1 ( .D(\u_DataPath/cw_tomem_i [4]), .CP(clk), 
        .Q(n9110) );
  HS65_LH_DFPQX4 clk_r_REG942_S5 ( .D(n8474), .CP(clk), .Q(n9428) );
  HS65_LH_DFPQX4 clk_r_REG940_S5 ( .D(n8524), .CP(clk), .Q(n9429) );
  HS65_LH_DFPQX4 clk_r_REG944_S5 ( .D(n8469), .CP(clk), .Q(n9433) );
  HS65_LH_DFPQX4 clk_r_REG568_S2 ( .D(\u_DataPath/u_execute/link_value_i [0]), 
        .CP(clk), .Q(n9315) );
  HS65_LH_DFPQX4 clk_r_REG930_S5 ( .D(n8506), .CP(clk), .Q(n9436) );
  HS65_LH_DFPQX4 clk_r_REG925_S5 ( .D(n8510), .CP(clk), .Q(n9435) );
  HS65_LH_DFPQX4 clk_r_REG708_S1 ( .D(n7649), .CP(clk), .Q(n9170) );
  HS65_LH_DFPQX4 clk_r_REG702_S1 ( .D(n7673), .CP(clk), .Q(n9173) );
  HS65_LH_DFPQX4 clk_r_REG114_S2 ( .D(\u_DataPath/pc_4_to_ex_i [31]), .CP(clk), 
        .Q(n9355) );
  HS65_LH_DFPQX4 clk_r_REG549_S2 ( .D(\u_DataPath/u_execute/link_value_i [1]), 
        .CP(clk), .Q(n9348) );
  HS65_LH_DFPQX4 clk_r_REG699_S1 ( .D(n7647), .CP(clk), .Q(n9172) );
  HS65_LH_DFPQX4 clk_r_REG900_S5 ( .D(n7978), .CP(clk), .Q(n8723) );
  HS65_LH_DFPQX4 clk_r_REG664_S7 ( .D(n8028), .CP(clk), .Q(n9058) );
  HS65_LH_DFPQX4 clk_r_REG670_S7 ( .D(n8029), .CP(clk), .Q(n9061) );
  HS65_LH_DFPQX4 clk_r_REG916_S5 ( .D(n8508), .CP(clk), .Q(n9452) );
  HS65_LH_DFPQX4 clk_r_REG914_S1 ( .D(n8467), .CP(clk), .Q(n8818) );
  HS65_LH_DFPQX4 clk_r_REG476_S1 ( .D(\u_DataPath/branch_target_i [3]), .CP(
        clk), .Q(n9365) );
  HS65_LH_DFPQX4 clk_r_REG666_S7 ( .D(n6488), .CP(clk), .Q(n9059) );
  HS65_LH_DFPQX4 clk_r_REG696_S1 ( .D(\u_DataPath/regfile_addr_out_towb_i [3]), 
        .CP(clk), .Q(n9270) );
  HS65_LH_DFPQX4 clk_r_REG200_S2 ( .D(\u_DataPath/pc_4_to_ex_i [30]), .CP(clk), 
        .Q(n9356) );
  HS65_LH_DFPQX4 clk_r_REG193_S2 ( .D(\u_DataPath/pc_4_to_ex_i [29]), .CP(clk), 
        .Q(n9357) );
  HS65_LH_DFPQX4 clk_r_REG709_S1 ( .D(\u_DataPath/regfile_addr_out_towb_i [4]), 
        .CP(clk), .Q(n9233) );
  HS65_LH_DFPQX4 clk_r_REG672_S7 ( .D(n7014), .CP(clk), .Q(n9092) );
  HS65_LH_DFPQX4 clk_r_REG679_S1 ( .D(n8162), .CP(clk), .Q(n9286) );
  HS65_LH_DFPQX4 clk_r_REG18_S2 ( .D(\u_DataPath/pc_4_to_ex_i [26]), .CP(clk), 
        .Q(n9354) );
  HS65_LH_DFPQX4 clk_r_REG881_S1 ( .D(\u_DataPath/idex_rt_i [2]), .CP(clk), 
        .Q(n9046) );
  HS65_LH_DFPQX4 clk_r_REG170_S2 ( .D(\u_DataPath/pc_4_to_ex_i [24]), .CP(clk), 
        .Q(n9353) );
  HS65_LH_DFPQX4 clk_r_REG52_S2 ( .D(\u_DataPath/pc_4_to_ex_i [22]), .CP(clk), 
        .Q(n9352) );
  HS65_LH_DFPQX4 clk_r_REG186_S2 ( .D(\u_DataPath/pc_4_to_ex_i [28]), .CP(clk), 
        .Q(n9361) );
  HS65_LH_DFPQX4 clk_r_REG878_S1 ( .D(\u_DataPath/idex_rt_i [4]), .CP(clk), 
        .Q(n8906) );
  HS65_LH_DFPQX4 clk_r_REG404_S3 ( .D(\u_DataPath/mem_writedata_out_i [9]), 
        .CP(clk), .Q(n8643) );
  HS65_LH_DFPQX4 clk_r_REG600_S6 ( .D(\u_DataPath/cw_memwb_i [2]), .CP(clk), 
        .Q(n9313) );
  HS65_LH_DFPQX4 clk_r_REG883_S1 ( .D(\u_DataPath/idex_rt_i [1]), .CP(clk), 
        .Q(n8819) );
  HS65_LH_DFPQX4 clk_r_REG700_S1 ( .D(n7015), .CP(clk), .Q(n9225) );
  HS65_LH_DFPQX4 clk_r_REG918_S5 ( .D(n8512), .CP(clk), .Q(n9360) );
  HS65_LH_DFPQX4 clk_r_REG703_S1 ( .D(n7216), .CP(clk), .Q(n9335) );
  HS65_LH_DFPQX4 clk_r_REG519_S1 ( .D(\u_DataPath/mem_writedata_out_i [29]), 
        .CP(clk), .Q(n9121) );
  HS65_LH_DFPQX4 clk_r_REG386_S2 ( .D(\u_DataPath/pc_4_to_ex_i [8]), .CP(clk), 
        .Q(n9358) );
  HS65_LH_DFPQX4 clk_r_REG411_S1 ( .D(\u_DataPath/mem_writedata_out_i [24]), 
        .CP(clk), .Q(n9123) );
  HS65_LH_DFPQX4 clk_r_REG38_S2 ( .D(\u_DataPath/pc_4_to_ex_i [10]), .CP(clk), 
        .Q(n9359) );
  HS65_LH_DFPQX4 clk_r_REG122_S1 ( .D(\u_DataPath/mem_writedata_out_i [27]), 
        .CP(clk), .Q(n9106) );
  HS65_LH_DFPQX4 clk_r_REG665_S7 ( .D(n8006), .CP(clk), .Q(n9184) );
  HS65_LH_DFPQX4 clk_r_REG671_S7 ( .D(n8003), .CP(clk), .Q(n9183) );
  HS65_LH_DFPQX4 clk_r_REG97_S1 ( .D(\u_DataPath/mem_writedata_out_i [11]), 
        .CP(clk), .Q(n8566) );
  HS65_LH_DFPQX4 clk_r_REG416_S4 ( .D(\u_DataPath/mem_writedata_out_i [21]), 
        .CP(clk), .Q(n8570) );
  HS65_LH_DFPQX4 clk_r_REG134_S2 ( .D(\u_DataPath/mem_writedata_out_i [20]), 
        .CP(clk), .Q(n8571) );
  HS65_LH_DFPQX4 clk_r_REG300_S1 ( .D(\u_DataPath/mem_writedata_out_i [8]), 
        .CP(clk), .Q(n8574) );
  HS65_LH_DFPQX4 clk_r_REG6_S3 ( .D(\u_DataPath/mem_writedata_out_i [7]), .CP(
        clk), .Q(n8578) );
  HS65_LH_DFPQX4 clk_r_REG65_S1 ( .D(\u_DataPath/mem_writedata_out_i [10]), 
        .CP(clk), .Q(n8573) );
  HS65_LH_DFPQX4 clk_r_REG139_S4 ( .D(\u_DataPath/mem_writedata_out_i [16]), 
        .CP(clk), .Q(n8579) );
  HS65_LH_DFPQX4 clk_r_REG130_S2 ( .D(\u_DataPath/mem_writedata_out_i [19]), 
        .CP(clk), .Q(n8580) );
  HS65_LH_DFPQX4 clk_r_REG523_S3 ( .D(\u_DataPath/mem_writedata_out_i [22]), 
        .CP(clk), .Q(n8581) );
  HS65_LH_DFPQX4 clk_r_REG256_S2 ( .D(n7632), .CP(clk), .Q(n9295) );
  HS65_LH_DFPQX4 clk_r_REG249_S2 ( .D(n7628), .CP(clk), .Q(n9292) );
  HS65_LH_DFPQX4 clk_r_REG2_S2 ( .D(\u_DataPath/u_execute/psw_status_i [0]), 
        .CP(clk), .Q(n8563) );
  HS65_LH_DFPQX4 clk_r_REG229_S2 ( .D(n7634), .CP(clk), .Q(n9293) );
  HS65_LH_DFPQX4 clk_r_REG921_S1 ( .D(n8522), .CP(clk), .Q(n9143) );
  HS65_LH_DFPSQX4 clk_r_REG725_S4 ( .D(opcode_i[4]), .CP(net3007), .SN(n7677), 
        .Q(n9118) );
  HS65_LH_DFPSQX4 clk_r_REG932_S4 ( .D(n8030), .CP(net3007), .SN(n2814), .Q(
        n9422) );
  HS65_LH_DFPSQX4 clk_r_REG920_S4 ( .D(n8077), .CP(net3007), .SN(n9554), .Q(
        n9389) );
  HS65_LH_DFPSQX4 clk_r_REG911_S4 ( .D(n7604), .CP(net3007), .SN(n9546), .Q(
        n9179) );
  HS65_LH_DFPSQX4 clk_r_REG905_S4 ( .D(n8031), .CP(net3007), .SN(n2814), .Q(
        n9311) );
  HS65_LH_DFPSQX4 clk_r_REG904_S4 ( .D(n7347), .CP(net3007), .SN(n2814), .Q(
        n8845) );
  HS65_LH_DFPSQX4 clk_r_REG938_S4 ( .D(n7965), .CP(net3007), .SN(n9557), .Q(
        n9303) );
  HS65_LH_DFPSQX4 clk_r_REG800_S4 ( .D(n7931), .CP(net3007), .SN(n9548), .Q(
        n9236) );
  HS65_LH_DFPSQX4 clk_r_REG912_S4 ( .D(n7412), .CP(net3007), .SN(n9555), .Q(
        n8898) );
  HS65_LH_DFPSQX4 clk_r_REG893_S4 ( .D(n8053), .CP(net3007), .SN(n2814), .Q(
        n9420) );
  HS65_LH_DFPSQX4 clk_r_REG869_S4 ( .D(n6479), .CP(net3007), .SN(n9557), .Q(
        n9467) );
  HS65_LH_DFPSQX4 clk_r_REG901_S4 ( .D(n8051), .CP(net3007), .SN(n2814), .Q(
        n9419) );
  HS65_LH_DFPSQX4 clk_r_REG888_S4 ( .D(n7982), .CP(net3007), .SN(n2814), .Q(
        n8990) );
  HS65_LH_DFPSQX4 clk_r_REG880_S4 ( .D(n8016), .CP(net3007), .SN(n9557), .Q(
        n9465) );
  HS65_LH_DFPSQX4 clk_r_REG877_S4 ( .D(n8017), .CP(net3007), .SN(n9557), .Q(
        n9384) );
  HS65_LH_DFPSQX4 clk_r_REG871_S4 ( .D(n8070), .CP(net3007), .SN(n9547), .Q(
        n8994) );
  HS65_LH_DFPSQX4 clk_r_REG891_S4 ( .D(n7350), .CP(net3007), .SN(n2814), .Q(
        n9182) );
  HS65_LH_DFPSQX4 clk_r_REG724_S4 ( .D(n7930), .CP(net3007), .SN(n9546), .Q(
        n9111) );
  HS65_LH_DFPSQX4 clk_r_REG719_S4 ( .D(n7934), .CP(net3007), .SN(n9554), .Q(
        n8739) );
  HS65_LH_DFPSQX4 clk_r_REG720_S4 ( .D(n7957), .CP(net3007), .SN(n9557), .Q(
        n8750) );
  HS65_LH_DFPSQX4 clk_r_REG623_S4 ( .D(n8072), .CP(net3007), .SN(n9545), .Q(
        n8703) );
  HS65_LH_DFPSQX4 clk_r_REG847_S4 ( .D(n6635), .CP(net3007), .SN(n9545), .Q(
        n9226) );
  HS65_LH_DFPSQX4 clk_r_REG722_S4 ( .D(n8020), .CP(net3007), .SN(n9548), .Q(
        n8725) );
  HS65_LH_DFPSQX4 clk_r_REG628_S4 ( .D(n7966), .CP(net3007), .SN(n9549), .Q(
        n8954) );
  HS65_LH_DFPSQX4 clk_r_REG621_S4 ( .D(n7951), .CP(net3007), .SN(n9545), .Q(
        n8586) );
  HS65_LH_DFPRQX4 clk_r_REG185_S1 ( .D(\u_DataPath/pc4_to_idexreg_i [28]), 
        .CP(net3007), .RN(n2814), .Q(n9447) );
  HS65_LH_DFPRQX4 clk_r_REG169_S1 ( .D(\u_DataPath/pc4_to_idexreg_i [24]), 
        .CP(net3007), .RN(n9549), .Q(n9372) );
  HS65_LH_DFPRQX4 clk_r_REG147_S1 ( .D(\u_DataPath/pc4_to_idexreg_i [17]), 
        .CP(net3007), .RN(n9549), .Q(n9405) );
  HS65_LH_DFPRQX4 clk_r_REG199_S1 ( .D(\u_DataPath/pc4_to_idexreg_i [30]), 
        .CP(net3007), .RN(n9549), .Q(n9327) );
  HS65_LH_DFPRQX4 clk_r_REG329_S1 ( .D(\u_DataPath/pc4_to_idexreg_i [15]), 
        .CP(net3007), .RN(n9549), .Q(n9451) );
  HS65_LH_DFPRQX4 clk_r_REG17_S1 ( .D(\u_DataPath/pc4_to_idexreg_i [26]), .CP(
        net3007), .RN(n9555), .Q(n9454) );
  HS65_LH_DFPRQX4 clk_r_REG342_S1 ( .D(\u_DataPath/pc4_to_idexreg_i [14]), 
        .CP(net3007), .RN(n9549), .Q(n9279) );
  HS65_LH_DFPRQX4 clk_r_REG319_S1 ( .D(\u_DataPath/pc4_to_idexreg_i [13]), 
        .CP(net3007), .RN(n9550), .Q(n9368) );
  HS65_LH_DFPRQX4 clk_r_REG267_S1 ( .D(\u_DataPath/pc4_to_idexreg_i [19]), 
        .CP(net3007), .RN(n9550), .Q(n9369) );
  HS65_LH_DFPRQX4 clk_r_REG155_S1 ( .D(\u_DataPath/pc4_to_idexreg_i [20]), 
        .CP(net3007), .RN(n9550), .Q(n9370) );
  HS65_LH_DFPRQX4 clk_r_REG51_S1 ( .D(\u_DataPath/pc4_to_idexreg_i [22]), .CP(
        net3007), .RN(n9549), .Q(n9371) );
  HS65_LH_DFPRQX4 clk_r_REG385_S1 ( .D(\u_DataPath/pc4_to_idexreg_i [8]), .CP(
        net3007), .RN(n9556), .Q(n9442) );
  HS65_LH_DFPRQX4 clk_r_REG481_S1 ( .D(\u_DataPath/pc4_to_idexreg_i [2]), .CP(
        net3007), .RN(n9551), .Q(n8833) );
  HS65_LH_DFPRQX4 clk_r_REG454_S1 ( .D(\u_DataPath/pc4_to_idexreg_i [5]), .CP(
        net3007), .RN(n9550), .Q(n8788) );
  HS65_LH_DFPRQX4 clk_r_REG440_S1 ( .D(\u_DataPath/pc4_to_idexreg_i [6]), .CP(
        net3007), .RN(n9551), .Q(n8830) );
  HS65_LH_DFPRQX4 clk_r_REG365_S1 ( .D(\u_DataPath/pc4_to_idexreg_i [11]), 
        .CP(net3007), .RN(n9550), .Q(n8786) );
  HS65_LH_DFPRQX4 clk_r_REG314_S1 ( .D(\u_DataPath/pc4_to_idexreg_i [12]), 
        .CP(net3007), .RN(n9551), .Q(n8827) );
  HS65_LH_DFPRQX4 clk_r_REG304_S1 ( .D(\u_DataPath/pc4_to_idexreg_i [9]), .CP(
        net3007), .RN(n9550), .Q(n8785) );
  HS65_LH_DFPRQX4 clk_r_REG281_S1 ( .D(\u_DataPath/pc4_to_idexreg_i [18]), 
        .CP(net3007), .RN(n9554), .Q(n8824) );
  HS65_LH_DFPRQX4 clk_r_REG240_S1 ( .D(\u_DataPath/pc4_to_idexreg_i [23]), 
        .CP(net3007), .RN(n9550), .Q(n8784) );
  HS65_LH_DFPRQX4 clk_r_REG192_S1 ( .D(\u_DataPath/pc4_to_idexreg_i [29]), 
        .CP(net3007), .RN(n9551), .Q(n8843) );
  HS65_LH_DFPRQX4 clk_r_REG179_S1 ( .D(\u_DataPath/pc4_to_idexreg_i [27]), 
        .CP(net3007), .RN(n9550), .Q(n8782) );
  HS65_LH_DFPRQX4 clk_r_REG162_S1 ( .D(\u_DataPath/pc4_to_idexreg_i [21]), 
        .CP(net3007), .RN(n2814), .Q(n8783) );
  HS65_LH_DFPRQX4 clk_r_REG44_S1 ( .D(\u_DataPath/pc4_to_idexreg_i [16]), .CP(
        net3007), .RN(n9551), .Q(n8835) );
  HS65_LH_DFPRQX4 clk_r_REG11_S1 ( .D(\u_DataPath/pc4_to_idexreg_i [25]), .CP(
        net3007), .RN(n9550), .Q(n8826) );
  HS65_LH_DFPRQX4 clk_r_REG430_S1 ( .D(\u_DataPath/pc4_to_idexreg_i [7]), .CP(
        net3007), .RN(n9556), .Q(n9441) );
  HS65_LH_DFPRQX4 clk_r_REG37_S1 ( .D(\u_DataPath/pc4_to_idexreg_i [10]), .CP(
        net3007), .RN(n9556), .Q(n9440) );
  HS65_LH_DFPRQX4 clk_r_REG113_S1 ( .D(\u_DataPath/pc4_to_idexreg_i [31]), 
        .CP(net3007), .RN(n9551), .Q(n8879) );
  HS65_LH_DFPRQX4 clk_r_REG567_S1 ( .D(\u_DataPath/pc4_to_idexreg_i [0]), .CP(
        net3007), .RN(n9549), .Q(n9344) );
  HS65_LH_DFPRQX4 clk_r_REG548_S1 ( .D(\u_DataPath/pc4_to_idexreg_i [1]), .CP(
        net3007), .RN(n9556), .Q(n9345) );
  HS65_LH_DFPRQX4 clk_r_REG422_S1 ( .D(\u_DataPath/pc4_to_idexreg_i [4]), .CP(
        net3007), .RN(n9554), .Q(n9439) );
  HS65_LH_DFPRQX4 clk_r_REG90_S1 ( .D(\u_DataPath/pc4_to_idexreg_i [3]), .CP(
        net3007), .RN(n9549), .Q(n9399) );
  HS65_LH_DFPRQX4 clk_r_REG946_S4 ( .D(\u_DataPath/immediate_ext_dec_i [9]), 
        .CP(net3007), .RN(n9556), .Q(n8793) );
  HS65_LH_DFPRQX4 clk_r_REG943_S4 ( .D(\u_DataPath/immediate_ext_dec_i [10]), 
        .CP(net3007), .RN(n9550), .Q(n8792) );
  HS65_LH_DFPRQX4 clk_r_REG941_S4 ( .D(\u_DataPath/immediate_ext_dec_i [7]), 
        .CP(net3007), .RN(n2814), .Q(n8791) );
  HS65_LH_DFPRQX4 clk_r_REG939_S4 ( .D(\u_DataPath/immediate_ext_dec_i [8]), 
        .CP(net3007), .RN(n9550), .Q(n8790) );
  HS65_LH_DFPRQX4 clk_r_REG929_S4 ( .D(\u_DataPath/immediate_ext_dec_i [11]), 
        .CP(net3007), .RN(n9554), .Q(n8815) );
  HS65_LH_DFPRQX4 clk_r_REG924_S4 ( .D(\u_DataPath/immediate_ext_dec_i [13]), 
        .CP(net3007), .RN(n9554), .Q(n8809) );
  HS65_LH_DFPRQX4 clk_r_REG922_S4 ( .D(\u_DataPath/immediate_ext_dec_i [14]), 
        .CP(net3007), .RN(n9554), .Q(n8808) );
  HS65_LH_DFPRQX4 clk_r_REG917_S4 ( .D(\u_DataPath/immediate_ext_dec_i [15]), 
        .CP(net3007), .RN(n9554), .Q(n8804) );
  HS65_LH_DFPRQX4 clk_r_REG915_S4 ( .D(\u_DataPath/immediate_ext_dec_i [12]), 
        .CP(net3007), .RN(n9550), .Q(n8803) );
  HS65_LH_DFPRQX4 clk_r_REG926_S4 ( .D(\u_DataPath/immediate_ext_dec_i [6]), 
        .CP(net3007), .RN(n2814), .Q(n8814) );
  HS65_LH_DFPRQX4 clk_r_REG931_S4 ( .D(\u_DataPath/immediate_ext_dec_i [2]), 
        .CP(net3007), .RN(n2814), .Q(n8817) );
  HS65_LH_DFPRQX4 clk_r_REG919_S4 ( .D(\u_DataPath/immediate_ext_dec_i [5]), 
        .CP(net3007), .RN(n9551), .Q(n8806) );
  HS65_LH_DFPRQX4 clk_r_REG910_S4 ( .D(\u_DataPath/immediate_ext_dec_i [4]), 
        .CP(net3007), .RN(n9550), .Q(n8802) );
  HS65_LH_DFPRQX4 clk_r_REG903_S4 ( .D(\u_DataPath/immediate_ext_dec_i [3]), 
        .CP(net3007), .RN(n2814), .Q(n8801) );
  HS65_LH_DFPRQX4 clk_r_REG937_S4 ( .D(opcode_i[5]), .CP(net3007), .RN(n9550), 
        .Q(n8789) );
  HS65_LH_DFPRQX4 clk_r_REG887_S4 ( .D(\u_DataPath/immediate_ext_dec_i [1]), 
        .CP(net3007), .RN(n2814), .Q(n8798) );
  HS65_LH_DFPRQX4 clk_r_REG799_S4 ( .D(n2804), .CP(net3007), .RN(n9555), .Q(
        n9464) );
  HS65_LH_DFPRQX4 clk_r_REG886_S4 ( .D(n2816), .CP(net3007), .RN(n9549), .Q(
        n9385) );
  HS65_LH_DFPRQX4 clk_r_REG868_S4 ( .D(\u_DataPath/jaddr_i [22]), .CP(net3007), 
        .RN(n9554), .Q(n8805) );
  HS65_LH_DFPRQX4 clk_r_REG897_S4 ( .D(\u_DataPath/immediate_ext_dec_i [0]), 
        .CP(net3007), .RN(n2814), .Q(n8799) );
  HS65_LH_DFPRQX4 clk_r_REG873_S4 ( .D(n2818), .CP(net3007), .RN(n9555), .Q(
        n9466) );
  HS65_LH_DFPRQX4 clk_r_REG879_S4 ( .D(\u_DataPath/jaddr_i [18]), .CP(net3007), 
        .RN(n9554), .Q(n8812) );
  HS65_LH_DFPRQX4 clk_r_REG731_S4 ( .D(\u_DataPath/jaddr_i [16]), .CP(net3007), 
        .RN(n9550), .Q(n8797) );
  HS65_LH_DFPRQX4 clk_r_REG882_S4 ( .D(\u_DataPath/jaddr_i [17]), .CP(net3007), 
        .RN(n9554), .Q(n8813) );
  HS65_LH_DFPRQX4 clk_r_REG876_S4 ( .D(\u_DataPath/jaddr_i [20]), .CP(net3007), 
        .RN(n9554), .Q(n8811) );
  HS65_LH_DFPRQX4 clk_r_REG835_S4 ( .D(n2812), .CP(net3007), .RN(n9555), .Q(
        n9462) );
  HS65_LH_DFPRQX4 clk_r_REG870_S4 ( .D(opcode_i[3]), .CP(net3007), .RN(n9554), 
        .Q(n8807) );
  HS65_LH_DFPRQX4 clk_r_REG898_S4 ( .D(n7954), .CP(net3007), .RN(n2814), .Q(
        n9052) );
  HS65_LH_DFPRQX4 clk_r_REG874_S4 ( .D(\u_DataPath/jaddr_i [24]), .CP(net3007), 
        .RN(n9554), .Q(n8810) );
  HS65_LH_DFPRQX4 clk_r_REG913_S4 ( .D(n7413), .CP(net3007), .RN(n9555), .Q(
        n9346) );
  HS65_LH_DFPRQX4 clk_r_REG894_S4 ( .D(n7995), .CP(net3007), .RN(n2814), .Q(
        n8901) );
  HS65_LH_DFPRQX4 clk_r_REG727_S4 ( .D(n7929), .CP(net3007), .RN(n9557), .Q(
        n8996) );
  HS65_LH_DFPRQX4 clk_r_REG730_S4 ( .D(n8321), .CP(net3007), .RN(n9555), .Q(
        n9418) );
  HS65_LH_DFPRQX4 clk_r_REG890_S4 ( .D(n7990), .CP(net3007), .RN(n2814), .Q(
        n9090) );
  HS65_LH_DFPRQX4 clk_r_REG721_S4 ( .D(n7964), .CP(net3007), .RN(n9554), .Q(
        n9045) );
  HS65_LH_DFPRQX4 clk_r_REG741_S4 ( .D(n6114), .CP(net3007), .RN(n9557), .Q(
        n9065) );
  HS65_LH_DFPRQX4 clk_r_REG726_S4 ( .D(n7933), .CP(net3007), .RN(n9555), .Q(
        n8737) );
  HS65_LH_DFPRQX4 clk_r_REG739_S4 ( .D(n6121), .CP(net3007), .RN(n9554), .Q(
        n9062) );
  HS65_LH_DFPRQX4 clk_r_REG763_S4 ( .D(n7587), .CP(net3007), .RN(n9548), .Q(
        n9113) );
  HS65_LH_DFPRQX4 clk_r_REG718_S4 ( .D(n8019), .CP(net3007), .RN(n9557), .Q(
        n9040) );
  HS65_LH_DFPRQX4 clk_r_REG755_S4 ( .D(n6017), .CP(net3007), .RN(n9557), .Q(
        n8951) );
  HS65_LH_DFPRQX4 clk_r_REG864_S4 ( .D(n6264), .CP(net3007), .RN(n9557), .Q(
        n8950) );
  HS65_LH_DFPRQX4 clk_r_REG753_S4 ( .D(n6109), .CP(net3007), .RN(n9548), .Q(
        n8868) );
  HS65_LH_DFPRQX4 clk_r_REG862_S4 ( .D(n6529), .CP(net3007), .RN(n9557), .Q(
        n8949) );
  HS65_LH_DFPRQX4 clk_r_REG747_S4 ( .D(n6101), .CP(net3007), .RN(n9546), .Q(
        n9100) );
  HS65_LH_DFPRQX4 clk_r_REG759_S4 ( .D(n6100), .CP(net3007), .RN(n9551), .Q(
        n9098) );
  HS65_LH_DFPRQX4 clk_r_REG745_S4 ( .D(n6129), .CP(net3007), .RN(n9557), .Q(
        n9070) );
  HS65_LH_DFPRQX4 clk_r_REG761_S4 ( .D(n6119), .CP(net3007), .RN(n9545), .Q(
        n9102) );
  HS65_LH_DFPRQX4 clk_r_REG757_S4 ( .D(n6128), .CP(net3007), .RN(n9547), .Q(
        n9097) );
  HS65_LH_DFPRQX4 clk_r_REG742_S4 ( .D(n7517), .CP(net3007), .RN(n9547), .Q(
        n9245) );
  HS65_LH_DFPRQX4 clk_r_REG794_S4 ( .D(n6131), .CP(net3007), .RN(n9556), .Q(
        n9159) );
  HS65_LH_DFPRQX4 clk_r_REG786_S4 ( .D(n6027), .CP(net3007), .RN(n9551), .Q(
        n8866) );
  HS65_LH_DFPRQX4 clk_r_REG796_S4 ( .D(n2822), .CP(net3007), .RN(n9545), .Q(
        n9166) );
  HS65_LH_DFPRQX4 clk_r_REG781_S4 ( .D(n6133), .CP(net3007), .RN(n9555), .Q(
        n8861) );
  HS65_LH_DFPRQX4 clk_r_REG792_S4 ( .D(n6103), .CP(net3007), .RN(n9556), .Q(
        n9158) );
  HS65_LH_DFPRQX4 clk_r_REG740_S4 ( .D(n7501), .CP(net3007), .RN(n9547), .Q(
        n9247) );
  HS65_LH_DFPRQX4 clk_r_REG764_S4 ( .D(n7293), .CP(net3007), .RN(n9547), .Q(
        n9242) );
  HS65_LH_DFPRQX4 clk_r_REG756_S4 ( .D(n7571), .CP(net3007), .RN(n9546), .Q(
        n9203) );
  HS65_LH_DFPRQX4 clk_r_REG736_S4 ( .D(n7572), .CP(net3007), .RN(n9547), .Q(
        n9204) );
  HS65_LH_DFPRQX4 clk_r_REG866_S4 ( .D(n6333), .CP(net3007), .RN(n9545), .Q(
        n9162) );
  HS65_LH_DFPRQX4 clk_r_REG860_S4 ( .D(n6312), .CP(net3007), .RN(n9551), .Q(
        n8852) );
  HS65_LH_DFPRQX4 clk_r_REG733_S4 ( .D(n6132), .CP(net3007), .RN(n9551), .Q(
        n8862) );
  HS65_LH_DFPRQX4 clk_r_REG771_S4 ( .D(n6120), .CP(net3007), .RN(n9548), .Q(
        n9101) );
  HS65_LH_DFPRQX4 clk_r_REG769_S4 ( .D(n6102), .CP(net3007), .RN(n9545), .Q(
        n9096) );
  HS65_LH_DFPRQX4 clk_r_REG767_S4 ( .D(n6130), .CP(net3007), .RN(n9547), .Q(
        n9064) );
  HS65_LH_DFPRQX4 clk_r_REG765_S4 ( .D(n6014), .CP(net3007), .RN(n9546), .Q(
        n8947) );
  HS65_LH_DFPRQX4 clk_r_REG865_S4 ( .D(n6982), .CP(net3007), .RN(n9545), .Q(
        n9191) );
  HS65_LH_DFPRQX4 clk_r_REG789_S4 ( .D(n7569), .CP(net3007), .RN(n9547), .Q(
        n9205) );
  HS65_LH_DFPRQX4 clk_r_REG754_S4 ( .D(n7510), .CP(net3007), .RN(n9547), .Q(
        n9243) );
  HS65_LH_DFPRQX4 clk_r_REG848_S4 ( .D(n6345), .CP(net3007), .RN(n9555), .Q(
        n9010) );
  HS65_LH_DFPRQX4 clk_r_REG863_S4 ( .D(n6916), .CP(net3007), .RN(n9545), .Q(
        n9185) );
  HS65_LH_DFPRQX4 clk_r_REG748_S4 ( .D(n7278), .CP(net3007), .RN(n9546), .Q(
        n9200) );
  HS65_LH_DFPRQX4 clk_r_REG760_S4 ( .D(n7475), .CP(net3007), .RN(n9547), .Q(
        n9208) );
  HS65_LH_DFPRQX4 clk_r_REG746_S4 ( .D(n7580), .CP(net3007), .RN(n9548), .Q(
        n9254) );
  HS65_LH_DFPRQX4 clk_r_REG762_S4 ( .D(n7578), .CP(net3007), .RN(n9549), .Q(
        n9261) );
  HS65_LH_DFPRQX4 clk_r_REG758_S4 ( .D(n7585), .CP(net3007), .RN(n9548), .Q(
        n9257) );
  HS65_LH_DFPRQX4 clk_r_REG815_S4 ( .D(n6528), .CP(net3007), .RN(n9557), .Q(
        n8940) );
  HS65_LH_DFPRQX4 clk_r_REG840_S4 ( .D(n6272), .CP(net3007), .RN(n9548), .Q(
        n9067) );
  HS65_LH_DFPRQX4 clk_r_REG779_S4 ( .D(n6113), .CP(net3007), .RN(n9545), .Q(
        n9165) );
  HS65_LH_DFPRQX4 clk_r_REG842_S4 ( .D(n6278), .CP(net3007), .RN(n9545), .Q(
        n9164) );
  HS65_LH_DFPRQX4 clk_r_REG844_S4 ( .D(n6277), .CP(net3007), .RN(n9551), .Q(
        n8849) );
  HS65_LH_DFPRQX4 clk_r_REG811_S4 ( .D(n6265), .CP(net3007), .RN(n9554), .Q(
        n8855) );
  HS65_LH_DFPRQX4 clk_r_REG795_S4 ( .D(n7503), .CP(net3007), .RN(n9548), .Q(
        n9250) );
  HS65_LH_DFPRQX4 clk_r_REG787_S4 ( .D(n7594), .CP(net3007), .RN(n9546), .Q(
        n9201) );
  HS65_LH_DFPRQX4 clk_r_REG823_S4 ( .D(n6338), .CP(net3007), .RN(n9556), .Q(
        n9155) );
  HS65_LH_DFPRQX4 clk_r_REG817_S4 ( .D(n6986), .CP(net3007), .RN(n9556), .Q(
        n9154) );
  HS65_LH_DFPRQX4 clk_r_REG819_S4 ( .D(n6266), .CP(net3007), .RN(n9551), .Q(
        n8854) );
  HS65_LH_DFPRQX4 clk_r_REG850_S4 ( .D(n6346), .CP(net3007), .RN(n9556), .Q(
        n9160) );
  HS65_LH_DFPRQX4 clk_r_REG813_S4 ( .D(n6267), .CP(net3007), .RN(n9551), .Q(
        n8853) );
  HS65_LH_DFPRQX4 clk_r_REG825_S4 ( .D(n6985), .CP(net3007), .RN(n9556), .Q(
        n9156) );
  HS65_LH_DFPRQX4 clk_r_REG838_S4 ( .D(n6245), .CP(net3007), .RN(n9551), .Q(
        n8850) );
  HS65_LH_DFPRQX4 clk_r_REG793_S4 ( .D(n7279), .CP(net3007), .RN(n9546), .Q(
        n9198) );
  HS65_LH_DFPRQX4 clk_r_REG836_S4 ( .D(n6299), .CP(net3007), .RN(n9551), .Q(
        n8848) );
  HS65_LH_DFPRQX4 clk_r_REG867_S4 ( .D(n6984), .CP(net3007), .RN(n9545), .Q(
        n9188) );
  HS65_LH_DFPRQX4 clk_r_REG861_S4 ( .D(n6910), .CP(net3007), .RN(n9546), .Q(
        n9194) );
  HS65_LH_DFPRQX4 clk_r_REG772_S4 ( .D(n7577), .CP(net3007), .RN(n9549), .Q(
        n9263) );
  HS65_LH_DFPRQX4 clk_r_REG770_S4 ( .D(n7280), .CP(net3007), .RN(n9546), .Q(
        n9199) );
  HS65_LH_DFPRQX4 clk_r_REG768_S4 ( .D(n7579), .CP(net3007), .RN(n9547), .Q(
        n9244) );
  HS65_LH_DFPRQX4 clk_r_REG766_S4 ( .D(n7570), .CP(net3007), .RN(n9547), .Q(
        n9206) );
  HS65_LH_DFPRQX4 clk_r_REG734_S4 ( .D(n7502), .CP(net3007), .RN(n9549), .Q(
        n9265) );
  HS65_LH_DFPRQX4 clk_r_REG777_S4 ( .D(n6108), .CP(net3007), .RN(n9556), .Q(
        n9161) );
  HS65_LH_DFPRQX4 clk_r_REG849_S4 ( .D(n6999), .CP(net3007), .RN(n9549), .Q(
        n9260) );
  HS65_LH_DFPRQX4 clk_r_REG784_S4 ( .D(n5981), .CP(net3007), .RN(n9551), .Q(
        n8864) );
  HS65_LH_DFPRQX4 clk_r_REG751_S4 ( .D(n6026), .CP(net3007), .RN(n9554), .Q(
        n8867) );
  HS65_LH_DFPRQX4 clk_r_REG737_S4 ( .D(n6110), .CP(net3007), .RN(n9557), .Q(
        n9009) );
  HS65_LH_DFPRQX4 clk_r_REG773_S4 ( .D(n6127), .CP(net3007), .RN(n9556), .Q(
        n9152) );
  HS65_LH_DFPRQX4 clk_r_REG822_S4 ( .D(n6918), .CP(net3007), .RN(n9548), .Q(
        n9251) );
  HS65_LH_DFPRQX4 clk_r_REG790_S4 ( .D(n7588), .CP(net3007), .RN(n9545), .Q(
        n9095) );
  HS65_LH_DFPRQX4 clk_r_REG743_S4 ( .D(n6112), .CP(net3007), .RN(n9557), .Q(
        n9068) );
  HS65_LH_DFPRQX4 clk_r_REG816_S4 ( .D(n6917), .CP(net3007), .RN(n9548), .Q(
        n9249) );
  HS65_LH_DFPRQX4 clk_r_REG808_S4 ( .D(n2821), .CP(net3007), .RN(n9557), .Q(
        n8938) );
  HS65_LH_DFPRQX4 clk_r_REG841_S4 ( .D(n6993), .CP(net3007), .RN(n9549), .Q(
        n9262) );
  HS65_LH_DFPRQX4 clk_r_REG780_S4 ( .D(n7518), .CP(net3007), .RN(n9548), .Q(
        n9258) );
  HS65_LH_DFPRQX4 clk_r_REG843_S4 ( .D(n7000), .CP(net3007), .RN(n9549), .Q(
        n9267) );
  HS65_LH_DFPRQX4 clk_r_REG845_S4 ( .D(n6998), .CP(net3007), .RN(n9545), .Q(
        n9189) );
  HS65_LH_DFPRQX4 clk_r_REG831_S4 ( .D(n6259), .CP(net3007), .RN(n9556), .Q(
        n9116) );
  HS65_LH_DFPRQX4 clk_r_REG812_S4 ( .D(n2801), .CP(net3007), .RN(n9555), .Q(
        n9471) );
  HS65_LH_DFPRQX4 clk_r_REG824_S4 ( .D(n6991), .CP(net3007), .RN(n9545), .Q(
        n9186) );
  HS65_LH_DFPRQX4 clk_r_REG818_S4 ( .D(n6911), .CP(net3007), .RN(n9545), .Q(
        n9187) );
  HS65_LH_DFPRQX4 clk_r_REG820_S4 ( .D(n6983), .CP(net3007), .RN(n9545), .Q(
        n9190) );
  HS65_LH_DFPRQX4 clk_r_REG814_S4 ( .D(n6908), .CP(net3007), .RN(n9555), .Q(
        n9475) );
  HS65_LH_DFPRQX4 clk_r_REG851_S4 ( .D(n7001), .CP(net3007), .RN(n9555), .Q(
        n9470) );
  HS65_LH_DFPRQX4 clk_r_REG839_S4 ( .D(n6992), .CP(net3007), .RN(n9549), .Q(
        n9264) );
  HS65_LH_DFPRQX4 clk_r_REG837_S4 ( .D(n7002), .CP(net3007), .RN(n9546), .Q(
        n9193) );
  HS65_LH_DFPRQX4 clk_r_REG826_S4 ( .D(n6909), .CP(net3007), .RN(n9555), .Q(
        n9469) );
  HS65_LH_DFPRQX4 clk_r_REG749_S4 ( .D(n5980), .CP(net3007), .RN(n9545), .Q(
        n8865) );
  HS65_LH_DFPRQX4 clk_r_REG806_S4 ( .D(n6340), .CP(net3007), .RN(n9546), .Q(
        n8937) );
  HS65_LH_DFPRQX4 clk_r_REG775_S4 ( .D(n6111), .CP(net3007), .RN(n9556), .Q(
        n9153) );
  HS65_LH_DFPRQX4 clk_r_REG774_S4 ( .D(n7586), .CP(net3007), .RN(n9550), .Q(
        n9363) );
  HS65_LH_DFPRQX4 clk_r_REG778_S4 ( .D(n7509), .CP(net3007), .RN(n9547), .Q(
        n9207) );
  HS65_LH_DFPRQX4 clk_r_REG785_S4 ( .D(n7595), .CP(net3007), .RN(n9548), .Q(
        n9256) );
  HS65_LH_DFPRQX4 clk_r_REG752_S4 ( .D(n7593), .CP(net3007), .RN(n9546), .Q(
        n9202) );
  HS65_LH_DFPRQX4 clk_r_REG738_S4 ( .D(n7555), .CP(net3007), .RN(n9546), .Q(
        n9197) );
  HS65_LH_DFPRQX4 clk_r_REG791_S4 ( .D(n7508), .CP(net3007), .RN(n9549), .Q(
        n9266) );
  HS65_LH_DFPRQX4 clk_r_REG744_S4 ( .D(n7515), .CP(net3007), .RN(n9548), .Q(
        n9253) );
  HS65_LH_DFPRQX4 clk_r_REG803_S4 ( .D(n6339), .CP(net3007), .RN(n9551), .Q(
        n8851) );
  HS65_LH_DFPRQX4 clk_r_REG833_S4 ( .D(n6258), .CP(net3007), .RN(n9556), .Q(
        n9157) );
  HS65_LH_DFPRQX4 clk_r_REG829_S4 ( .D(n6497), .CP(net3007), .RN(n9547), .Q(
        n8860) );
  HS65_LH_DFPRQX4 clk_r_REG827_S4 ( .D(n6498), .CP(net3007), .RN(n9547), .Q(
        n8859) );
  HS65_LH_DFPRQX4 clk_r_REG856_S4 ( .D(n6975), .CP(net3007), .RN(n9547), .Q(
        n8858) );
  HS65_LH_DFPRQX4 clk_r_REG852_S4 ( .D(n6976), .CP(net3007), .RN(n9548), .Q(
        n8856) );
  HS65_LH_DFPRQX4 clk_r_REG832_S4 ( .D(n6972), .CP(net3007), .RN(n9546), .Q(
        n9195) );
  HS65_LH_DFPRQX4 clk_r_REG809_S4 ( .D(n6348), .CP(net3007), .RN(n9545), .Q(
        n9163) );
  HS65_LH_DFPRQX4 clk_r_REG750_S4 ( .D(n7560), .CP(net3007), .RN(n9548), .Q(
        n9259) );
  HS65_LH_DFPRQX4 clk_r_REG805_S4 ( .D(n6895), .CP(net3007), .RN(n9548), .Q(
        n9248) );
  HS65_LH_DFPRQX4 clk_r_REG807_S4 ( .D(n6890), .CP(net3007), .RN(n9547), .Q(
        n9246) );
  HS65_LH_DFPRQX4 clk_r_REG776_S4 ( .D(n7516), .CP(net3007), .RN(n9550), .Q(
        n9364) );
  HS65_LH_DFPRQX4 clk_r_REG834_S4 ( .D(n6724), .CP(net3007), .RN(n9546), .Q(
        n9192) );
  HS65_LH_DFPRQX4 clk_r_REG830_S4 ( .D(n6457), .CP(net3007), .RN(n9546), .Q(
        n9196) );
  HS65_LH_DFPRQX4 clk_r_REG828_S4 ( .D(n6973), .CP(net3007), .RN(n9548), .Q(
        n9255) );
  HS65_LH_DFPRQX4 clk_r_REG855_S4 ( .D(n6974), .CP(net3007), .RN(n9555), .Q(
        n9468) );
  HS65_LH_DFPRQX4 clk_r_REG853_S4 ( .D(n6726), .CP(net3007), .RN(n9555), .Q(
        n9474) );
  HS65_LH_DFPRQX4 clk_r_REG810_S4 ( .D(n6943), .CP(net3007), .RN(n9547), .Q(
        n9240) );
  HS65_LH_DFPRQX4 clk_r_REG594_S4 ( .D(n7992), .CP(net3007), .RN(n9550), .Q(
        n8766) );
  HS65_LH_DFPRQX4 clk_r_REG596_S4 ( .D(n7958), .CP(net3007), .RN(n9555), .Q(
        n8603) );
  HS65_LH_DFPRQX4 clk_r_REG615_S4 ( .D(n8038), .CP(net3007), .RN(n9549), .Q(
        n9318) );
  HS65_LL_DFPQX4 clk_r_REG640_S5 ( .D(\u_DataPath/u_idexreg/N10 ), .CP(clk), 
        .Q(n8732) );
  HS65_LL_DFPQX4 clk_r_REG576_S2 ( .D(n8306), .CP(clk), .Q(n8767) );
  HS65_LH_DFPQX4 clk_r_REG289_S2 ( .D(n5632), .CP(clk), .Q(n9005) );
  HS65_LH_DFPQX9 clk_r_REG634_S6 ( .D(write_byte_snps_wire), .CP(clk), .Q(
        n8874) );
  HS65_LH_DFPQX9 clk_r_REG111_S4 ( .D(addr_to_iram_29), .CP(net3007), .Q(n8562) );
  HS65_LH_DFPQX9 clk_r_REG204_S5 ( .D(addr_to_iram_28), .CP(net3007), .Q(n8561) );
  HS65_LH_DFPQX9 clk_r_REG197_S5 ( .D(addr_to_iram_27), .CP(net3007), .Q(n8560) );
  HS65_LH_DFPQX9 clk_r_REG190_S5 ( .D(addr_to_iram_26), .CP(net3007), .Q(n8559) );
  HS65_LH_DFPQX9 clk_r_REG145_S3 ( .D(addr_to_iram_15), .CP(net3007), .Q(n8558) );
  HS65_LH_DFPQX9 clk_r_REG183_S5 ( .D(addr_to_iram_25), .CP(net3007), .Q(n8557) );
  HS65_LH_DFPQX18 clk_r_REG244_S5 ( .D(addr_to_iram_21), .CP(net3007), .Q(
        n8556) );
  HS65_LH_DFPQX18 clk_r_REG160_S2 ( .D(addr_to_iram_19), .CP(net3007), .Q(
        n8555) );
  HS65_LH_DFPQX9 clk_r_REG324_S5 ( .D(addr_to_iram_14), .CP(net3007), .Q(n8554) );
  HS65_LH_DFPQX9 clk_r_REG177_S5 ( .D(addr_to_iram_24), .CP(net3007), .Q(n8552) );
  HS65_LH_DFPQX18 clk_r_REG167_S5 ( .D(addr_to_iram_20), .CP(net3007), .Q(
        n8551) );
  HS65_LH_DFPQX18 clk_r_REG49_S4 ( .D(addr_to_iram_18), .CP(net3007), .Q(n8550) );
  HS65_LH_DFPQX18 clk_r_REG420_S4 ( .D(addr_to_iram_1), .CP(net3007), .Q(n8549) );
  HS65_LH_DFPQX18 clk_r_REG88_S4 ( .D(addr_to_iram_0), .CP(net3007), .Q(n8548)
         );
  HS65_LH_DFPQX18 clk_r_REG463_S4 ( .D(addr_to_iram_2), .CP(net3007), .Q(n8545) );
  HS65_LH_DFPQX18 clk_r_REG452_S4 ( .D(addr_to_iram_3), .CP(net3007), .Q(n8544) );
  HS65_LH_DFPQX18 clk_r_REG428_S4 ( .D(addr_to_iram_4), .CP(net3007), .Q(n8543) );
  HS65_LH_DFPQX18 clk_r_REG35_S4 ( .D(addr_to_iram_5), .CP(net3007), .Q(n8542)
         );
  HS65_LH_DFPQX18 clk_r_REG312_S4 ( .D(addr_to_iram_8), .CP(net3007), .Q(n8541) );
  HS65_LH_DFPQX18 clk_r_REG302_S4 ( .D(addr_to_iram_6), .CP(net3007), .Q(n8540) );
  HS65_LH_DFPQX18 clk_r_REG317_S4 ( .D(addr_to_iram_10), .CP(net3007), .Q(
        n8539) );
  HS65_LH_DFPQX9 clk_r_REG15_S5 ( .D(addr_to_iram_23), .CP(net3007), .Q(n8538)
         );
  HS65_LH_DFPQX18 clk_r_REG369_S4 ( .D(addr_to_iram_9), .CP(net3007), .Q(n8537) );
  HS65_LH_DFPQX9 clk_r_REG308_S4 ( .D(addr_to_iram_7), .CP(net3007), .Q(n8536)
         );
  HS65_LH_DFPQX18 clk_r_REG279_S2 ( .D(addr_to_iram_16), .CP(net3007), .Q(
        n8535) );
  HS65_LH_DFPQX9 clk_r_REG327_S5 ( .D(addr_to_iram_12), .CP(net3007), .Q(n8534) );
  HS65_LH_DFPQX9 clk_r_REG42_S4 ( .D(addr_to_iram_13), .CP(net3007), .Q(n8533)
         );
  HS65_LH_DFPQX9 clk_r_REG175_S5 ( .D(addr_to_iram_22), .CP(net3007), .Q(n8531) );
  HS65_LH_DFPQX18 clk_r_REG153_S2 ( .D(addr_to_iram_17), .CP(net3007), .Q(
        n8530) );
  HS65_LH_DFPQX4 clk_r_REG311_S1 ( .D(\u_DataPath/branch_target_i [10]), .CP(
        clk), .Q(n9449) );
  HS65_LH_DFPQX4 clk_r_REG469_S2 ( .D(n5654), .CP(clk), .Q(n9414) );
  HS65_LH_DFPQX4 clk_r_REG275_S2 ( .D(n5829), .CP(clk), .Q(n9396) );
  HS65_LH_DFPQX4 clk_r_REG48_S3 ( .D(\u_DataPath/jump_address_i [20]), .CP(clk), .Q(n9377) );
  HS65_LH_DFPQX4 clk_r_REG398_S3 ( .D(n3025), .CP(clk), .Q(n9336) );
  HS65_LH_DFPQX4 clk_r_REG661_S7 ( .D(n7309), .CP(clk), .Q(n9316) );
  HS65_LH_DFPQX4 clk_r_REG496_S3 ( .D(n2926), .CP(clk), .Q(n9294) );
  HS65_LH_DFPQX4 clk_r_REG535_S2 ( .D(n5620), .CP(clk), .Q(n9274) );
  HS65_LH_DFPQX4 clk_r_REG695_S1 ( .D(n8027), .CP(clk), .Q(n9230) );
  HS65_LH_DFPQX4 clk_r_REG691_S1 ( .D(n7976), .CP(clk), .Q(n9211) );
  HS65_LH_DFPQX4 clk_r_REG711_S1 ( .D(\u_DataPath/cw_to_ex_i [19]), .CP(clk), 
        .Q(n9142) );
  HS65_LH_DFPQX4 clk_r_REG60_S4 ( .D(n7655), .CP(clk), .Q(n9124) );
  HS65_LH_DFPQX4 clk_r_REG333_S2 ( .D(n5580), .CP(clk), .Q(n9091) );
  HS65_LH_DFPQX4 clk_r_REG423_S2 ( .D(\u_DataPath/u_execute/link_value_i [5]), 
        .CP(clk), .Q(n9073) );
  HS65_LH_DFPQX4 clk_r_REG374_S2 ( .D(n5540), .CP(clk), .Q(n9038) );
  HS65_LH_DFPQX4 clk_r_REG395_S3 ( .D(n8338), .CP(clk), .Q(n9023) );
  HS65_LH_DFPQX4 clk_r_REG461_S2 ( .D(n5909), .CP(clk), .Q(n9006) );
  HS65_LH_DFPQX4 clk_r_REG218_S2 ( .D(n5929), .CP(clk), .Q(n8986) );
  HS65_LH_DFPQX4 clk_r_REG441_S2 ( .D(n5700), .CP(clk), .Q(n8971) );
  HS65_LH_DFPQX4 clk_r_REG10_S4 ( .D(\u_DataPath/pc_4_i [25]), .CP(net3007), 
        .Q(n8955) );
  HS65_LH_DFPQX4 clk_r_REG271_S2 ( .D(n5637), .CP(clk), .Q(n8927) );
  HS65_LH_DFPQX4 clk_r_REG315_S2 ( .D(n5791), .CP(clk), .Q(n8912) );
  HS65_LH_DFPQX4 clk_r_REG194_S2 ( .D(n5672), .CP(clk), .Q(n8893) );
  HS65_LH_DFPQX4 clk_r_REG570_S2 ( .D(\u_DataPath/toPC2_i [0]), .CP(clk), .Q(
        n8872) );
  HS65_LH_DFPQX4 clk_r_REG443_S1 ( .D(\u_DataPath/branch_target_i [6]), .CP(
        clk), .Q(n8829) );
  HS65_LH_DFPQX4 clk_r_REG106_S1 ( .D(n8040), .CP(clk), .Q(n8774) );
  HS65_LH_DFPQX4 clk_r_REG21_S1 ( .D(n7659), .CP(clk), .Q(n8741) );
  HS65_LH_DFPQX4 clk_r_REG58_S1 ( .D(n8445), .CP(clk), .Q(n8721) );
  HS65_LH_DFPQX4 clk_r_REG490_S1 ( .D(\u_DataPath/mem_writedata_out_i [2]), 
        .CP(clk), .Q(n8704) );
  HS65_LH_DFPQX4 clk_r_REG123_S3 ( .D(\u_DataPath/data_read_ex_1_i [27]), .CP(
        clk), .Q(n8672) );
  HS65_LH_DFPQX4 clk_r_REG108_S2 ( .D(\u_DataPath/data_read_ex_2_i [31]), .CP(
        clk), .Q(n8657) );
  HS65_LH_DFPQX4 clk_r_REG499_S2 ( .D(\u_DataPath/data_read_ex_1_i [30]), .CP(
        clk), .Q(n8641) );
  HS65_LH_DFPQX4 clk_r_REG70_S3 ( .D(\u_DataPath/data_read_ex_1_i [14]), .CP(
        clk), .Q(n8626) );
  HS65_LH_DFPQX4 clk_r_REG381_S3 ( .D(\u_DataPath/jump_address_i [9]), .CP(clk), .Q(n8611) );
  HS65_LH_DFPQX4 clk_r_REG265_S3 ( .D(n8290), .CP(clk), .Q(n8593) );
  HS65_LH_DFPQX4 clk_r_REG694_S1 ( .D(n7997), .CP(clk), .Q(n8569) );
  HS65_LH_IVX2 U9389 ( .A(Data_out_fromRAM[19]), .Z(n8197) );
  HS65_LH_IVX2 U9392 ( .A(Data_out_fromRAM[22]), .Z(n8284) );
  HS65_LH_IVX4 U4668 ( .A(Data_out_fromRAM[28]), .Z(n8294) );
  HS65_LHS_XNOR2X6 U4150 ( .A(n9337), .B(n9148), .Z(
        \u_DataPath/u_execute/link_value_i [8]) );
  HS65_LH_IVX9 U6534 ( .A(n8675), .Z(\u_DataPath/jump_address_i [6]) );
  HS65_LL_AOI13X4 U5065 ( .A(n8899), .B(n9151), .C(n8925), .D(n8941), .Z(n2989) );
  HS65_LH_IVX9 U6589 ( .A(n8606), .Z(\u_DataPath/jump_address_i [5]) );
  HS65_LL_AO31X18 U4142 ( .A(n8945), .B(n9094), .C(n9114), .D(n3107), .Z(n3149) );
  HS65_LH_NAND2X2 U5036 ( .A(n2989), .B(n9103), .Z(n2949) );
  HS65_LL_OR2X9 U3576 ( .A(n8760), .B(n3107), .Z(n3236) );
  HS65_LHS_XNOR2X3 U6722 ( .A(n9224), .B(n7443), .Z(
        \u_DataPath/u_execute/link_value_i [19]) );
  HS65_LH_NOR2X5 U4141 ( .A(n9380), .B(n7428), .Z(n7429) );
  HS65_LHS_XOR2X3 U4138 ( .A(n9333), .B(n7629), .Z(
        \u_DataPath/u_execute/link_value_i [12]) );
  HS65_LH_IVX4 U5146 ( .A(\u_DataPath/dataOut_exe_i [27]), .Z(n3104) );
  HS65_LH_IVX4 U4190 ( .A(n5633), .Z(n5634) );
  HS65_LH_NAND2X5 U4582 ( .A(n8976), .B(n5820), .Z(n5752) );
  HS65_LHS_XNOR2X6 U7592 ( .A(n9466), .B(n9046), .Z(n7200) );
  HS65_LHS_XNOR2X3 U7447 ( .A(n8813), .B(n9092), .Z(n6491) );
  HS65_LH_OR2X4 U7320 ( .A(\u_DataPath/dataOut_exe_i [13]), .B(n9012), .Z(
        n3063) );
  HS65_LHS_XNOR2X6 U7584 ( .A(n9467), .B(n9339), .Z(n7197) );
  HS65_LH_OAI12X3 U5941 ( .A(n9003), .B(n5573), .C(n8716), .Z(n5545) );
  HS65_LH_NAND2X4 U6769 ( .A(n8679), .B(n2800), .Z(n8413) );
  HS65_LHS_XNOR2X6 U6832 ( .A(n9462), .B(n8906), .Z(n7198) );
  HS65_LH_OR2X4 U5887 ( .A(\u_DataPath/dataOut_exe_i [15]), .B(n9012), .Z(
        n2840) );
  HS65_LL_OAI12X2 U6766 ( .A(n9055), .B(n5646), .C(n8775), .Z(n5572) );
  HS65_LH_NAND2X4 U5879 ( .A(n3017), .B(n2800), .Z(n8402) );
  HS65_LHS_XNOR2X6 U7595 ( .A(n8810), .B(n9112), .Z(n7199) );
  HS65_LHS_XOR2X6 U8450 ( .A(n9217), .B(n7625), .Z(
        \u_DataPath/u_execute/link_value_i [11]) );
  HS65_LHS_XOR2X6 U7509 ( .A(n8811), .B(n8906), .Z(n7203) );
  HS65_LL_NOR2X3 U5921 ( .A(n7206), .B(n7205), .Z(n7207) );
  HS65_LH_AOI12X2 U3451 ( .A(n9109), .B(n5705), .C(n8710), .Z(n5699) );
  HS65_LH_NAND2X7 U5923 ( .A(n7198), .B(n7197), .Z(n7214) );
  HS65_LH_NOR2X6 U4285 ( .A(\u_DataPath/dataOut_exe_i [1]), .B(
        \u_DataPath/dataOut_exe_i [0]), .Z(n3564) );
  HS65_LL_NOR2X3 U4540 ( .A(n9292), .B(n7627), .Z(n6758) );
  HS65_LH_NAND2X5 U4167 ( .A(n9175), .B(n6487), .Z(n6495) );
  HS65_LH_NOR2X6 U4594 ( .A(n7203), .B(n7202), .Z(n7208) );
  HS65_LL_NAND3X3 U6790 ( .A(n7201), .B(n7200), .C(n7199), .Z(n7213) );
  HS65_LH_NOR2X3 U4135 ( .A(\u_DataPath/dataOut_exe_i [0]), .B(n3178), .Z(
        n2954) );
  HS65_LH_IVX7 U4665 ( .A(\u_DataPath/dataOut_exe_i [0]), .Z(n8156) );
  HS65_LH_AOI12X2 U4567 ( .A(n9302), .B(n5705), .C(n9414), .Z(n5655) );
  HS65_LH_IVX4 U7415 ( .A(n8263), .Z(n2938) );
  HS65_LH_NOR2X5 U5815 ( .A(\u_DataPath/dataOut_exe_i [21]), .B(n3178), .Z(
        n3179) );
  HS65_LL_NOR2X2 U6734 ( .A(\u_DataPath/dataOut_exe_i [18]), .B(n3178), .Z(
        n3153) );
  HS65_LH_NOR2X5 U4557 ( .A(\u_DataPath/dataOut_exe_i [31]), .B(n3980), .Z(
        n8452) );
  HS65_LH_NOR2X5 U4554 ( .A(\u_DataPath/dataOut_exe_i [22]), .B(n3980), .Z(
        n8438) );
  HS65_LH_NOR2X5 U5023 ( .A(\u_DataPath/dataOut_exe_i [29]), .B(n3178), .Z(
        n3121) );
  HS65_LH_NOR2X5 U5030 ( .A(\u_DataPath/dataOut_exe_i [30]), .B(n3178), .Z(
        n2886) );
  HS65_LH_NOR2X5 U5812 ( .A(\u_DataPath/dataOut_exe_i [28]), .B(n3178), .Z(
        n3116) );
  HS65_LH_IVX7 U5829 ( .A(n3056), .Z(n8406) );
  HS65_LL_OAI21X3 U5878 ( .A(n8727), .B(n9115), .C(n3565), .Z(n2813) );
  HS65_LH_NAND2X5 U4899 ( .A(n9287), .B(n2797), .Z(n8404) );
  HS65_LH_IVX7 U4131 ( .A(n3009), .Z(n8405) );
  HS65_LH_IVX4 U7583 ( .A(n8158), .Z(n2943) );
  HS65_LH_OAI21X3 U6771 ( .A(n8727), .B(n9115), .C(n3565), .Z(n8457) );
  HS65_LH_NAND2AX7 U4134 ( .A(n8709), .B(n2712), .Z(n3023) );
  HS65_LH_NAND2X7 U4122 ( .A(n3109), .B(n2712), .Z(n3110) );
  HS65_LH_AOI21X2 U5014 ( .A(n7654), .B(n2710), .C(n2886), .Z(n2891) );
  HS65_LH_IVX7 U4196 ( .A(n8159), .Z(n8376) );
  HS65_LH_NAND2X5 U5579 ( .A(n9283), .B(n2797), .Z(n8412) );
  HS65_LH_OAI21X3 U6702 ( .A(n8656), .B(n3149), .C(n3063), .Z(n3064) );
  HS65_LL_NAND2X2 U5808 ( .A(n8278), .B(n2798), .Z(n3216) );
  HS65_LH_NAND2X4 U5799 ( .A(n3090), .B(n8406), .Z(n3060) );
  HS65_LHS_XNOR2X6 U3705 ( .A(n8924), .B(n5693), .Z(\u_DataPath/toPC2_i [9])
         );
  HS65_LL_NAND2X2 U4217 ( .A(n3184), .B(n8730), .Z(n3186) );
  HS65_LH_NOR2X5 U6677 ( .A(n8637), .B(n3181), .Z(n3166) );
  HS65_LL_NAND2X7 U7296 ( .A(n7302), .B(n6496), .Z(n6861) );
  HS65_LH_IVX2 U8197 ( .A(n5328), .Z(n4927) );
  HS65_LH_NAND2AX7 U4125 ( .A(n8680), .B(n2778), .Z(n3150) );
  HS65_LL_AOI112X4 U4528 ( .A(n8694), .B(n2712), .C(n3127), .D(n3126), .Z(
        n3128) );
  HS65_LH_AOI22X6 U4538 ( .A(n2710), .B(n8717), .C(n9331), .D(n2778), .Z(n3146) );
  HS65_LL_AO112X4 U3750 ( .A(n8278), .B(n2712), .C(n2954), .D(n2953), .Z(n2774) );
  HS65_LH_NOR2X5 U5773 ( .A(n8632), .B(n3181), .Z(n3171) );
  HS65_LH_OAI21X3 U3548 ( .A(n3983), .B(n2772), .C(n3982), .Z(n3984) );
  HS65_LH_AOI12X2 U4547 ( .A(n5820), .B(n5884), .C(n5819), .Z(n5821) );
  HS65_LH_AOI22X3 U5015 ( .A(n3104), .B(n2800), .C(n8696), .D(n2798), .Z(n3105) );
  HS65_LL_AOI12X2 U5825 ( .A(n3090), .B(n8444), .C(n3089), .Z(n3093) );
  HS65_LH_NAND2AX7 U5025 ( .A(n8634), .B(n2778), .Z(n2935) );
  HS65_LH_AOI22X6 U5007 ( .A(n2710), .B(n8697), .C(n9340), .D(n2778), .Z(n3097) );
  HS65_LL_NAND2X2 U5115 ( .A(n3184), .B(n9435), .Z(n3069) );
  HS65_LH_AOI12X2 U5029 ( .A(n5613), .B(n5682), .C(n5612), .Z(n5614) );
  HS65_LL_IVX13 U5009 ( .A(n2798), .Z(n2794) );
  HS65_LHS_XNOR2X3 U6711 ( .A(n9000), .B(n5884), .Z(
        \u_DataPath/u_execute/resAdd1_i [16]) );
  HS65_LH_AOI12X2 U3441 ( .A(n9150), .B(n5884), .C(n8715), .Z(n5878) );
  HS65_LH_AOI22X1 U5789 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][7] ), .B(n9208), 
        .C(n9100), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][7] ), .Z(n6043)
         );
  HS65_LH_AOI22X1 U5787 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][7] ), .B(n9196), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][7] ), .D(
        n9192), .Z(n6461) );
  HS65_LL_OAI21X2 U3781 ( .A(n8649), .B(n2772), .C(n3105), .Z(n8448) );
  HS65_LL_NAND3X2 U5810 ( .A(n3090), .B(n8383), .C(n8382), .Z(n2951) );
  HS65_LL_OAI112X3 U4465 ( .A(n2794), .B(n3100), .C(n3099), .D(n2843), .Z(
        n7676) );
  HS65_LL_NOR2X5 U6613 ( .A(n3088), .B(n3087), .Z(\lte_x_57/B[25] ) );
  HS65_LL_IVX7 U4939 ( .A(n3138), .Z(\sub_x_51/A[16] ) );
  HS65_LL_NAND2X2 U5072 ( .A(n9229), .B(n2976), .Z(n2977) );
  HS65_LL_OAI21X2 U3749 ( .A(n8648), .B(n2772), .C(n3125), .Z(n2773) );
  HS65_LL_NAND2X4 U6614 ( .A(n3182), .B(n2826), .Z(n4918) );
  HS65_LH_IVX2 U7492 ( .A(n5365), .Z(n5173) );
  HS65_LH_NAND3X2 U7488 ( .A(\u_DataPath/cw_to_ex_i [1]), .B(n4019), .C(n5327), 
        .Z(n4020) );
  HS65_LL_NOR2X6 U5113 ( .A(n2862), .B(n3245), .Z(n4774) );
  HS65_LL_IVX7 U4530 ( .A(n3950), .Z(\sub_x_51/A[5] ) );
  HS65_LH_AOI12X2 U3442 ( .A(n9391), .B(n5872), .C(n9276), .Z(n5782) );
  HS65_LH_IVX9 U5126 ( .A(n3301), .Z(n5161) );
  HS65_LH_AOI22X1 U4946 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][17] ), .B(n9162), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][17] ), .D(
        n9190), .Z(n6363) );
  HS65_LH_AOI22X1 U5737 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][11] ), .B(n9199), 
        .C(n9198), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][11] ), .Z(n6803)
         );
  HS65_LH_AOI22X1 U5748 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][17] ), .B(n9196), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][17] ), .D(
        n9192), .Z(n6360) );
  HS65_LH_AOI22X1 U5705 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][17] ), .B(n9208), 
        .C(n9100), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][17] ), .Z(n5943)
         );
  HS65_LL_IVX7 U4462 ( .A(n3588), .Z(n3241) );
  HS65_LH_AOI22X1 U5738 ( .A(n9207), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][16] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][16] ), .D(n9266), 
        .Z(n6067) );
  HS65_LH_AOI22X1 U6635 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][24] ), .B(n9162), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][24] ), .D(
        n9190), .Z(n6270) );
  HS65_LH_AOI22X1 U6633 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][24] ), .B(n9196), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][24] ), .D(
        n9192), .Z(n6263) );
  HS65_LH_AOI22X1 U7265 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][22] ), .B(n9162), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][22] ), .D(
        n8854), .Z(n6549) );
  HS65_LH_AOI22X1 U6640 ( .A(n9207), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][24] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][24] ), .D(n9266), 
        .Z(n5979) );
  HS65_LH_AOI22X1 U5659 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][23] ), .B(n9208), 
        .C(n9100), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][23] ), .Z(n7119)
         );
  HS65_LH_AOI22X1 U6657 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][23] ), .B(n9196), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][23] ), .D(
        n9192), .Z(n6332) );
  HS65_LH_NAND2X4 U5537 ( .A(n3239), .B(n7321), .Z(n4680) );
  HS65_LH_AOI22X1 U5709 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][18] ), .B(n9208), 
        .C(n9100), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][18] ), .Z(n7221)
         );
  HS65_LH_NAND2X7 U8167 ( .A(\sub_x_51/A[13] ), .B(n2786), .Z(n5232) );
  HS65_LHS_XOR2X3 U7159 ( .A(n5311), .B(n5312), .Z(n4964) );
  HS65_LH_AOI22X1 U6641 ( .A(n9207), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][18] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][18] ), .D(n9266), 
        .Z(n7225) );
  HS65_LH_AOI22X1 U5651 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][19] ), .B(n9208), 
        .C(n9100), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][19] ), .Z(n6764)
         );
  HS65_LH_AOI22X3 U4508 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][31] ), .B(n9247), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][31] ), .D(
        n9227), .Z(n7507) );
  HS65_LH_AOI22X1 U7246 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][30] ), .B(n9162), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][30] ), .D(
        n8854), .Z(n6569) );
  HS65_LHS_XOR2X3 U4501 ( .A(n9047), .B(n5782), .Z(
        \u_DataPath/u_execute/resAdd1_i [15]) );
  HS65_LH_AOI22X1 U4524 ( .A(n9207), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][20] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][20] ), .D(n9095), 
        .Z(n7103) );
  HS65_LH_AOI22X1 U4525 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][20] ), .B(n9208), 
        .C(n9100), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][20] ), .Z(n7099)
         );
  HS65_LH_AOI22X1 U4497 ( .A(n9201), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][30] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][30] ), .D(n9202), 
        .Z(n7540) );
  HS65_LH_AOI22X1 U5677 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][15] ), .B(n9199), 
        .C(n9198), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][15] ), .Z(n7260)
         );
  HS65_LH_AOI22X1 U7247 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][28] ), .B(n9162), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][28] ), .D(
        n8854), .Z(n6526) );
  HS65_LH_AOI22X1 U5698 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][10] ), .B(n9208), 
        .C(n9100), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][10] ), .Z(n7039)
         );
  HS65_LH_AOI22X1 U6659 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][13] ), .B(n9208), 
        .C(n9100), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][13] ), .Z(n7019)
         );
  HS65_LH_AOI22X1 U6655 ( .A(n9207), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][13] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][13] ), .D(n9266), 
        .Z(n7023) );
  HS65_LH_AOI22X1 U5722 ( .A(n9207), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][10] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][10] ), .D(n9266), 
        .Z(n7043) );
  HS65_LH_AOI22X1 U6672 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][12] ), .B(n9199), 
        .C(n9198), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][12] ), .Z(n7138)
         );
  HS65_LH_AOI22X1 U4977 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][13] ), .B(n9162), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][13] ), .D(
        n9190), .Z(n6403) );
  HS65_LH_AOI22X1 U4959 ( .A(n9161), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][8] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][8] ), .D(n9266), 
        .Z(n6848) );
  HS65_LH_AOI22X1 U6670 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][19] ), .B(n9196), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][19] ), .D(
        n9192), .Z(n6290) );
  HS65_LH_NOR2X5 U5420 ( .A(\lte_x_57/B[10] ), .B(n5386), .Z(n3676) );
  HS65_LH_AOI22X1 U5694 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][13] ), .B(n9196), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][13] ), .D(
        n9192), .Z(n6400) );
  HS65_LL_NOR2X3 U5561 ( .A(n4901), .B(n4902), .Z(n5454) );
  HS65_LH_AOI22X1 U4932 ( .A(n9201), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][28] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][28] ), .D(n9202), 
        .Z(n7597) );
  HS65_LH_AOI22X1 U6649 ( .A(n9207), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][25] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][25] ), .D(n9266), 
        .Z(n7483) );
  HS65_LH_AOI22X1 U5623 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][8] ), .B(n9199), 
        .C(n9198), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][8] ), .Z(n6843)
         );
  HS65_LH_AOI22X1 U4961 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][16] ), .B(n9196), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][16] ), .D(
        n9157), .Z(n6168) );
  HS65_LL_NOR2X2 U6545 ( .A(\lte_x_57/B[7] ), .B(n4346), .Z(n4336) );
  HS65_LH_AOI22X1 U5724 ( .A(n9201), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][31] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][31] ), .D(n9202), 
        .Z(n7520) );
  HS65_LH_AOI22X1 U5666 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][21] ), .B(n9196), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][21] ), .D(
        n9192), .Z(n6380) );
  HS65_LH_AOI22X1 U6651 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][25] ), .B(n9208), 
        .C(n9100), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][25] ), .Z(n7479)
         );
  HS65_LH_AOI22X1 U4953 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][21] ), .B(n9162), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][21] ), .D(
        n9190), .Z(n6383) );
  HS65_LH_AOI22X1 U6625 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][22] ), .B(n9199), 
        .C(n9198), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][22] ), .Z(n7178)
         );
  HS65_LH_AOI22X1 U5617 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][26] ), .B(n9199), 
        .C(n9198), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][26] ), .Z(n6783)
         );
  HS65_LH_AOI22X1 U6664 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][27] ), .B(n9196), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][27] ), .D(
        n9192), .Z(n6311) );
  HS65_LH_AOI22X1 U5649 ( .A(n9207), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][14] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][14] ), .D(n9266), 
        .Z(n6087) );
  HS65_LH_AOI22X1 U4976 ( .A(n9161), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][6] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][6] ), .D(n9266), 
        .Z(n6828) );
  HS65_LH_AOI22X3 U8092 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][0] ), .B(n9098), 
        .C(n9200), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][0] ), .Z(n7284)
         );
  HS65_LH_AOI22X1 U5001 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][2] ), .B(n9196), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][2] ), .D(
        n9157), .Z(n6220) );
  HS65_LH_AOI22X1 U4929 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][0] ), .B(n9196), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][0] ), .D(
        n9157), .Z(n6200) );
  HS65_LH_AOI22X1 U5780 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][4] ), .B(n9196), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][4] ), .D(
        n9192), .Z(n6420) );
  HS65_LH_AOI22X1 U6647 ( .A(n9207), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][1] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][1] ), .D(n9266), 
        .Z(n7245) );
  HS65_LH_AOI22X1 U5753 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][1] ), .B(n9208), 
        .C(n9100), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][1] ), .Z(n7241)
         );
  HS65_LH_IVX2 U8116 ( .A(n5356), .Z(n5384) );
  HS65_LH_IVX2 U7094 ( .A(n5455), .Z(n4006) );
  HS65_LH_NOR2X5 U6576 ( .A(n4203), .B(n3338), .Z(n3861) );
  HS65_LL_OAI12X2 U6419 ( .A(n5284), .B(n4998), .C(n5303), .Z(n4999) );
  HS65_LL_OAI12X2 U7113 ( .A(n4725), .B(n4718), .C(n4720), .Z(n3268) );
  HS65_LL_NAND2X5 U3540 ( .A(n3186), .B(n3185), .Z(n5066) );
  HS65_LH_IVX2 U8147 ( .A(n4958), .Z(n4959) );
  HS65_LH_IVX2 U8150 ( .A(n4964), .Z(n4965) );
  HS65_LH_NOR2X3 U3972 ( .A(n5036), .B(n5335), .Z(n5407) );
  HS65_LH_IVX2 U7110 ( .A(n3896), .Z(n3897) );
  HS65_LH_IVX2 U7132 ( .A(n5361), .Z(n4888) );
  HS65_LH_IVX2 U7147 ( .A(n5366), .Z(n4887) );
  HS65_LH_IVX2 U7609 ( .A(n5335), .Z(n4876) );
  HS65_LL_NAND2X4 U6530 ( .A(\lte_x_57/B[25] ), .B(n3247), .Z(n5259) );
  HS65_LH_IVX4 U4455 ( .A(n3756), .Z(n3757) );
  HS65_LL_OAI12X2 U8195 ( .A(n5453), .B(n5011), .C(n5445), .Z(n4929) );
  HS65_LH_IVX2 U8186 ( .A(n5375), .Z(n5035) );
  HS65_LH_NOR2X6 U6523 ( .A(\lte_x_57/B[25] ), .B(n3247), .Z(n3372) );
  HS65_LH_IVX7 U3991 ( .A(n4578), .Z(n3420) );
  HS65_LH_NAND2X4 U8773 ( .A(\lte_x_57/B[29] ), .B(n3204), .Z(n5147) );
  HS65_LH_AOI21X2 U6505 ( .A(n5284), .B(n5004), .C(n5304), .Z(n4002) );
  HS65_LL_NAND2X5 U4445 ( .A(n3834), .B(n3241), .Z(n4147) );
  HS65_LH_NOR2X3 U8143 ( .A(\lte_x_57/B[28] ), .B(n2791), .Z(n5141) );
  HS65_LL_NAND2X4 U6496 ( .A(\lte_x_57/B[6] ), .B(n5089), .Z(n4820) );
  HS65_LH_NOR2X3 U4479 ( .A(n5311), .B(n3338), .Z(n3329) );
  HS65_LH_IVX4 U6427 ( .A(n4023), .Z(n4024) );
  HS65_LH_NAND2X7 U4851 ( .A(\sub_x_51/A[5] ), .B(n2787), .Z(n3767) );
  HS65_LH_NAND2X5 U6506 ( .A(n3951), .B(n5089), .Z(n5350) );
  HS65_LH_NOR2X3 U4055 ( .A(n5016), .B(n3338), .Z(n3820) );
  HS65_LH_NOR2X3 U4463 ( .A(n3160), .B(n3322), .Z(n3489) );
  HS65_LLS_XOR2X3 U8209 ( .A(\lte_x_57/B[25] ), .B(n5072), .Z(n4988) );
  HS65_LH_IVX2 U7702 ( .A(n4775), .Z(n4776) );
  HS65_LL_OAI12X2 U7099 ( .A(n3673), .B(n4258), .C(n3675), .Z(n3260) );
  HS65_LH_IVX2 U7091 ( .A(n4799), .Z(n4800) );
  HS65_LH_CNIVX3 U4461 ( .A(n3580), .Z(n3582) );
  HS65_LL_NOR2X2 U3773 ( .A(n5371), .B(n5372), .Z(n5427) );
  HS65_LL_CNIVX3 U3593 ( .A(n4594), .Z(n5451) );
  HS65_LL_NAND2X4 U5429 ( .A(\lte_x_57/B[6] ), .B(n2998), .Z(n4861) );
  HS65_LH_IVX4 U4886 ( .A(n4316), .Z(n3400) );
  HS65_LH_IVX4 U4021 ( .A(n3888), .Z(n3614) );
  HS65_LH_NAND2X7 U4798 ( .A(\lte_x_57/B[3] ), .B(n2995), .Z(n4767) );
  HS65_LL_IVX7 U5503 ( .A(n5092), .Z(n2994) );
  HS65_LH_IVX4 U4856 ( .A(n5259), .Z(n5316) );
  HS65_LH_NAND2X5 U4830 ( .A(n3758), .B(n3757), .Z(n3763) );
  HS65_LL_OAI12X2 U5464 ( .A(n5131), .B(n4701), .C(n4703), .Z(n5253) );
  HS65_LH_NAND2X7 U4844 ( .A(n5517), .B(n4958), .Z(n4331) );
  HS65_LL_AOI12X2 U8330 ( .A(n4687), .B(n4686), .C(n4685), .Z(n4688) );
  HS65_LL_NOR2X2 U5478 ( .A(n5066), .B(\sub_x_51/A[21] ), .Z(n4486) );
  HS65_LH_NAND2X4 U6452 ( .A(n4602), .B(n3246), .Z(n4608) );
  HS65_LL_OAI12X2 U8223 ( .A(n3372), .B(n4552), .C(n5259), .Z(n5261) );
  HS65_LH_IVX2 U7605 ( .A(n5354), .Z(n5023) );
  HS65_LH_IVX4 U3986 ( .A(n5371), .Z(n5024) );
  HS65_LH_IVX4 U8365 ( .A(n4541), .Z(n4398) );
  HS65_LL_IVX9 U5531 ( .A(n3225), .Z(n2796) );
  HS65_LH_IVX2 U4002 ( .A(n5009), .Z(n5317) );
  HS65_LH_NAND2X7 U6349 ( .A(n5232), .B(n5355), .Z(n4096) );
  HS65_LL_IVX13 U3556 ( .A(n2829), .Z(n3742) );
  HS65_LL_OAI12X2 U8129 ( .A(n5219), .B(n4270), .C(n4272), .Z(n5101) );
  HS65_LH_IVX4 U8350 ( .A(n4701), .Z(n4702) );
  HS65_LH_AOI31X2 U4006 ( .A(n2780), .B(n5487), .C(n5417), .D(n5343), .Z(n5345) );
  HS65_LL_NAND2X2 U5444 ( .A(n5259), .B(n4594), .Z(n5439) );
  HS65_LL_NOR2X2 U6464 ( .A(n5191), .B(n4592), .Z(n3201) );
  HS65_LH_OAI12X2 U3997 ( .A(n5141), .B(n5009), .C(n5140), .Z(n5142) );
  HS65_LH_IVX2 U8317 ( .A(n4190), .Z(n4196) );
  HS65_LH_IVX2 U7072 ( .A(n3955), .Z(n3956) );
  HS65_LH_CNIVX3 U4766 ( .A(n4259), .Z(n4262) );
  HS65_LL_NAND2X4 U8645 ( .A(n2780), .B(n4208), .Z(n5502) );
  HS65_LH_NAND2X7 U4009 ( .A(n4725), .B(n2783), .Z(n4139) );
  HS65_LL_OAI12X2 U8144 ( .A(n5259), .B(n5139), .C(n4594), .Z(n5144) );
  HS65_LH_NOR2X3 U4872 ( .A(n4533), .B(n3322), .Z(n3594) );
  HS65_LH_AOI22X1 U5624 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][3] ), .B(n9162), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][3] ), .D(
        n9190), .Z(n6443) );
  HS65_LH_AOI22X1 U6609 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][3] ), .B(n9196), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][3] ), .D(
        n9192), .Z(n6440) );
  HS65_LL_NAND2AX4 U5349 ( .A(n4738), .B(n3593), .Z(n4292) );
  HS65_LH_NAND2X5 U6430 ( .A(n5140), .B(n4398), .Z(n4404) );
  HS65_LH_NAND2X2 U6593 ( .A(n4781), .B(n9538), .Z(n3799) );
  HS65_LH_OAI12X3 U4804 ( .A(n5266), .B(n5436), .C(n5446), .Z(n5267) );
  HS65_LH_CNIVX3 U5518 ( .A(n4187), .Z(n4188) );
  HS65_LH_NAND2X2 U4416 ( .A(n5074), .B(n5143), .Z(n5075) );
  HS65_LH_CNIVX3 U4795 ( .A(n5439), .Z(n5012) );
  HS65_LH_IVX7 U3990 ( .A(n4859), .Z(n4860) );
  HS65_LL_AOI12X2 U8178 ( .A(n5453), .B(n5317), .C(n5454), .Z(n5319) );
  HS65_LH_IVX2 U8171 ( .A(n5427), .Z(n5390) );
  HS65_LH_IVX4 U4812 ( .A(n4448), .Z(n4449) );
  HS65_LL_AOI12X2 U6395 ( .A(n5446), .B(n5314), .C(n5313), .Z(n5322) );
  HS65_LH_IVX2 U7086 ( .A(n5412), .Z(n5414) );
  HS65_LH_NAND2X5 U6402 ( .A(n4703), .B(n4702), .Z(n4717) );
  HS65_LH_IVX9 U5387 ( .A(n3453), .Z(n4490) );
  HS65_LH_IVX2 U8346 ( .A(n4238), .Z(n4241) );
  HS65_LH_IVX4 U3980 ( .A(n4637), .Z(n3206) );
  HS65_LH_NAND2X4 U8138 ( .A(n3128), .B(n3187), .Z(n5126) );
  HS65_LH_CNIVX3 U4393 ( .A(n4640), .Z(n3205) );
  HS65_LH_IVX2 U7707 ( .A(n3714), .Z(n3408) );
  HS65_LL_AOI12X2 U7079 ( .A(\sub_x_51/A[13] ), .B(n4208), .C(n3740), .Z(n3744) );
  HS65_LH_NAND2X5 U4361 ( .A(n4272), .B(n4271), .Z(n4274) );
  HS65_LH_NAND2X2 U4432 ( .A(n3465), .B(n4988), .Z(n3385) );
  HS65_LL_AOI12X2 U7114 ( .A(\lte_x_57/B[14] ), .B(n3742), .C(n3741), .Z(n3743) );
  HS65_LH_NAND2X2 U8702 ( .A(n4781), .B(n5208), .Z(n3856) );
  HS65_LL_NOR2X2 U4763 ( .A(n3664), .B(n5200), .Z(n3077) );
  HS65_LH_NAND2X7 U4396 ( .A(n5234), .B(n5030), .Z(n3894) );
  HS65_LL_OAI12X3 U3846 ( .A(n5109), .B(n5391), .C(n5232), .Z(n3885) );
  HS65_LH_NAND2X5 U6412 ( .A(n3842), .B(n3841), .Z(n3843) );
  HS65_LH_NOR2X5 U4444 ( .A(n3848), .B(n3860), .Z(n4125) );
  HS65_LH_CNIVX3 U3994 ( .A(n4984), .Z(n4991) );
  HS65_LH_NAND2X4 U4417 ( .A(n5151), .B(n5071), .Z(n5154) );
  HS65_LH_NAND2X4 U4855 ( .A(\lte_x_57/B[15] ), .B(n3742), .Z(n3581) );
  HS65_LH_IVX2 U8217 ( .A(n4209), .Z(n4210) );
  HS65_LL_AOI12X2 U8298 ( .A(n3379), .B(n4027), .C(n4032), .Z(n4028) );
  HS65_LL_NOR2X5 U3510 ( .A(n4440), .B(n4147), .Z(n4743) );
  HS65_LH_IVX2 U8341 ( .A(n4126), .Z(n3227) );
  HS65_LH_IVX2 U8255 ( .A(n4125), .Z(n3226) );
  HS65_LH_IVX2 U8747 ( .A(n5342), .Z(n4875) );
  HS65_LH_IVX2 U8782 ( .A(n5434), .Z(n5291) );
  HS65_LH_IVX2 U7695 ( .A(n5347), .Z(n4874) );
  HS65_LH_IVX2 U8607 ( .A(n3484), .Z(n3288) );
  HS65_LH_IVX2 U5422 ( .A(n3926), .Z(n3927) );
  HS65_LH_IVX2 U8253 ( .A(n4127), .Z(n3231) );
  HS65_LH_AOI211X1 U7040 ( .A(n5417), .B(n4872), .C(n5342), .D(n5415), .Z(
        n4873) );
  HS65_LH_IVX2 U8254 ( .A(n4128), .Z(n3230) );
  HS65_LH_IVX2 U8261 ( .A(n3917), .Z(n3918) );
  HS65_LH_IVX2 U3772 ( .A(n5387), .Z(n5025) );
  HS65_LH_NAND3X3 U4823 ( .A(n3488), .B(n3575), .C(n3295), .Z(n4616) );
  HS65_LL_AOI12X2 U5282 ( .A(n5320), .B(n5319), .C(n5318), .Z(n5321) );
  HS65_LH_OAI21X2 U3966 ( .A(n3954), .B(n3953), .C(n3952), .Z(n3958) );
  HS65_LH_OAI21X3 U4433 ( .A(n4901), .B(n3322), .C(n3398), .Z(n3712) );
  HS65_LH_NAND2X7 U3959 ( .A(n4861), .B(n4860), .Z(n4866) );
  HS65_LH_NAND2X7 U3842 ( .A(n3744), .B(n3743), .Z(n4038) );
  HS65_LL_AOI12X2 U5362 ( .A(n3255), .B(n4821), .C(n3254), .Z(n3256) );
  HS65_LH_NOR2X2 U4391 ( .A(n5085), .B(n4427), .Z(n5117) );
  HS65_LH_IVX2 U8201 ( .A(n3992), .Z(n3999) );
  HS65_LH_AOI12X4 U5468 ( .A(\lte_x_57/B[30] ), .B(n5496), .C(n3482), .Z(n3483) );
  HS65_LH_IVX2 U8321 ( .A(n4375), .Z(n4378) );
  HS65_LH_CNIVX3 U4382 ( .A(n4376), .Z(n4377) );
  HS65_LH_IVX9 U5368 ( .A(n4184), .Z(n4769) );
  HS65_LH_NAND2X5 U3960 ( .A(n4488), .B(n4490), .Z(n3457) );
  HS65_LH_NOR2X2 U6383 ( .A(n5247), .B(n5184), .Z(n5129) );
  HS65_LL_OAI12X2 U8139 ( .A(n4460), .B(n4709), .C(n5131), .Z(n5135) );
  HS65_LL_NOR2AX3 U6477 ( .A(n5496), .B(n3951), .Z(n3845) );
  HS65_LH_CNIVX3 U8278 ( .A(n4821), .Z(n4340) );
  HS65_LH_AOI211X1 U3491 ( .A(n5404), .B(n4894), .C(n5332), .D(n4893), .Z(
        n4900) );
  HS65_LL_OAI12X2 U8225 ( .A(n5433), .B(n4458), .C(n4460), .Z(n5254) );
  HS65_LH_IVX2 U8698 ( .A(n3806), .Z(n3809) );
  HS65_LH_NAND3X3 U4380 ( .A(n5449), .B(n4009), .C(n4008), .Z(n4010) );
  HS65_LL_IVX9 U5331 ( .A(n4321), .Z(n4225) );
  HS65_LL_OAI12X3 U3754 ( .A(n5433), .B(n4458), .C(n4460), .Z(n4707) );
  HS65_LH_NAND2X4 U5415 ( .A(n4367), .B(n4366), .Z(n4373) );
  HS65_LH_OAI21X3 U5274 ( .A(n4753), .B(n4468), .C(n4467), .Z(n4469) );
  HS65_LH_AOI12X2 U4363 ( .A(n4366), .B(n4369), .C(n5294), .Z(n3634) );
  HS65_LL_IVX4 U8697 ( .A(n3760), .Z(n4822) );
  HS65_LH_OAI21X3 U6331 ( .A(n3330), .B(n4326), .C(n4673), .Z(n4327) );
  HS65_LH_IVX2 U6337 ( .A(n4368), .Z(n4371) );
  HS65_LH_OAI21X3 U7016 ( .A(n5240), .B(n5239), .C(n5238), .Z(n5241) );
  HS65_LH_NAND2AX4 U5403 ( .A(n3403), .B(n3402), .Z(n3405) );
  HS65_LL_NOR2X2 U3797 ( .A(n3467), .B(n4750), .Z(n4471) );
  HS65_LH_NAND2X7 U7102 ( .A(n3730), .B(n4777), .Z(n3339) );
  HS65_LL_NAND3X3 U3811 ( .A(n3581), .B(n3646), .C(n3471), .Z(n4567) );
  HS65_LL_AOI12X2 U3495 ( .A(n4707), .B(n3197), .C(n3196), .Z(n3198) );
  HS65_LH_CBI4I6X2 U4338 ( .A(n4900), .B(n4899), .C(n4898), .D(n4897), .Z(
        n4908) );
  HS65_LL_NAND2X5 U3532 ( .A(n4411), .B(n3326), .Z(n4659) );
  HS65_LL_NAND3X3 U3511 ( .A(n3460), .B(n3851), .C(n3459), .Z(n3836) );
  HS65_LL_OAI12X2 U6343 ( .A(n4818), .B(n4340), .C(n4820), .Z(n4341) );
  HS65_LH_IVX2 U7703 ( .A(n4793), .Z(n4798) );
  HS65_LH_NOR2X3 U3948 ( .A(n4007), .B(n5260), .Z(n4013) );
  HS65_LH_OAI21X2 U5283 ( .A(n2855), .B(n3918), .C(n4743), .Z(n3919) );
  HS65_LH_IVX2 U7037 ( .A(n5250), .Z(n3997) );
  HS65_LL_NOR2X2 U3975 ( .A(n4812), .B(n4514), .Z(n3796) );
  HS65_LH_AOI211X1 U6308 ( .A(n5420), .B(n4875), .C(n4874), .D(n4873), .Z(
        n4891) );
  HS65_LH_IVX2 U7025 ( .A(n5462), .Z(n5464) );
  HS65_LHS_XNOR2X3 U5325 ( .A(n4806), .B(n4805), .Z(n4807) );
  HS65_LL_NAND2X7 U8687 ( .A(n4433), .B(n4842), .Z(n4792) );
  HS65_LH_OAI21X3 U5300 ( .A(n5272), .B(n5271), .C(n5270), .Z(n5273) );
  HS65_LH_IVX2 U6360 ( .A(n4707), .Z(n4708) );
  HS65_LH_NOR2X5 U4407 ( .A(n3827), .B(n3570), .Z(n3571) );
  HS65_LL_NOR2X3 U3790 ( .A(n3689), .B(n3688), .Z(n4308) );
  HS65_LH_OAI21X3 U8290 ( .A(n3193), .B(n4846), .C(n4471), .Z(n4472) );
  HS65_LL_IVX7 U6286 ( .A(n4659), .Z(n5510) );
  HS65_LL_NAND2X4 U3782 ( .A(n4368), .B(n3191), .Z(n4104) );
  HS65_LL_IVX9 U4340 ( .A(n4792), .Z(n5484) );
  HS65_LH_OAI12X3 U8267 ( .A(n4840), .B(n5499), .C(n4248), .Z(n4249) );
  HS65_LL_NAND2X2 U5246 ( .A(n3379), .B(n3294), .Z(n4500) );
  HS65_LL_NOR2X5 U3786 ( .A(n3340), .B(n3339), .Z(n4332) );
  HS65_LH_NOR2X2 U3927 ( .A(n5087), .B(n5121), .Z(n5124) );
  HS65_LH_OAI211X3 U3912 ( .A(n3079), .B(n4846), .C(n4150), .D(n3577), .Z(
        n3578) );
  HS65_LH_OAI21X2 U4746 ( .A(n5121), .B(n5120), .C(n5119), .Z(n5122) );
  HS65_LH_IVX7 U4351 ( .A(n4905), .Z(n4923) );
  HS65_LL_OAI12X3 U7017 ( .A(n4262), .B(n2823), .C(n4261), .Z(n4263) );
  HS65_LH_NOR3X3 U4742 ( .A(n5022), .B(n5021), .C(n5020), .Z(n5058) );
  HS65_LH_NOR2X2 U4354 ( .A(n5069), .B(n5138), .Z(n5076) );
  HS65_LL_IVX7 U5238 ( .A(n5499), .Z(n4836) );
  HS65_LL_AOI12X2 U5242 ( .A(n3285), .B(n4119), .C(n4750), .Z(n4405) );
  HS65_LH_NAND2X4 U3909 ( .A(n4294), .B(n4066), .Z(n4067) );
  HS65_LH_NAND2X5 U4744 ( .A(n4671), .B(n4567), .Z(n3833) );
  HS65_LH_IVX7 U4764 ( .A(n4381), .Z(n4617) );
  HS65_LH_IVX4 U4740 ( .A(n2823), .Z(n3607) );
  HS65_LH_OAI21X3 U5290 ( .A(n4292), .B(n4034), .C(n4033), .Z(n4035) );
  HS65_LHS_XNOR2X6 U3698 ( .A(n3843), .B(n4863), .Z(n3881) );
  HS65_LL_NOR2X2 U5263 ( .A(n2830), .B(n5499), .Z(n4197) );
  HS65_LL_OAI12X3 U3638 ( .A(n4275), .B(n2823), .C(n4277), .Z(n4049) );
  HS65_LL_OAI13X1 U4722 ( .A(n4891), .B(n4899), .C(n4890), .D(n4889), .Z(n4909) );
  HS65_LH_OAI22X3 U3905 ( .A(n5499), .B(n4624), .C(n4665), .D(n4623), .Z(n4625) );
  HS65_LL_OAI22X1 U7001 ( .A(n4747), .B(n4332), .C(n5499), .D(n4791), .Z(n3707) );
  HS65_LH_NAND2X7 U4326 ( .A(n4836), .B(n4793), .Z(n4318) );
  HS65_LL_OAI12X2 U6232 ( .A(n4838), .B(n4837), .C(n4836), .Z(n4839) );
  HS65_LL_AOI22X1 U3896 ( .A(n5510), .B(n4742), .C(n5505), .D(n3693), .Z(n3703) );
  HS65_LL_NAND2X2 U3596 ( .A(n5511), .B(n5510), .Z(n5512) );
  HS65_LH_CBI4I1X3 U3898 ( .A(n2792), .B(\u_DataPath/u_execute/A_inALU_i[26] ), 
        .C(n4509), .D(n5510), .Z(n4510) );
  HS65_LL_AOI12X2 U7007 ( .A(n5157), .B(n5156), .C(n5155), .Z(n5158) );
  HS65_LL_IVX2 U6228 ( .A(n5165), .Z(n5167) );
  HS65_LL_IVX2 U4730 ( .A(n4692), .Z(n4579) );
  HS65_LH_NAND2X4 U3894 ( .A(n5484), .B(n4290), .Z(n4157) );
  HS65_LL_NAND2AX4 U6326 ( .A(n3850), .B(n3849), .Z(n5479) );
  HS65_LL_AOI12X2 U5250 ( .A(n4577), .B(n4692), .C(n3420), .Z(n3421) );
  HS65_LH_IVX9 U4758 ( .A(n4745), .Z(n4672) );
  HS65_LL_OAI12X2 U3776 ( .A(n3809), .B(n3808), .C(n4836), .Z(n3810) );
  HS65_LL_AOI12X2 U3494 ( .A(n4721), .B(n4729), .C(n4724), .Z(n4136) );
  HS65_LL_AOI12X2 U4329 ( .A(n5510), .B(n4569), .C(n4568), .Z(n4586) );
  HS65_LH_IVX2 U4331 ( .A(n4197), .Z(n3804) );
  HS65_LL_AOI12X2 U4743 ( .A(n4490), .B(n4729), .C(n4489), .Z(n4491) );
  HS65_LH_NAND2X4 U3911 ( .A(n5211), .B(n3837), .Z(n3838) );
  HS65_LH_NAND2X2 U5233 ( .A(n5484), .B(n4477), .Z(n4069) );
  HS65_LL_AOI12X2 U6257 ( .A(n4604), .B(n4692), .C(n4603), .Z(n4605) );
  HS65_LH_OA12X9 U3906 ( .A(n4659), .B(n4332), .C(n4331), .Z(n2827) );
  HS65_LL_OAI12X2 U5296 ( .A(n4381), .B(n4747), .C(n4117), .Z(n4123) );
  HS65_LL_AOI12X2 U8289 ( .A(n5510), .B(n4473), .C(n4472), .Z(n4474) );
  HS65_LL_AOI12X2 U8336 ( .A(n4294), .B(n3801), .C(n3800), .Z(n3815) );
  HS65_LL_OAI12X2 U8647 ( .A(n4613), .B(n3494), .C(n3493), .Z(n3495) );
  HS65_LH_NOR2X5 U4323 ( .A(n4738), .B(n4737), .Z(n4760) );
  HS65_LL_AOI12X2 U8783 ( .A(n5331), .B(n5380), .C(n5330), .Z(n5478) );
  HS65_LL_AOI12X2 U8240 ( .A(n5124), .B(n5123), .C(n5122), .Z(n5159) );
  HS65_LH_OAI21X2 U5204 ( .A(n4292), .B(n4070), .C(n4069), .Z(n4071) );
  HS65_LL_AOI12X2 U4322 ( .A(n5243), .B(n5242), .C(n5241), .Z(n5277) );
  HS65_LH_NAND3X3 U6962 ( .A(n4670), .B(n4669), .C(n4668), .Z(n4678) );
  HS65_LL_OAI12X2 U6217 ( .A(n4909), .B(n4908), .C(n4907), .Z(n4941) );
  HS65_LL_OAI12X2 U3879 ( .A(n4378), .B(n4695), .C(n4377), .Z(n4379) );
  HS65_LL_AOI12X2 U4328 ( .A(n4836), .B(n3801), .C(n3739), .Z(n3748) );
  HS65_LL_OAI12X2 U3814 ( .A(n4659), .B(n4441), .C(n3745), .Z(n3746) );
  HS65_LL_AOI12X2 U3505 ( .A(n5510), .B(n4466), .C(n4040), .Z(n4041) );
  HS65_LL_OAI12X2 U5198 ( .A(n3279), .B(n4695), .C(n3278), .Z(n3280) );
  HS65_LL_OAI12X2 U6169 ( .A(n4580), .B(n4695), .C(n4579), .Z(n4581) );
  HS65_LH_NAND2X4 U3883 ( .A(n5048), .B(n5047), .Z(n5049) );
  HS65_LL_OAI12X2 U6957 ( .A(n4241), .B(n4273), .C(n4240), .Z(n4242) );
  HS65_LL_OAI12X2 U6936 ( .A(n4606), .B(n4695), .C(n4605), .Z(n4607) );
  HS65_LL_OAI12X2 U4313 ( .A(n3422), .B(n4695), .C(n3421), .Z(n3423) );
  HS65_LL_OAI21X2 U3833 ( .A(n4408), .B(n4901), .C(n4407), .Z(n4409) );
  HS65_LL_OAI12X2 U8715 ( .A(n4094), .B(n4273), .C(n4093), .Z(n4095) );
  HS65_LL_OAI12X2 U6961 ( .A(n4177), .B(n4273), .C(n4176), .Z(n4178) );
  HS65_LL_NOR2AX13 U3504 ( .A(n3085), .B(n3084), .Z(n4714) );
  HS65_LH_AO22X9 U6227 ( .A(n4950), .B(n5517), .C(n4433), .D(n5485), .Z(n3653)
         );
  HS65_LL_OAI12X2 U5197 ( .A(n4416), .B(n4695), .C(n4415), .Z(n4417) );
  HS65_LH_NOR2X3 U3633 ( .A(n4665), .B(n4563), .Z(n3474) );
  HS65_LL_OAI12X2 U6939 ( .A(n4371), .B(n4714), .C(n4370), .Z(n4372) );
  HS65_LL_NAND3X2 U3760 ( .A(n3815), .B(n3814), .C(n3813), .Z(n3816) );
  HS65_LL_OAI12X2 U4695 ( .A(n4714), .B(n4598), .C(n4597), .Z(n4599) );
  HS65_LL_NAND2X2 U3877 ( .A(n5050), .B(n5049), .Z(n5056) );
  HS65_LL_OAI12X2 U4696 ( .A(n4715), .B(n4714), .C(n4713), .Z(n4716) );
  HS65_LL_NAND2X2 U3871 ( .A(n4267), .B(n4266), .Z(n4268) );
  HS65_LL_AO112X4 U3775 ( .A(n7325), .B(n4633), .C(n4632), .D(n4631), .Z(n4634) );
  HS65_LL_NAND2X2 U4308 ( .A(n7325), .B(n3365), .Z(n3366) );
  HS65_LL_NAND2X2 U4304 ( .A(n4699), .B(n4698), .Z(n4700) );
  HS65_LH_IVX9 U5183 ( .A(n5524), .Z(n5525) );
  HS65_LL_IVX2 U4676 ( .A(n4100), .Z(n4101) );
  HS65_LH_IVX9 U6543 ( .A(n8645), .Z(\u_DataPath/jump_address_i [12]) );
  HS65_LH_NOR2X6 U5919 ( .A(n8975), .B(n9050), .Z(n5820) );
  HS65_LH_NAND2X7 U5047 ( .A(n9358), .B(n9148), .Z(n7622) );
  HS65_LH_IVX7 U4569 ( .A(n8741), .Z(n3109) );
  HS65_LH_AOI22X3 U9617 ( .A(n8687), .B(n9426), .C(n9252), .D(n9079), .Z(n8283) );
  HS65_LH_NAND2X5 U8386 ( .A(n9359), .B(n9181), .Z(n7625) );
  HS65_LH_AOI12X6 U3570 ( .A(n9425), .B(\u_DataPath/from_mem_data_out_i [0]), 
        .C(n8935), .Z(n8278) );
  HS65_LHS_XOR2X6 U6830 ( .A(n9464), .B(n9112), .Z(n7206) );
  HS65_LH_IVX7 U5902 ( .A(n5646), .Z(n5705) );
  HS65_LH_AOI12X2 U3515 ( .A(n8976), .B(n5819), .C(n9307), .Z(n5751) );
  HS65_LL_IVX13 U4143 ( .A(n3107), .Z(n3178) );
  HS65_LH_AOI12X2 U7325 ( .A(n8988), .B(n5908), .C(n8712), .Z(n5902) );
  HS65_LH_IVX4 U8393 ( .A(n8278), .Z(n2955) );
  HS65_LH_IVX18 U3567 ( .A(n3149), .Z(n2778) );
  HS65_LH_NAND2X4 U4476 ( .A(n9332), .B(n2797), .Z(n3059) );
  HS65_LH_NOR2X5 U4532 ( .A(n8625), .B(n3181), .Z(n3123) );
  HS65_LL_NAND3X5 U5899 ( .A(n7209), .B(n7208), .C(n7207), .Z(n7212) );
  HS65_LH_NAND2AX4 U7527 ( .A(n8657), .B(n3090), .Z(n3983) );
  HS65_LL_AOI12X2 U4548 ( .A(n9030), .B(n5717), .C(n9298), .Z(n5641) );
  HS65_LH_NAND2X4 U4106 ( .A(n3090), .B(n8443), .Z(n3165) );
  HS65_LH_NOR2X3 U4128 ( .A(n3174), .B(n8438), .Z(n3168) );
  HS65_LH_NOR2X5 U6730 ( .A(n3174), .B(n8390), .Z(n2932) );
  HS65_LH_NAND2X7 U4220 ( .A(n3174), .B(n9428), .Z(n2933) );
  HS65_LL_OAI112X4 U7259 ( .A(n9336), .B(n3149), .C(n3024), .D(n3023), .Z(
        \sub_x_51/A[8] ) );
  HS65_LL_AOI12X2 U8211 ( .A(n8702), .B(n2798), .C(n3035), .Z(n3036) );
  HS65_LH_IVX7 U3770 ( .A(n8412), .Z(n3070) );
  HS65_LH_NAND2X7 U4286 ( .A(\u_DataPath/cw_to_ex_i [2]), .B(
        \u_DataPath/cw_to_ex_i [1]), .Z(n2862) );
  HS65_LL_NAND2X7 U3806 ( .A(n2806), .B(n3110), .Z(
        \u_DataPath/u_execute/A_inALU_i[26] ) );
  HS65_LL_NAND2X4 U4984 ( .A(n8374), .B(n5183), .Z(n2963) );
  HS65_LH_AOI12X2 U7290 ( .A(n9235), .B(n5888), .C(n9275), .Z(n5806) );
  HS65_LH_NAND2X7 U7307 ( .A(n9110), .B(n8457), .Z(n8046) );
  HS65_LH_NOR2X5 U4983 ( .A(n2955), .B(n2794), .Z(n8369) );
  HS65_LH_IVX9 U4998 ( .A(\sub_x_51/A[8] ), .Z(n4283) );
  HS65_LL_AOI21X2 U3681 ( .A(Data_out_fromRAM[15]), .B(n8165), .C(n7312), .Z(
        n7313) );
  HS65_LL_NAND2X5 U5133 ( .A(n3283), .B(n4018), .Z(n3245) );
  HS65_LH_IVX9 U3690 ( .A(n3245), .Z(n3292) );
  HS65_LL_AOI12X2 U5766 ( .A(n8889), .B(n5725), .C(n9305), .Z(n5584) );
  HS65_LL_NAND2X5 U3817 ( .A(n3022), .B(n3021), .Z(n5386) );
  HS65_LL_NOR2X3 U3675 ( .A(n3213), .B(n3245), .Z(n3834) );
  HS65_LL_CNIVX3 U4875 ( .A(n3949), .Z(n2787) );
  HS65_LH_NAND2X7 U4042 ( .A(n5312), .B(n5311), .Z(n5309) );
  HS65_LH_NAND2X7 U7172 ( .A(n2825), .B(n5251), .Z(n5298) );
  HS65_LH_NAND2X5 U6488 ( .A(n3039), .B(n3073), .Z(n5227) );
  HS65_LH_NOR2X5 U8707 ( .A(n3950), .B(n3949), .Z(n5334) );
  HS65_LL_NAND2X4 U5559 ( .A(n4383), .B(n5063), .Z(n5295) );
  HS65_LH_AOI22X3 U8096 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][0] ), .B(n9159), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][0] ), .D(n8862), .Z(n7295) );
  HS65_LH_AOI22X3 U8089 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][0] ), .B(n9062), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][0] ), .D(n8863), .Z(n7289) );
  HS65_LH_AOI22X3 U8091 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][0] ), .B(n8865), 
        .C(n8864), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][0] ), .Z(n7290)
         );
  HS65_LH_NAND2X7 U5399 ( .A(n4048), .B(n4047), .Z(n4050) );
  HS65_LH_IVX7 U3785 ( .A(n4727), .Z(n2783) );
  HS65_LH_NOR2X5 U8111 ( .A(n5192), .B(n3200), .Z(n5132) );
  HS65_LH_IVX9 U5379 ( .A(n3676), .Z(n4257) );
  HS65_LH_IVX7 U3595 ( .A(n5454), .Z(n5008) );
  HS65_LH_NOR2X5 U8168 ( .A(\lte_x_57/B[10] ), .B(n3074), .Z(n5200) );
  HS65_LH_IVX4 U4033 ( .A(n3903), .Z(n3606) );
  HS65_LH_NAND2X5 U8137 ( .A(\sub_x_51/A[18] ), .B(n3188), .Z(n5125) );
  HS65_LH_IVX4 U8370 ( .A(n4275), .Z(n4276) );
  HS65_LHS_XNOR2X3 U5604 ( .A(n8993), .B(n5729), .Z(\u_DataPath/toPC2_i [25])
         );
  HS65_LH_NOR2X5 U5461 ( .A(n5139), .B(n5191), .Z(n5262) );
  HS65_LH_IVX7 U4012 ( .A(n4709), .Z(n4103) );
  HS65_LH_NOR2X5 U5463 ( .A(n5264), .B(n5141), .Z(n5197) );
  HS65_LL_NOR2X6 U3798 ( .A(n5148), .B(n4784), .Z(n4750) );
  HS65_LH_NOR2X6 U5524 ( .A(n5148), .B(n3322), .Z(n3482) );
  HS65_LH_CNIVX3 U8342 ( .A(n3673), .Z(n3674) );
  HS65_LH_OAI21X2 U3969 ( .A(n4703), .B(n5132), .C(n4552), .Z(n5133) );
  HS65_LH_IVX7 U4864 ( .A(n4374), .Z(n3540) );
  HS65_LH_NAND2X7 U5475 ( .A(\sub_x_51/A[21] ), .B(n5066), .Z(n4487) );
  HS65_LH_NAND2X7 U4791 ( .A(n5227), .B(n4024), .Z(n4026) );
  HS65_LH_IVX7 U7071 ( .A(n4260), .Z(n4261) );
  HS65_LH_NOR2X5 U8231 ( .A(n2793), .B(n3078), .Z(n5204) );
  HS65_LH_NAND2X7 U4017 ( .A(n3901), .B(n3606), .Z(n3612) );
  HS65_LH_IVX4 U4016 ( .A(n4592), .Z(n4593) );
  HS65_LL_AOI22X1 U4049 ( .A(\u_DataPath/u_execute/A_inALU_i[26] ), .B(n3826), 
        .C(n2792), .D(\add_x_50/A[23] ), .Z(n3295) );
  HS65_LL_IVX7 U8613 ( .A(n4738), .Z(n4433) );
  HS65_LH_CNIVX3 U8301 ( .A(n3820), .Z(n3821) );
  HS65_LL_OAI12X3 U3691 ( .A(n8982), .B(n5768), .C(n9029), .Z(n5928) );
  HS65_LL_NOR2X3 U3794 ( .A(n5204), .B(n5391), .Z(n3883) );
  HS65_LH_NAND2X5 U3973 ( .A(n4594), .B(n4593), .Z(n4600) );
  HS65_LL_AOI12X2 U5560 ( .A(n8983), .B(n5928), .C(n9301), .Z(n5763) );
  HS65_LH_NOR2X5 U5580 ( .A(n4431), .B(n3338), .Z(n4503) );
  HS65_LH_NAND2X7 U3977 ( .A(n5219), .B(n4348), .Z(n4354) );
  HS65_LH_NAND2X4 U8693 ( .A(n2793), .B(n3742), .Z(n3683) );
  HS65_LHS_XNOR2X3 U4877 ( .A(n8992), .B(n5721), .Z(\u_DataPath/toPC2_i [27])
         );
  HS65_LH_NAND3X5 U3607 ( .A(n5286), .B(n5298), .C(n5285), .Z(n5306) );
  HS65_LH_NAND2X5 U6365 ( .A(n3675), .B(n3674), .Z(n3681) );
  HS65_LL_IVX2 U6436 ( .A(n4486), .Z(n3250) );
  HS65_LH_IVX9 U5411 ( .A(n5367), .Z(n5395) );
  HS65_LH_NAND2X7 U4404 ( .A(n5131), .B(n4103), .Z(n4109) );
  HS65_LH_NAND2X7 U6410 ( .A(\add_x_50/A[19] ), .B(n3189), .Z(n5434) );
  HS65_LH_NAND3X5 U5391 ( .A(n5388), .B(n3961), .C(n5237), .Z(n3969) );
  HS65_LH_IVX2 U8249 ( .A(n4595), .Z(n3312) );
  HS65_LH_NAND2X4 U8212 ( .A(n3128), .B(n3742), .Z(n3286) );
  HS65_LH_CNIVX3 U8618 ( .A(n3629), .Z(n3348) );
  HS65_LH_NAND2X5 U3937 ( .A(n5233), .B(n4175), .Z(n4179) );
  HS65_LH_NAND2X7 U4365 ( .A(n5111), .B(n3665), .Z(n3671) );
  HS65_LL_NOR2AX3 U3853 ( .A(n3250), .B(n3453), .Z(n4721) );
  HS65_LH_AOI211X2 U7009 ( .A(n4888), .B(n4887), .C(n5396), .D(n4886), .Z(
        n4889) );
  HS65_LL_NAND2X4 U3832 ( .A(n3478), .B(n3477), .Z(n4571) );
  HS65_LH_OAI21X3 U7117 ( .A(n4383), .B(n3322), .C(n3687), .Z(n3688) );
  HS65_LL_AOI22X1 U5462 ( .A(n2793), .B(n5496), .C(n5498), .D(\sub_x_51/A[13] ), .Z(n3224) );
  HS65_LH_AOI21X2 U3600 ( .A(n5114), .B(n5113), .C(n5112), .Z(n5120) );
  HS65_LH_NOR2X5 U5347 ( .A(n4859), .B(n4349), .Z(n4352) );
  HS65_LH_NAND2X4 U5412 ( .A(n4802), .B(n4217), .Z(n4218) );
  HS65_LH_OAI12X3 U6366 ( .A(n4804), .B(n4803), .C(n4802), .Z(n4805) );
  HS65_LL_AOI22X1 U8302 ( .A(\u_DataPath/u_execute/A_inALU_i[26] ), .B(n5496), 
        .C(n5498), .D(\sub_x_51/A[27] ), .Z(n3822) );
  HS65_LL_OAI12X3 U5510 ( .A(n8984), .B(n5763), .C(n9028), .Z(n5868) );
  HS65_LH_AOI22X1 U8238 ( .A(n5498), .B(n5497), .C(\lte_x_57/B[2] ), .D(n5496), 
        .Z(n5500) );
  HS65_LH_OAI12X3 U3499 ( .A(n4727), .B(n4726), .C(n4725), .Z(n4728) );
  HS65_LH_NAND2X4 U5333 ( .A(n5250), .B(n5188), .Z(n5189) );
  HS65_LH_OAI12X3 U6351 ( .A(n4770), .B(n4769), .C(n4768), .Z(n4771) );
  HS65_LH_IVX7 U3765 ( .A(n4643), .Z(n4399) );
  HS65_LHS_XNOR2X6 U7085 ( .A(n9133), .B(n5868), .Z(
        \u_DataPath/u_execute/resAdd1_i [30]) );
  HS65_LH_IVX7 U4782 ( .A(n3795), .Z(n3798) );
  HS65_LL_NAND2X4 U3851 ( .A(n3269), .B(n4721), .Z(n3271) );
  HS65_LH_NAND2X5 U6355 ( .A(n4460), .B(n4459), .Z(n4465) );
  HS65_LH_CNIVX3 U8251 ( .A(n4741), .Z(n3349) );
  HS65_LH_NOR3X4 U3984 ( .A(n3348), .B(n3716), .C(n3347), .Z(n4657) );
  HS65_LL_NAND2X2 U5245 ( .A(n3792), .B(n3791), .Z(n3793) );
  HS65_LH_OAI12X3 U6296 ( .A(n3679), .B(n2823), .C(n3678), .Z(n3680) );
  HS65_LH_OAI21X2 U6297 ( .A(n5138), .B(n5137), .C(n5136), .Z(n5157) );
  HS65_LH_OAI21X3 U6277 ( .A(n4838), .B(n4837), .C(n4294), .Z(n4215) );
  HS65_LL_AOI12X2 U7004 ( .A(n5505), .B(n4066), .C(n3728), .Z(n3751) );
  HS65_LH_NOR2X5 U5293 ( .A(n4727), .B(n4722), .Z(n4730) );
  HS65_LH_NOR2X5 U5302 ( .A(n5258), .B(n5189), .Z(n5199) );
  HS65_LL_NAND3X2 U6997 ( .A(n4152), .B(n4151), .C(n4150), .Z(n4154) );
  HS65_LH_NAND2X2 U4350 ( .A(n5492), .B(n4807), .Z(n4808) );
  HS65_LL_OAI12X3 U6392 ( .A(n8978), .B(n5668), .C(n9034), .Z(n5670) );
  HS65_LL_OAI12X2 U3804 ( .A(n5481), .B(n4333), .C(n3928), .Z(n3929) );
  HS65_LH_OAI12X3 U5275 ( .A(n5370), .B(n5369), .C(n5368), .Z(n5381) );
  HS65_LL_AOI13X2 U4724 ( .A(n5502), .B(n5501), .C(n5500), .D(n5499), .Z(n5503) );
  HS65_LH_NOR2X3 U3636 ( .A(n4659), .B(n4386), .Z(n4223) );
  HS65_LL_IVX9 U3839 ( .A(n4732), .Z(n4695) );
  HS65_LL_AOI12X2 U8373 ( .A(n5517), .B(n4848), .C(n4847), .Z(n4853) );
  HS65_LLS_XOR2X3 U3809 ( .A(n4825), .B(n4824), .Z(n4826) );
  HS65_LH_NAND2X4 U4729 ( .A(n5492), .B(n3877), .Z(n3878) );
  HS65_LH_NOR2X6 U4325 ( .A(n4329), .B(n4328), .Z(n4737) );
  HS65_LH_IVX9 U5273 ( .A(n5479), .Z(n5480) );
  HS65_LH_NOR2X5 U5195 ( .A(n4526), .B(n4695), .Z(n4527) );
  HS65_LL_AOI12X2 U8360 ( .A(n5510), .B(n4512), .C(n3409), .Z(n3410) );
  HS65_LL_NAND3X2 U3812 ( .A(n4060), .B(n4059), .C(n4058), .Z(n4061) );
  HS65_LL_OAI12X2 U3805 ( .A(n5481), .B(n4840), .C(n4839), .Z(n4841) );
  HS65_LH_NAND2X4 U3769 ( .A(n4596), .B(n4639), .Z(n4598) );
  HS65_LH_IVX9 U5212 ( .A(n4560), .Z(n4561) );
  HS65_LL_OAI21X2 U6202 ( .A(n4111), .B(n4659), .C(n4110), .Z(n4124) );
  HS65_LL_AOI21X2 U3834 ( .A(n4836), .B(n4573), .C(n4406), .Z(n4407) );
  HS65_LL_NAND3X2 U3838 ( .A(n4043), .B(n4042), .C(n4041), .Z(n4044) );
  HS65_LL_IVX2 U3622 ( .A(n3616), .Z(n3617) );
  HS65_LL_AOI21X2 U4700 ( .A(n4017), .B(n4016), .C(n4015), .Z(n4021) );
  HS65_LH_NAND2X4 U8282 ( .A(n4411), .B(n4535), .Z(n4074) );
  HS65_LL_AOI21X2 U6164 ( .A(n5492), .B(n3936), .C(n3935), .Z(n3937) );
  HS65_LL_NAND2X2 U3854 ( .A(n3415), .B(n3414), .Z(n3427) );
  HS65_LH_IVX7 U3872 ( .A(n3749), .Z(n3750) );
  HS65_LL_IVX2 U4681 ( .A(n3752), .Z(n3753) );
  HS65_LH_IVX2 U9391 ( .A(Data_out_fromRAM[17]), .Z(n8193) );
  HS65_LH_IVX2 U9388 ( .A(Data_out_fromRAM[21]), .Z(n8202) );
  HS65_LH_NOR2X3 U5861 ( .A(n9232), .B(n9403), .Z(n7443) );
  HS65_LH_IVX9 U3732 ( .A(n8655), .Z(\u_DataPath/jump_address_i [8]) );
  HS65_LH_NAND2X7 U3658 ( .A(n9042), .B(n9181), .Z(n7428) );
  HS65_LH_NAND2X7 U3673 ( .A(n9180), .B(n9181), .Z(n7629) );
  HS65_LL_IVX9 U4564 ( .A(n9012), .Z(n3107) );
  HS65_LL_IVX9 U3566 ( .A(n2800), .Z(n3980) );
  HS65_LH_NOR2X3 U7417 ( .A(n9541), .B(n2782), .Z(n8384) );
  HS65_LH_NOR2X5 U6765 ( .A(n9448), .B(n3980), .Z(n8390) );
  HS65_LL_CNBFX14 U4107 ( .A(n3149), .Z(n3181) );
  HS65_LH_NOR2X5 U4925 ( .A(n8659), .B(n2772), .Z(n8427) );
  HS65_LH_IVX9 U3714 ( .A(n3162), .Z(n8443) );
  HS65_LL_IVX18 U3568 ( .A(n3090), .Z(n3174) );
  HS65_LH_NOR2X2 U4630 ( .A(n3090), .B(n8730), .Z(n3089) );
  HS65_LH_NOR3X4 U4570 ( .A(n8898), .B(n9182), .C(n7349), .Z(n7945) );
  HS65_LH_NAND2X7 U3652 ( .A(n8701), .B(n2710), .Z(n3040) );
  HS65_LH_NAND2X4 U5008 ( .A(n8700), .B(n2798), .Z(n8416) );
  HS65_LH_OAI21X3 U4978 ( .A(n8626), .B(n3181), .C(n3045), .Z(n3046) );
  HS65_LL_NAND2X2 U4213 ( .A(n3184), .B(n8730), .Z(n3155) );
  HS65_LH_NAND2X5 U7458 ( .A(n3174), .B(n9433), .Z(n3022) );
  HS65_LH_NOR2X6 U3672 ( .A(n9458), .B(n7635), .Z(n7303) );
  HS65_LH_IVX18 U4079 ( .A(n3103), .Z(\sub_x_51/A[27] ) );
  HS65_LL_AOI12X2 U4534 ( .A(n9035), .B(n5932), .C(n9297), .Z(n5787) );
  HS65_LL_OAI13X5 U3791 ( .A(n5934), .B(n2940), .C(n8385), .D(n2939), .Z(n3949) );
  HS65_LL_IVX2 U5547 ( .A(n5251), .Z(n3194) );
  HS65_LL_NOR2X3 U6521 ( .A(n3160), .B(n5252), .Z(n5304) );
  HS65_LH_NOR2X3 U7608 ( .A(n3039), .B(n3073), .Z(n5080) );
  HS65_LH_AO22X9 U8093 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][0] ), .B(n9204), 
        .C(n9203), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][0] ), .Z(n7281)
         );
  HS65_LH_AO22X9 U8090 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][0] ), .B(n9102), 
        .C(n9101), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][0] ), .Z(n7292) );
  HS65_LH_NAND2X5 U8228 ( .A(\lte_x_57/B[15] ), .B(n2788), .Z(n5234) );
  HS65_LH_NAND2X7 U8772 ( .A(\lte_x_57/B[28] ), .B(n2791), .Z(n5140) );
  HS65_LL_AOI12X2 U5602 ( .A(n8973), .B(n5729), .C(n9308), .Z(n5565) );
  HS65_LH_NOR2X6 U8169 ( .A(\sub_x_51/A[27] ), .B(n4005), .Z(n5191) );
  HS65_LH_NOR2X5 U3592 ( .A(n5336), .B(n5335), .Z(n5403) );
  HS65_LH_NOR2X5 U8145 ( .A(\u_DataPath/u_execute/A_inALU_i[26] ), .B(n4622), 
        .Z(n5139) );
  HS65_LL_CNIVX3 U3641 ( .A(n4601), .Z(n3246) );
  HS65_LH_OR2X9 U4054 ( .A(n3103), .B(n3338), .Z(n3485) );
  HS65_LL_NAND2X4 U8140 ( .A(\sub_x_51/A[22] ), .B(n3194), .Z(n5131) );
  HS65_LH_IVX9 U3647 ( .A(n4812), .Z(n5486) );
  HS65_LH_IVX7 U5433 ( .A(n5070), .Z(n4540) );
  HS65_LH_NOR2X5 U6465 ( .A(n4918), .B(n5066), .Z(n5297) );
  HS65_LH_OAI12X3 U5375 ( .A(n4006), .B(n4594), .C(n5009), .Z(n5260) );
  HS65_LH_NAND2X4 U6507 ( .A(n5092), .B(n4192), .Z(n5043) );
  HS65_LH_NAND2X4 U8121 ( .A(n2793), .B(n3078), .Z(n5109) );
  HS65_LH_NAND2X7 U5479 ( .A(\sub_x_51/A[20] ), .B(n5064), .Z(n4488) );
  HS65_LH_OAI12X2 U3999 ( .A(n5147), .B(n5146), .C(n5145), .Z(n5150) );
  HS65_LH_NAND2X7 U8166 ( .A(n2793), .B(n3078), .Z(n5233) );
  HS65_LH_IVX2 U8327 ( .A(n4943), .Z(n4848) );
  HS65_LH_NOR2X6 U8110 ( .A(n2793), .B(n3078), .Z(n5110) );
  HS65_LH_NOR2X5 U8136 ( .A(\lte_x_57/B[11] ), .B(n3075), .Z(n5078) );
  HS65_LH_IVX4 U4005 ( .A(n5415), .Z(n5344) );
  HS65_LH_AOI21X2 U7708 ( .A(n4781), .B(n5186), .C(n4750), .Z(n3642) );
  HS65_LH_NAND2X2 U8695 ( .A(\sub_x_51/A[16] ), .B(n3742), .Z(n3687) );
  HS65_LH_NAND2X5 U6435 ( .A(n4820), .B(n4819), .Z(n4825) );
  HS65_LH_IVX2 U8214 ( .A(n4804), .Z(n4217) );
  HS65_LH_NAND3X3 U4770 ( .A(n5427), .B(n5426), .C(n5425), .Z(n5429) );
  HS65_LH_IVX7 U4402 ( .A(n5438), .Z(n5459) );
  HS65_LH_AOI21X2 U8320 ( .A(n4781), .B(n5063), .C(n4750), .Z(n4385) );
  HS65_LH_NAND2X4 U4848 ( .A(\lte_x_57/B[7] ), .B(n3742), .Z(n4214) );
  HS65_LH_NAND2X4 U4013 ( .A(n4214), .B(n4213), .Z(n4837) );
  HS65_LH_NAND2X7 U3956 ( .A(n3875), .B(n3874), .Z(n3876) );
  HS65_LH_OAI21X2 U3946 ( .A(n4794), .B(n2789), .C(n3379), .Z(n4795) );
  HS65_LH_NAND3X5 U3947 ( .A(n4973), .B(n4972), .C(n4971), .Z(n4978) );
  HS65_LH_NOR3X4 U3934 ( .A(n5062), .B(n4812), .C(n4284), .Z(n4309) );
  HS65_LL_AOI21X2 U3845 ( .A(n3081), .B(n3885), .C(n3080), .Z(n3082) );
  HS65_LH_NAND2X7 U6321 ( .A(n5433), .B(n4461), .Z(n3500) );
  HS65_LL_OAI12X2 U6266 ( .A(n3206), .B(n4643), .C(n3205), .Z(n3207) );
  HS65_LL_NOR2X2 U3925 ( .A(n5414), .B(n5413), .Z(n5423) );
  HS65_LH_CNIVX3 U8250 ( .A(n4742), .Z(n3337) );
  HS65_LL_OAI21X2 U4337 ( .A(n4084), .B(n2823), .C(n4083), .Z(n4085) );
  HS65_LH_IVX9 U3645 ( .A(n4105), .Z(n4711) );
  HS65_LL_AOI12X2 U8284 ( .A(n4525), .B(n4692), .C(n4524), .Z(n4528) );
  HS65_LL_NOR2X2 U6995 ( .A(n5499), .B(n4039), .Z(n4040) );
  HS65_LL_AOI22X1 U3835 ( .A(n4618), .B(n4831), .C(n4667), .D(n4617), .Z(n4627) );
  HS65_LH_IVX9 U3639 ( .A(n4667), .Z(n4744) );
  HS65_LH_NAND2X4 U3848 ( .A(n3314), .B(n4639), .Z(n3316) );
  HS65_LH_NAND2X4 U3847 ( .A(n4400), .B(n4639), .Z(n4402) );
  HS65_LH_NAND2X5 U4330 ( .A(n5492), .B(n4826), .Z(n4858) );
  HS65_LL_OAI12X2 U7717 ( .A(n5278), .B(n5277), .C(n5276), .Z(n5528) );
  HS65_LH_NAND2X7 U3679 ( .A(n4858), .B(n4857), .Z(n4869) );
  HS65_LH_NAND2X5 U6920 ( .A(n4774), .B(n4548), .Z(n4549) );
  HS65_LL_AOI21X2 U6139 ( .A(n7327), .B(n4307), .C(n4306), .Z(n8347) );
  HS65_LL_DFPQX9 clk_r_REG601_S6 ( .D(n3234), .CP(clk), .Q(n9012) );
  HS65_LL_DFPQNX18 clk_r_REG602_S6 ( .D(n2781), .CP(clk), .QN(n2782) );
  HS65_LL_IVX9 U3579 ( .A(n3236), .Z(n2712) );
  HS65_LH_IVX9 U3644 ( .A(\u_DataPath/cw_to_ex_i [2]), .Z(n5329) );
  HS65_LH_AOI21X2 U4094 ( .A(n8718), .B(n2712), .C(n3151), .Z(n3152) );
  HS65_LH_IVX9 U4082 ( .A(n3993), .Z(\add_x_50/A[19] ) );
  HS65_LL_CNIVX7 U6406 ( .A(n5211), .Z(n2789) );
  HS65_LL_NOR3X4 U4938 ( .A(n3038), .B(n2842), .C(n3037), .Z(n3039) );
  HS65_LH_IVX9 U5418 ( .A(n5203), .Z(n3078) );
  HS65_LH_AOI21X2 U3802 ( .A(\sub_x_51/A[21] ), .B(n5498), .C(n3489), .Z(n3492) );
  HS65_LH_IVX9 U7130 ( .A(n4147), .Z(n4411) );
  HS65_LH_IVX9 U8596 ( .A(n2825), .Z(\sub_x_51/A[22] ) );
  HS65_LH_IVX9 U6526 ( .A(n5190), .Z(n4622) );
  HS65_LL_OAI12X3 U6575 ( .A(n3165), .B(n8442), .C(n3164), .Z(n5252) );
  HS65_LH_OAI12X3 U5372 ( .A(n4272), .B(n4023), .C(n5108), .Z(n4239) );
  HS65_LH_AOI21X2 U4734 ( .A(n4168), .B(n4082), .C(n4081), .Z(n4083) );
  HS65_LH_AOI21X2 U8796 ( .A(n8713), .B(n9048), .C(n8773), .Z(n5847) );
  HS65_LH_AOI21X2 U8259 ( .A(n5507), .B(n5084), .C(n5506), .Z(n3913) );
  HS65_LH_AOI21X2 U7120 ( .A(n4781), .B(n5187), .C(n4750), .Z(n4438) );
  HS65_LH_AOI21X2 U5232 ( .A(n4543), .B(n4646), .C(n4542), .Z(n4544) );
  HS65_LH_AOI21X2 U7133 ( .A(n4781), .B(n5246), .C(n4750), .Z(n3546) );
  HS65_LL_AOI21X2 U6918 ( .A(n7327), .B(n4056), .C(n4055), .Z(n8351) );
  HS65_LL_AOI21X2 U5176 ( .A(n7327), .B(n4499), .C(n4498), .Z(n8331) );
  HS65_LL_AOI21X2 U6125 ( .A(n7327), .B(n3371), .C(n3370), .Z(n8329) );
  HS65_LH_DFPRQX9 clk_r_REG857_S4 ( .D(n6725), .CP(net3007), .RN(n9555), .Q(
        n9472) );
  HS65_LL_AOI21X2 U3371 ( .A(n4774), .B(n7316), .C(n4700), .Z(n8337) );
  HS65_LH_AOI21X2 U3372 ( .A(n4294), .B(n5504), .C(n4293), .Z(n4298) );
  HS65_LH_IVX9 U3376 ( .A(n4871), .Z(n5497) );
  HS65_LL_NOR4ABX2 U3379 ( .A(n8772), .B(n8729), .C(n8569), .D(n8585), .Z(
        n8001) );
  HS65_LL_MX41X4 U3381 ( .D0(n8770), .S0(n9482), .D1(n8623), .S1(n9496), .D2(
        n9503), .S2(n8767), .D3(n9081), .S3(n9489), .Z(
        \u_DataPath/from_mem_data_out_i [6]) );
  HS65_LH_NAND2X2 U3384 ( .A(\lte_x_57/B[29] ), .B(n4208), .Z(n3396) );
  HS65_LL_IVX9 U3385 ( .A(n2830), .Z(n4208) );
  HS65_LL_OAI21X3 U3392 ( .A(n3316), .B(n4714), .C(n3315), .Z(n3317) );
  HS65_LH_AOI22X1 U3394 ( .A(n4673), .B(n4742), .C(n4225), .D(n4672), .Z(n4675) );
  HS65_LH_AOI21X2 U3402 ( .A(n4225), .B(n3824), .C(n5208), .Z(n3832) );
  HS65_LH_NAND3X2 U3405 ( .A(n4796), .B(n4411), .C(n4225), .Z(n3294) );
  HS65_LH_NAND2X2 U3407 ( .A(n4225), .B(n4290), .Z(n3493) );
  HS65_LL_NOR2AX3 U3408 ( .A(n4225), .B(n4224), .Z(n4226) );
  HS65_LL_MUX21I1X3 U3411 ( .D0(n2773), .D1(n8730), .S0(
        \u_DataPath/cw_to_ex_i [14]), .Z(n5196) );
  HS65_LL_IVX9 U3413 ( .A(n2772), .Z(n2797) );
  HS65_LLS_XNOR2X3 U3417 ( .A(n4429), .B(n4428), .Z(n4457) );
  HS65_LL_CNIVX3 U3420 ( .A(n5201), .Z(n3072) );
  HS65_LH_CBI4I6X2 U3427 ( .A(n3231), .B(n3230), .C(n4842), .D(n3229), .Z(
        n3232) );
  HS65_LL_AO12X4 U3428 ( .A(n4843), .B(n4842), .C(n4841), .Z(n4854) );
  HS65_LH_NOR2AX3 U3432 ( .A(n4842), .B(n4674), .Z(n4618) );
  HS65_LL_AO12X4 U3436 ( .A(n8698), .B(n2798), .C(n3068), .Z(n2839) );
  HS65_LL_NAND4ABX3 U3437 ( .A(n8349), .B(n4361), .C(n8347), .D(n4360), .Z(
        n4362) );
  HS65_LL_AOI21X3 U3438 ( .A(n7327), .B(n4236), .C(n4235), .Z(n8342) );
  HS65_LL_AOI21X3 U3439 ( .A(n5492), .B(n3505), .C(n3504), .Z(n8355) );
  HS65_LL_NAND2X2 U3444 ( .A(n3503), .B(n3502), .Z(n3504) );
  HS65_LL_AOI21X2 U3457 ( .A(n4411), .B(n3605), .C(n3604), .Z(n3623) );
  HS65_LL_NOR2X2 U3458 ( .A(n4167), .B(n4166), .Z(n4183) );
  HS65_LL_NOR3X1 U3485 ( .A(n3305), .B(n3304), .C(n3303), .Z(n3306) );
  HS65_LL_AOI21X2 U3492 ( .A(\lte_x_57/B[29] ), .B(n4508), .C(n4507), .Z(n4518) );
  HS65_LH_OAI21X2 U3502 ( .A(n4794), .B(n3204), .C(n4501), .Z(n4508) );
  HS65_LL_AOI211X1 U3517 ( .A(n4667), .B(n4742), .C(n3548), .D(n3547), .Z(
        n3549) );
  HS65_LL_AOI12X2 U3531 ( .A(n5353), .B(n5352), .C(n5351), .Z(n5358) );
  HS65_LL_NOR2X6 U3534 ( .A(n4147), .B(n2776), .Z(n4667) );
  HS65_LH_NOR2X6 U3555 ( .A(n3325), .B(n3324), .Z(n4746) );
  HS65_LH_NOR2X3 U3590 ( .A(n5347), .B(n5341), .Z(n5413) );
  HS65_LL_AOI12X3 U3598 ( .A(n4216), .B(n3253), .C(n3252), .Z(n3760) );
  HS65_LH_IVX9 U3610 ( .A(n4440), .Z(n4671) );
  HS65_LH_NOR3X4 U3612 ( .A(n5281), .B(n5280), .C(n5318), .Z(n5325) );
  HS65_LL_NAND2X4 U3620 ( .A(n3273), .B(n4604), .Z(n4682) );
  HS65_LH_NOR2X3 U3632 ( .A(n5211), .B(n4189), .Z(n5342) );
  HS65_LH_CNIVX3 U3642 ( .A(n5043), .Z(n5420) );
  HS65_LH_IVX7 U3654 ( .A(n5233), .Z(n4091) );
  HS65_LH_NAND3X3 U3695 ( .A(n5227), .B(n4876), .C(n4895), .Z(n4899) );
  HS65_LL_OAI12X3 U3722 ( .A(n3842), .B(n3765), .C(n3767), .Z(n4862) );
  HS65_LH_NAND2X7 U3723 ( .A(\sub_x_51/A[16] ), .B(n4796), .Z(n3646) );
  HS65_LH_NAND2X5 U3731 ( .A(n3993), .B(n5246), .Z(n5003) );
  HS65_LH_OAI12X3 U3735 ( .A(n5396), .B(n3886), .C(n5234), .Z(n5235) );
  HS65_LL_NAND2X7 U3739 ( .A(n3587), .B(n3241), .Z(n4738) );
  HS65_LL_CNIVX3 U3747 ( .A(n4653), .Z(n4620) );
  HS65_LH_NOR2X5 U3753 ( .A(n3054), .B(n5203), .Z(n5371) );
  HS65_LH_NAND2X7 U3766 ( .A(\sub_x_51/A[18] ), .B(n5063), .Z(n4374) );
  HS65_LH_AO22X9 U3780 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][0] ), .B(n9202), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][0] ), .D(
        n9201), .Z(n7291) );
  HS65_LL_CNIVX3 U3813 ( .A(n5252), .Z(n3195) );
  HS65_LH_NAND2X7 U3830 ( .A(\u_DataPath/cw_to_ex_i [1]), .B(n5329), .Z(n3240)
         );
  HS65_LL_OAI211X3 U3899 ( .A(n8816), .B(n7986), .C(n7985), .D(n7984), .Z(
        \u_DataPath/cw_to_ex_i [3]) );
  HS65_LH_NAND2X7 U3902 ( .A(n9134), .B(\u_DataPath/cw_to_ex_i [14]), .Z(n2992) );
  HS65_LH_NOR2X6 U3917 ( .A(n6483), .B(n6482), .Z(n6484) );
  HS65_LL_NAND3X13 U3932 ( .A(n9373), .B(n9374), .C(n8362), .Z(
        \u_DataPath/cw_to_ex_i [14]) );
  HS65_LL_NOR4ABX4 U4008 ( .A(n4365), .B(n4364), .C(n4363), .D(n4362), .Z(
        n8357) );
  HS65_LL_NAND2X2 U4039 ( .A(n8342), .B(n8350), .Z(n4361) );
  HS65_LL_NAND3X3 U4050 ( .A(n3623), .B(n3622), .C(n3621), .Z(n8346) );
  HS65_LL_NAND2X4 U4090 ( .A(n3938), .B(n3937), .Z(n8345) );
  HS65_LL_NOR2AX3 U4092 ( .A(n5523), .B(n5522), .Z(n5524) );
  HS65_LL_NOR2X2 U4140 ( .A(n4760), .B(n4759), .Z(n4761) );
  HS65_LL_IVX2 U4144 ( .A(n3603), .Z(n3604) );
  HS65_LL_NAND4ABX3 U4189 ( .A(n5521), .B(n5520), .C(n5519), .D(n5518), .Z(
        n5522) );
  HS65_LL_NAND3X2 U4203 ( .A(n4299), .B(n4298), .C(n4297), .Z(n4300) );
  HS65_LH_AOI21X2 U4222 ( .A(n5484), .B(n5483), .C(n5482), .Z(n5523) );
  HS65_LL_OAI112X1 U4296 ( .A(n4476), .B(n2776), .C(n4475), .D(n4474), .Z(
        n4485) );
  HS65_LL_AOI21X2 U4298 ( .A(n5517), .B(n5516), .C(n5515), .Z(n5518) );
  HS65_LL_AOI21X2 U4302 ( .A(n5171), .B(\u_DataPath/cw_to_ex_i [2]), .C(n5170), 
        .Z(n5172) );
  HS65_LL_NAND3X2 U4356 ( .A(n4287), .B(n4286), .C(n4285), .Z(n4288) );
  HS65_LL_AOI12X2 U4369 ( .A(n5517), .B(n4984), .C(n3470), .Z(n3473) );
  HS65_LH_OAI12X3 U4371 ( .A(n5468), .B(n5467), .C(n5466), .Z(n5469) );
  HS65_LH_AOI22X3 U4385 ( .A(n5517), .B(n4974), .C(n5510), .D(n4609), .Z(n4251) );
  HS65_LL_OAI112X1 U4390 ( .A(n4623), .B(n4321), .C(n3233), .D(n3232), .Z(
        n3605) );
  HS65_LH_AOI21X2 U4400 ( .A(n4836), .B(n5483), .C(n4296), .Z(n4297) );
  HS65_LH_IVX4 U4411 ( .A(n4748), .Z(n4749) );
  HS65_LH_NAND3X5 U4425 ( .A(n4130), .B(n4129), .C(n4471), .Z(n4131) );
  HS65_LH_IVX7 U4454 ( .A(n3390), .Z(n4441) );
  HS65_LH_NOR2X3 U4458 ( .A(n5290), .B(n5002), .Z(n5052) );
  HS65_LH_NOR2X5 U4470 ( .A(n4523), .B(n4682), .Z(n4525) );
  HS65_LH_NOR2X6 U4486 ( .A(n3691), .B(n3690), .Z(n4333) );
  HS65_LL_NAND2X4 U4495 ( .A(n3720), .B(n3719), .Z(n4844) );
  HS65_LH_CNIVX3 U4504 ( .A(n4427), .Z(n3650) );
  HS65_LL_OAI12X2 U4509 ( .A(n4592), .B(n3312), .C(n4594), .Z(n3313) );
  HS65_LH_CNIVX3 U4515 ( .A(n3969), .Z(n3974) );
  HS65_LL_NAND2X4 U4517 ( .A(n3492), .B(n3491), .Z(n4290) );
  HS65_LHS_XNOR2X6 U4523 ( .A(n5490), .B(n3785), .Z(n9505) );
  HS65_LL_NAND2X4 U4556 ( .A(n3926), .B(n3925), .Z(n4742) );
  HS65_LL_NOR2X3 U4566 ( .A(n3416), .B(n3419), .Z(n4604) );
  HS65_LH_NAND3X5 U4578 ( .A(n4944), .B(n4943), .C(n4942), .Z(n5166) );
  HS65_LH_IVX9 U4670 ( .A(n4613), .Z(n4673) );
  HS65_LH_NOR2X5 U4675 ( .A(n4032), .B(n3322), .Z(n4212) );
  HS65_LH_IVX4 U4689 ( .A(n4270), .Z(n4271) );
  HS65_LH_CNIVX3 U4698 ( .A(n4784), .Z(n3720) );
  HS65_LH_NOR2X5 U4699 ( .A(n5092), .B(n4192), .Z(n5415) );
  HS65_LH_AOI22X3 U4708 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][1] ), .B(n9473), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][1] ), .D(
        n9474), .Z(n6239) );
  HS65_LL_NAND2X5 U4739 ( .A(n3284), .B(n3301), .Z(n4794) );
  HS65_LH_OAI12X3 U4751 ( .A(n8886), .B(n5878), .C(n9107), .Z(n5880) );
  HS65_LH_IVX9 U4762 ( .A(n3962), .Z(\lte_x_57/B[15] ) );
  HS65_LH_OR2X9 U4789 ( .A(n8407), .B(n2794), .Z(n9543) );
  HS65_LH_OAI12X3 U4854 ( .A(n9049), .B(n5894), .C(n8777), .Z(n5813) );
  HS65_LH_NOR2X5 U4858 ( .A(n9408), .B(n7641), .Z(n7425) );
  HS65_LH_NOR2X5 U4913 ( .A(n8624), .B(n2772), .Z(n8391) );
  HS65_LH_NAND2X5 U4919 ( .A(n2947), .B(n2800), .Z(n8383) );
  HS65_LH_NOR2X5 U4920 ( .A(\u_DataPath/dataOut_exe_i [30]), .B(n3980), .Z(
        n2919) );
  HS65_LL_OAI112X4 U4962 ( .A(n8800), .B(n8002), .C(n8001), .D(n8000), .Z(
        \u_DataPath/cw_to_ex_i [0]) );
  HS65_LL_OAI12X3 U4963 ( .A(n9421), .B(n7986), .C(n7977), .Z(
        \u_DataPath/cw_to_ex_i [4]) );
  HS65_LH_OAI12X3 U4971 ( .A(n8980), .B(n5633), .C(n9027), .Z(n5612) );
  HS65_LH_IVX4 U4985 ( .A(n9330), .Z(n3008) );
  HS65_LL_AO312X9 U5016 ( .A(n9177), .B(n9444), .C(n9504), .D(n9023), .E(n9278), .F(n8781), .Z(\u_DataPath/dataOut_exe_i [1]) );
  HS65_LH_NAND3X5 U5032 ( .A(n8900), .B(n9310), .C(n8821), .Z(n7971) );
  HS65_LH_OAI12X3 U5042 ( .A(n8998), .B(n8777), .C(n8708), .Z(n5746) );
  HS65_LL_NAND4ABX6 U5160 ( .A(n5182), .B(n5181), .C(n8337), .D(n5180), .Z(
        n7664) );
  HS65_LL_NOR3AX4 U5162 ( .A(n3939), .B(n8345), .C(n8346), .Z(n4102) );
  HS65_LL_NAND3AX3 U5166 ( .A(n4539), .B(n4538), .C(n4537), .Z(n4550) );
  HS65_LL_NAND2AX4 U5168 ( .A(n3879), .B(n3878), .Z(n3880) );
  HS65_LL_NAND2AX4 U5178 ( .A(n4869), .B(n4868), .Z(n8322) );
  HS65_LLS_XNOR2X3 U5179 ( .A(n4531), .B(n4530), .Z(n4532) );
  HS65_LL_AOI211X3 U5180 ( .A(n4774), .B(n3428), .C(n3427), .D(n3426), .Z(
        n8330) );
  HS65_LL_OAI21X2 U5184 ( .A(n4305), .B(n9544), .C(n4303), .Z(n4306) );
  HS65_LL_NOR2AX3 U5186 ( .A(n3751), .B(n3750), .Z(n3752) );
  HS65_LHS_XNOR2X6 U5192 ( .A(n4109), .B(n4108), .Z(n4145) );
  HS65_LL_NAND2X2 U5199 ( .A(n4518), .B(n4517), .Z(n4539) );
  HS65_LL_NAND3X2 U5205 ( .A(n4165), .B(n4164), .C(n4163), .Z(n4166) );
  HS65_LL_NAND2AX4 U5208 ( .A(n3840), .B(n3839), .Z(n8340) );
  HS65_LL_AOI21X2 U5215 ( .A(n5517), .B(n4975), .C(n4288), .Z(n4299) );
  HS65_LL_NAND3X2 U5221 ( .A(n5514), .B(n5513), .C(n5512), .Z(n5515) );
  HS65_LLS_XOR2X3 U5222 ( .A(n4695), .B(n3660), .Z(n3661) );
  HS65_LL_NAND2X2 U5225 ( .A(n4065), .B(n4064), .Z(n4535) );
  HS65_LL_AOI12X2 U5229 ( .A(n3805), .B(n3804), .C(n4871), .Z(n3812) );
  HS65_LH_NOR2AX3 U5230 ( .A(n4470), .B(n4469), .Z(n4475) );
  HS65_LHS_XNOR2X6 U5269 ( .A(n4050), .B(n4049), .Z(n4051) );
  HS65_LL_AOI21X2 U5287 ( .A(n5517), .B(n4986), .C(n4131), .Z(n4132) );
  HS65_LH_NAND2X4 U5289 ( .A(n5510), .B(n4789), .Z(n4790) );
  HS65_LH_OAI21X3 U5297 ( .A(n3913), .B(n3962), .C(n3912), .Z(n3914) );
  HS65_LH_NAND2X4 U5305 ( .A(n4175), .B(n4090), .Z(n4094) );
  HS65_LH_OAI21X3 U5310 ( .A(n4613), .B(n4514), .C(n3399), .Z(n4045) );
  HS65_LL_OAI12X2 U5321 ( .A(n4662), .B(n5499), .C(n4655), .Z(n4656) );
  HS65_LL_OAI12X2 U5330 ( .A(n4784), .B(n4783), .C(n4782), .Z(n4785) );
  HS65_LH_AOI31X3 U5337 ( .A(n4662), .B(n4661), .C(n4660), .D(n4659), .Z(n4663) );
  HS65_LL_AOI12X2 U5340 ( .A(n4433), .B(n4432), .C(n4503), .Z(n4476) );
  HS65_LL_NAND2X2 U5342 ( .A(n4673), .B(n4843), .Z(n4245) );
  HS65_LL_NAND3X3 U5345 ( .A(n3401), .B(n3735), .C(n3400), .Z(n4479) );
  HS65_LH_CBI4I1X5 U5358 ( .A(n3592), .B(n3591), .C(n4812), .D(n3590), .Z(
        n4843) );
  HS65_LHS_XNOR2X6 U5370 ( .A(n3779), .B(n3778), .Z(n9542) );
  HS65_LH_NAND2X4 U5371 ( .A(n5259), .B(n3373), .Z(n3378) );
  HS65_LL_OR2X9 U5390 ( .A(n5092), .B(n5211), .Z(n4321) );
  HS65_LL_OAI12X2 U5394 ( .A(n4802), .B(n4799), .C(n4801), .Z(n3252) );
  HS65_LL_NAND2X5 U5421 ( .A(n3239), .B(n5211), .Z(n4284) );
  HS65_LH_AOI21X2 U5437 ( .A(\lte_x_57/B[11] ), .B(n3826), .C(n4313), .Z(n3925) );
  HS65_LH_OAI12X3 U5453 ( .A(n4552), .B(n3372), .C(n5259), .Z(n4595) );
  HS65_LH_IVX4 U5456 ( .A(n3782), .Z(n3783) );
  HS65_LH_NOR2X3 U5490 ( .A(n3951), .B(n3338), .Z(n4775) );
  HS65_LH_NAND2X5 U5491 ( .A(\lte_x_57/B[4] ), .B(n3241), .Z(n3842) );
  HS65_LL_NAND2X4 U5496 ( .A(\add_x_50/A[23] ), .B(n3195), .Z(n4703) );
  HS65_LL_NAND2AX14 U5501 ( .A(n5062), .B(n2802), .Z(n4846) );
  HS65_LL_OR2X9 U5516 ( .A(n2991), .B(n7670), .Z(n2844) );
  HS65_LL_NOR2X6 U5539 ( .A(n3015), .B(n3014), .Z(\lte_x_57/B[10] ) );
  HS65_LH_OAI21X3 U5549 ( .A(n8652), .B(n2772), .C(n2920), .Z(n8450) );
  HS65_LH_OAI21X3 U5550 ( .A(n9330), .B(n3178), .C(n3004), .Z(n3005) );
  HS65_LH_NAND2X4 U5563 ( .A(n8701), .B(n2798), .Z(n8419) );
  HS65_LHS_XNOR2X6 U5608 ( .A(n8913), .B(n5904), .Z(
        \u_DataPath/u_execute/resAdd1_i [7]) );
  HS65_LHS_XNOR2X6 U5660 ( .A(n8819), .B(n8813), .Z(n7209) );
  HS65_LL_MUXI21X2 U5684 ( .D0(n8794), .D1(\u_DataPath/from_mem_data_out_i [6]), .S0(n9415), .Z(n8245) );
  HS65_LHS_XNOR2X6 U5752 ( .A(n9167), .B(n9061), .Z(n6482) );
  HS65_LL_OAI12X3 U5833 ( .A(n9044), .B(n8753), .C(n8593), .Z(
        \u_DataPath/dataOut_exe_i [20]) );
  HS65_LL_OAI12X3 U5912 ( .A(n9044), .B(n8749), .C(n8599), .Z(
        \u_DataPath/dataOut_exe_i [27]) );
  HS65_LH_OAI12X6 U5916 ( .A(n9044), .B(n8763), .C(n9077), .Z(
        \u_DataPath/dataOut_exe_i [4]) );
  HS65_LH_IVX2 U5924 ( .A(n5343), .Z(n5041) );
  HS65_LH_IVX2 U5925 ( .A(n4118), .Z(n3595) );
  HS65_LH_OR2X4 U5926 ( .A(n2854), .B(n3595), .Z(n3596) );
  HS65_LH_NAND2X2 U5975 ( .A(n3090), .B(n8389), .Z(n2925) );
  HS65_LH_NAND2X2 U6114 ( .A(\lte_x_57/B[10] ), .B(n4796), .Z(n4202) );
  HS65_LH_OAI21X2 U6120 ( .A(n5108), .B(n5107), .C(n5426), .Z(n5113) );
  HS65_LL_NOR2X2 U6123 ( .A(n4701), .B(n5132), .Z(n5134) );
  HS65_LH_IVX2 U6128 ( .A(n3900), .Z(n3902) );
  HS65_LH_NOR2X2 U6137 ( .A(\sub_x_51/A[5] ), .B(n2787), .Z(n5218) );
  HS65_LH_AND3X4 U6140 ( .A(n5053), .B(n5052), .C(n5461), .Z(n2834) );
  HS65_LH_OAI31X1 U6146 ( .A(n4913), .B(n5367), .C(n5296), .D(n5003), .Z(n4916) );
  HS65_LH_NAND2X2 U6148 ( .A(n5356), .B(n5337), .Z(n3955) );
  HS65_LHS_XNOR2X3 U6154 ( .A(n4803), .B(n4218), .Z(n9540) );
  HS65_LH_AOI22X1 U6155 ( .A(n5505), .B(n4828), .C(n5484), .D(n4832), .Z(n4244) );
  HS65_LH_NOR2X2 U6162 ( .A(n5078), .B(n5200), .Z(n5231) );
  HS65_LH_OAI21X2 U6163 ( .A(n5106), .B(n5105), .C(n5104), .Z(n5123) );
  HS65_LH_IVX2 U6165 ( .A(n4931), .Z(n4935) );
  HS65_LL_NOR4ABX4 U6167 ( .A(n8355), .B(n4102), .C(n8339), .D(n4101), .Z(
        n4364) );
  HS65_LH_AOI21X2 U6170 ( .A(n4781), .B(n5072), .C(n4750), .Z(n3382) );
  HS65_LL_OAI12X2 U6176 ( .A(n3362), .B(n4695), .C(n3361), .Z(n3363) );
  HS65_LH_AOI22X1 U6181 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][2] ), .B(n9199), 
        .C(n9198), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][2] ), .Z(n6144)
         );
  HS65_LH_AOI22X1 U6183 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][7] ), .B(n8938), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][7] ), .D(n9264), .Z(n6467) );
  HS65_LH_AOI22X1 U6184 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][13] ), .B(n9247), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][13] ), .D(
        n9227), .Z(n7024) );
  HS65_LH_AOI22X1 U6185 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][3] ), .B(n9199), 
        .C(n9198), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][3] ), .Z(n6106)
         );
  HS65_LH_AO22X4 U6186 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][11] ), .B(n9254), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][11] ), .D(
        n9244), .Z(n6815) );
  HS65_LH_AO22X4 U6190 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][26] ), .B(n9470), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][26] ), .D(
        n9164), .Z(n6946) );
  HS65_LH_AOI22X1 U6200 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][8] ), .B(n9242), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][8] ), .D(n8861), .Z(n6853) );
  HS65_LH_AOI22X1 U6201 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][6] ), .B(n9242), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][6] ), .D(n8861), .Z(n6833) );
  HS65_LH_AOI22X1 U6203 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][6] ), .B(n9199), 
        .C(n9198), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][6] ), .Z(n6823)
         );
  HS65_LH_AO22X4 U6204 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][19] ), .B(n9469), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][19] ), .D(
        n8853), .Z(n6292) );
  HS65_LH_AO22X4 U6212 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][12] ), .B(n9261), 
        .C(n9263), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][12] ), .Z(n7147)
         );
  HS65_LH_AO22X4 U6218 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][8] ), .B(n8939), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][8] ), .D(
        n9186), .Z(n6654) );
  HS65_LH_AOI22X1 U6219 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][24] ), .B(n8851), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][24] ), .D(
        n9264), .Z(n6274) );
  HS65_LH_AO22X4 U6226 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][17] ), .B(n9261), 
        .C(n9263), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][17] ), .Z(n5956)
         );
  HS65_LH_AO22X4 U6240 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][10] ), .B(n9364), 
        .C(n9253), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][10] ), .Z(n7041)
         );
  HS65_LH_AOI22X1 U6243 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][1] ), .B(n9259), 
        .C(n9256), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][1] ), .Z(n7247)
         );
  HS65_LH_AOI22X1 U6249 ( .A(n9207), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][19] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][19] ), .D(n9266), 
        .Z(n6768) );
  HS65_LH_AOI22X1 U6253 ( .A(n9207), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][7] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][7] ), .D(n9266), 
        .Z(n6047) );
  HS65_LH_AO22X4 U6260 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][29] ), .B(n9251), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][29] ), .D(
        n9186), .Z(n6921) );
  HS65_LH_AOI22X1 U6264 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][14] ), .B(n8938), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][14] ), .D(
        n9264), .Z(n6871) );
  HS65_LH_AOI22X1 U6278 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][25] ), .B(n8938), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][25] ), .D(
        n9264), .Z(n6961) );
  HS65_LH_AO22X4 U6287 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][12] ), .B(n9470), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][12] ), .D(
        n9267), .Z(n6698) );
  HS65_LH_AO22X4 U6288 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][15] ), .B(n9470), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][15] ), .D(
        n9267), .Z(n6898) );
  HS65_LH_AOI22X1 U6289 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][21] ), .B(n9159), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][21] ), .D(
        n9265), .Z(n6007) );
  HS65_LH_AOI22X1 U6294 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][21] ), .B(n9208), 
        .C(n9100), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][21] ), .Z(n5997)
         );
  HS65_LH_AOI22X1 U6299 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][9] ), .B(n9255), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][9] ), .D(
        n9195), .Z(n6980) );
  HS65_LH_AO22X4 U6303 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][20] ), .B(n8858), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][20] ), .D(
        n9468), .Z(n6584) );
  HS65_LH_AO22X4 U6304 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][20] ), .B(n9204), 
        .C(n9203), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][20] ), .Z(n7096)
         );
  HS65_LH_AOI22X1 U6305 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][5] ), .B(n8950), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][5] ), .D(
        n8855), .Z(n6630) );
  HS65_LH_AOI22X1 U6306 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][10] ), .B(n9188), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][10] ), .D(
        n9190), .Z(n6710) );
  HS65_LH_AOI22X1 U6310 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][6] ), .B(n9188), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][6] ), .D(
        n9190), .Z(n6734) );
  HS65_LH_AO22X4 U6312 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][22] ), .B(n9469), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][22] ), .D(
        n9475), .Z(n6548) );
  HS65_LH_AO22X4 U6316 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][15] ), .B(n9261), 
        .C(n9101), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][15] ), .Z(n7269)
         );
  HS65_LH_AO22X4 U6318 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][28] ), .B(n9251), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][28] ), .D(
        n9155), .Z(n6533) );
  HS65_LH_AO22X4 U6345 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][30] ), .B(n9251), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][30] ), .D(
        n9155), .Z(n6573) );
  HS65_LH_AO22X4 U6347 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][31] ), .B(n9251), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][31] ), .D(
        n9155), .Z(n6613) );
  HS65_LH_AOI22X1 U6362 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][5] ), .B(n9199), 
        .C(n9198), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][5] ), .Z(n7078)
         );
  HS65_LH_AOI22X1 U6364 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][9] ), .B(n9199), 
        .C(n9198), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][9] ), .Z(n7058)
         );
  HS65_LH_AO22X4 U6369 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][29] ), .B(n9261), 
        .C(n9263), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][29] ), .Z(n7552)
         );
  HS65_LH_AOI22X1 U6374 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][27] ), .B(n9208), 
        .C(n9100), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][27] ), .Z(n7159)
         );
  HS65_LH_AO22X4 U6396 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][23] ), .B(n9261), 
        .C(n9263), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][23] ), .Z(n7127)
         );
  HS65_LH_AO22X4 U6399 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][28] ), .B(n9363), 
        .C(n9257), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][28] ), .Z(n7592)
         );
  HS65_LH_AO22X4 U6401 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][30] ), .B(n9152), 
        .C(n9257), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][30] ), .Z(n7538)
         );
  HS65_LH_AO22X4 U6404 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][26] ), .B(n9261), 
        .C(n9263), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][26] ), .Z(n6792)
         );
  HS65_LH_AOI22X1 U6429 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][13] ), .B(n8851), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][13] ), .D(
        n9264), .Z(n6406) );
  HS65_LH_AOI22X1 U6432 ( .A(n9207), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][31] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][31] ), .D(n9266), 
        .Z(n7512) );
  HS65_LH_AOI22X1 U6447 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][21] ), .B(n8851), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][21] ), .D(
        n9264), .Z(n6386) );
  HS65_LH_AOI22X1 U6450 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][18] ), .B(n9250), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][18] ), .D(
        n9265), .Z(n7231) );
  HS65_LH_AOI22X1 U6458 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][24] ), .B(n9250), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][24] ), .D(
        n9265), .Z(n5987) );
  HS65_LH_AOI22X1 U6469 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][24] ), .B(n9208), 
        .C(n9100), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][24] ), .Z(n5975)
         );
  HS65_LH_AOI22X1 U6478 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][16] ), .B(n9208), 
        .C(n9100), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][16] ), .Z(n6063)
         );
  HS65_LH_AOI22X1 U6483 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][17] ), .B(n8851), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][17] ), .D(
        n9264), .Z(n6366) );
  HS65_LH_AOI22X1 U6487 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][23] ), .B(n9226), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][23] ), .D(
        n9193), .Z(n6350) );
  HS65_LH_AOI22X1 U6491 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][11] ), .B(n9226), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][11] ), .D(
        n9193), .Z(n6513) );
  HS65_LH_AOI22X1 U6509 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][1] ), .B(n8851), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][1] ), .D(n9264), .Z(n6247) );
  HS65_LH_AO22X4 U6512 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][4] ), .B(n9472), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][4] ), .D(
        n9468), .Z(n6418) );
  HS65_LH_AO22X4 U6520 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][16] ), .B(n9473), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][16] ), .D(
        n9474), .Z(n6165) );
  HS65_LH_AOI22X1 U6539 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][27] ), .B(n9191), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][27] ), .D(
        n9471), .Z(n6316) );
  HS65_LH_AOI22X1 U6563 ( .A(n9207), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][4] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][4] ), .D(n9266), 
        .Z(n6025) );
  HS65_LH_AO22X4 U6566 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][2] ), .B(n9154), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][2] ), .D(
        n9194), .Z(n6221) );
  HS65_LH_AO22X4 U6568 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][3] ), .B(n9010), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][3] ), .D(n8849), .Z(n6452) );
  HS65_LH_AOI22X1 U6578 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][0] ), .B(n9226), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][0] ), .D(n9193), .Z(n6210) );
  HS65_LH_AOI22X1 U6590 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][18] ), .B(n8938), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][18] ), .D(
        n9264), .Z(n6673) );
  HS65_LH_AO22X4 U6591 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][22] ), .B(n9363), 
        .C(n9097), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][22] ), .Z(n7191)
         );
  HS65_LH_AOI22X1 U6592 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][25] ), .B(n9250), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][25] ), .D(
        n9265), .Z(n7489) );
  HS65_LH_AOI22X1 U6597 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][14] ), .B(n9242), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][14] ), .D(
        n9166), .Z(n6092) );
  HS65_LHS_XOR2X3 U6623 ( .A(n3103), .B(n3106), .Z(n4970) );
  HS65_LHS_XOR2X3 U6639 ( .A(\lte_x_57/B[28] ), .B(n4902), .Z(n4993) );
  HS65_LL_NAND3X2 U6648 ( .A(n9362), .B(n2989), .C(n9103), .Z(n3028) );
  HS65_LL_NAND2X2 U6658 ( .A(n8157), .B(n2961), .Z(n5183) );
  HS65_LH_AOI21X2 U6671 ( .A(n8751), .B(n2710), .C(n3116), .Z(n3118) );
  HS65_LL_MUXI21X2 U6692 ( .D0(n9289), .D1(n2941), .S0(n9415), .Z(n8158) );
  HS65_LHS_XOR2X3 U6696 ( .A(n8991), .B(n5758), .Z(
        \u_DataPath/u_execute/resAdd1_i [31]) );
  HS65_LL_AOI112X1 U6704 ( .A(n8821), .B(n9089), .C(n8731), .D(n8602), .Z(
        n8002) );
  HS65_LL_AOI22X1 U6706 ( .A(n8942), .B(n9252), .C(n9278), .D(n8873), .Z(n8296) );
  HS65_LL_NAND2X4 U6717 ( .A(n3663), .B(n3662), .Z(n8352) );
  HS65_LL_AOI21X4 U6889 ( .A(n7327), .B(n3881), .C(n3880), .Z(n8341) );
  HS65_LH_AO22X4 U6890 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][4] ), .B(n9202), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][4] ), .D(
        n9201), .Z(n6030) );
  HS65_LH_AO22X4 U6897 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][5] ), .B(n9202), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][5] ), .D(
        n9201), .Z(n7086) );
  HS65_LH_AO22X4 U6898 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][15] ), .B(n9202), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][15] ), .D(
        n9201), .Z(n7268) );
  HS65_LH_AO22X4 U6899 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][26] ), .B(n9202), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][26] ), .D(
        n9201), .Z(n6791) );
  HS65_LH_AO22X4 U6900 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][23] ), .B(n9202), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][23] ), .D(
        n9201), .Z(n7126) );
  HS65_LH_AO22X4 U6901 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][9] ), .B(n9202), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][9] ), .D(
        n9201), .Z(n7066) );
  HS65_LH_AO22X4 U6902 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][27] ), .B(n9202), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][27] ), .D(
        n9201), .Z(n7166) );
  HS65_LH_AO22X4 U6903 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][20] ), .B(n9202), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][20] ), .D(
        n9201), .Z(n7106) );
  HS65_LH_AO22X4 U6905 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][22] ), .B(n9202), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][22] ), .D(
        n9201), .Z(n7186) );
  HS65_LH_AO22X4 U6906 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][11] ), .B(n9202), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][11] ), .D(
        n9201), .Z(n6811) );
  HS65_LH_AO22X4 U6911 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][6] ), .B(n9202), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][6] ), .D(
        n9201), .Z(n6831) );
  HS65_LH_AO22X4 U6916 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][8] ), .B(n9202), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][8] ), .D(
        n9201), .Z(n6851) );
  HS65_LH_AO22X4 U6925 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][3] ), .B(n9202), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][3] ), .D(
        n9201), .Z(n6125) );
  HS65_LH_AO22X4 U6929 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][12] ), .B(n9202), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][12] ), .D(
        n9201), .Z(n7146) );
  HS65_LH_AO22X4 U6934 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][2] ), .B(n9202), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][2] ), .D(
        n9201), .Z(n6152) );
  HS65_LH_AO22X4 U6940 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][8] ), .B(n9472), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][8] ), .D(
        n9468), .Z(n6645) );
  HS65_LH_AO22X4 U6942 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][7] ), .B(n9472), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][7] ), .D(
        n9468), .Z(n6459) );
  HS65_LH_AO22X4 U6946 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][24] ), .B(n9472), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][24] ), .D(
        n8857), .Z(n6261) );
  HS65_LH_AO22X4 U6953 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][19] ), .B(n9472), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][19] ), .D(
        n8857), .Z(n6288) );
  HS65_LH_AO22X4 U6955 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][18] ), .B(n9472), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][18] ), .D(
        n9468), .Z(n6665) );
  HS65_LH_AO22X4 U6965 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][8] ), .B(n9473), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][8] ), .D(
        n9474), .Z(n6644) );
  HS65_LH_AO22X4 U6968 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][7] ), .B(n9473), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][7] ), .D(
        n9474), .Z(n6458) );
  HS65_LH_AO22X4 U6973 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][24] ), .B(n9473), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][24] ), .D(
        n9474), .Z(n6260) );
  HS65_LH_AO22X4 U6976 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][19] ), .B(n9473), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][19] ), .D(
        n9474), .Z(n6287) );
  HS65_LH_AO22X4 U6988 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][18] ), .B(n9473), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][18] ), .D(
        n9474), .Z(n6664) );
  HS65_LL_NAND2AX4 U6999 ( .A(n4653), .B(n3588), .Z(n4784) );
  HS65_LL_NAND3X2 U7010 ( .A(n9089), .B(n8800), .C(n8821), .Z(n7986) );
  HS65_LLS_XNOR2X3 U7014 ( .A(n4651), .B(n4650), .Z(n7316) );
  HS65_LL_MX41X4 U7022 ( .D0(n8623), .S0(n9491), .D1(n8770), .S1(n9477), .D2(
        n8767), .S2(n9498), .D3(n9081), .S3(n9484), .Z(
        \u_DataPath/from_mem_data_out_i [1]) );
  HS65_LL_MX41X7 U7027 ( .D0(n8770), .S0(n9476), .D1(n8623), .S1(n9490), .D2(
        n9497), .S2(n8767), .D3(n9081), .S3(n9483), .Z(
        \u_DataPath/from_mem_data_out_i [0]) );
  HS65_LL_MX41X4 U7049 ( .D0(n8770), .S0(n9480), .D1(n8623), .S1(n9494), .D2(
        n9501), .S2(n8767), .D3(n9081), .S3(n9487), .Z(
        \u_DataPath/from_mem_data_out_i [4]) );
  HS65_LH_MX41X7 U7051 ( .D0(n8770), .S0(n9481), .D1(n8623), .S1(n9495), .D2(
        n9502), .S2(n8767), .D3(n9081), .S3(n9488), .Z(
        \u_DataPath/from_mem_data_out_i [5]) );
  HS65_LL_MX41X4 U7059 ( .D0(n8770), .S0(n9479), .D1(n8623), .S1(n9493), .D2(
        n9500), .S2(n8767), .D3(n9081), .S3(n9486), .Z(
        \u_DataPath/from_mem_data_out_i [3]) );
  HS65_LL_NAND2X4 U7076 ( .A(n5497), .B(n9538), .Z(n3784) );
  HS65_LL_NOR2X2 U7080 ( .A(\u_DataPath/dataOut_exe_i [1]), .B(n2782), .Z(
        n8373) );
  HS65_LL_NAND2X2 U7089 ( .A(n2830), .B(n4750), .Z(n3590) );
  HS65_LL_NAND2X4 U7095 ( .A(\u_DataPath/cw_to_ex_i [0]), .B(n3587), .Z(n4653)
         );
  HS65_LL_NAND3X2 U7104 ( .A(n3300), .B(n3299), .C(n3298), .Z(n3304) );
  HS65_LL_AOI22X1 U7119 ( .A(n4610), .B(n4571), .C(n4830), .D(n4570), .Z(n4576) );
  HS65_LL_AOI22X1 U7128 ( .A(n4830), .B(n3836), .C(n4743), .D(n4571), .Z(n3655) );
  HS65_LL_NAND2X2 U7154 ( .A(n4830), .B(n4512), .Z(n4513) );
  HS65_LL_OAI12X2 U7157 ( .A(n2784), .B(n3927), .C(n4830), .Z(n3928) );
  HS65_LL_AOI22X1 U7179 ( .A(n5510), .B(n4616), .C(n4830), .D(n4615), .Z(n4628) );
  HS65_LL_AOI22X1 U7180 ( .A(n4830), .B(n4382), .C(n5510), .D(n4617), .Z(n4389) );
  HS65_LL_NAND2X2 U7182 ( .A(n4830), .B(n4616), .Z(n3299) );
  HS65_LL_AOI22X1 U7186 ( .A(n5517), .B(n4952), .C(n4830), .D(n4480), .Z(n4481) );
  HS65_LL_IVX4 U7189 ( .A(n4830), .Z(n4747) );
  HS65_LL_NAND2X4 U7223 ( .A(n3834), .B(n5208), .Z(n4674) );
  HS65_LH_NAND2X2 U7235 ( .A(n4743), .B(n4479), .Z(n3412) );
  HS65_LL_AOI22X1 U7264 ( .A(n4740), .B(n3390), .C(n4667), .D(n4479), .Z(n4482) );
  HS65_LL_AO12X4 U7266 ( .A(n4733), .B(n4732), .C(n4731), .Z(n4734) );
  HS65_LLS_XNOR2X3 U7286 ( .A(n2968), .B(n4871), .Z(n4942) );
  HS65_LL_NAND3X2 U7298 ( .A(n5347), .B(n5412), .C(n5346), .Z(n5352) );
  HS65_LL_MUXI21X2 U7308 ( .D0(n9457), .D1(n2970), .S0(n9415), .Z(n8159) );
  HS65_LH_IVX9 U7336 ( .A(\u_DataPath/from_mem_data_out_i [2]), .Z(n2970) );
  HS65_LL_NAND2X2 U7414 ( .A(n4245), .B(n4244), .Z(n4250) );
  HS65_LL_NAND3AX6 U7427 ( .A(n3387), .B(n3386), .C(n3736), .Z(n4466) );
  HS65_LL_OAI12X3 U7448 ( .A(n5490), .B(n3782), .C(n3784), .Z(n4216) );
  HS65_LL_NOR2X2 U7531 ( .A(n5497), .B(n9538), .Z(n3782) );
  HS65_LH_OAI21X2 U7537 ( .A(n3227), .B(n3226), .C(n4673), .Z(n3233) );
  HS65_LL_IVX7 U7570 ( .A(n2830), .Z(n3826) );
  HS65_LL_OAI12X3 U7594 ( .A(n9044), .B(n8744), .C(n8597), .Z(
        \u_DataPath/dataOut_exe_i [23]) );
  HS65_LL_OAI12X3 U7711 ( .A(n9044), .B(n8754), .C(n8620), .Z(
        \u_DataPath/dataOut_exe_i [30]) );
  HS65_LL_NAND2X4 U8112 ( .A(n4620), .B(n4619), .Z(n4748) );
  HS65_LH_IVX9 U8154 ( .A(n4284), .Z(n4619) );
  HS65_LL_NAND3X3 U8191 ( .A(n5177), .B(n8325), .C(n8324), .Z(n5181) );
  HS65_LL_NAND2X2 U8256 ( .A(n4788), .B(n4787), .Z(n4811) );
  HS65_LL_OAI12X3 U8273 ( .A(n7983), .B(n8585), .C(n8816), .Z(n7984) );
  HS65_LH_BFX18 U8288 ( .A(n2802), .Z(n5507) );
  HS65_LL_AO22X4 U8295 ( .A(n4671), .B(n4392), .C(n4433), .D(n4391), .Z(n4393)
         );
  HS65_LL_NAND4ABX6 U8305 ( .A(n8731), .B(n8585), .C(n7972), .D(n7971), .Z(
        \u_DataPath/cw_to_ex_i [1]) );
  HS65_LL_NAND3X2 U8311 ( .A(n3469), .B(n3468), .C(n4471), .Z(n3470) );
  HS65_LH_BFX4 U8312 ( .A(n7677), .Z(n9557) );
  HS65_LH_BFX4 U8313 ( .A(n9556), .Z(n9548) );
  HS65_LLS_XOR2X3 U8314 ( .A(n4556), .B(n4555), .Z(n9539) );
  HS65_LL_AO22X4 U8315 ( .A(n9072), .B(n9252), .C(n9278), .D(n8735), .Z(n9541)
         );
  HS65_LH_BFX4 U8357 ( .A(n9556), .Z(n9555) );
  HS65_LH_BFX4 U8368 ( .A(n9555), .Z(n9554) );
  HS65_LH_BFX4 U8369 ( .A(n9557), .Z(n9553) );
  HS65_LH_BFX4 U8503 ( .A(n9554), .Z(n9550) );
  HS65_LH_BFX4 U8564 ( .A(n9546), .Z(n9551) );
  HS65_LH_BFX4 U8568 ( .A(n9556), .Z(n9549) );
  HS65_LH_BFX4 U8602 ( .A(n9546), .Z(n9547) );
  HS65_LH_BFX4 U8603 ( .A(n9548), .Z(n9546) );
  HS65_LH_BFX4 U8604 ( .A(n9547), .Z(n9545) );
  HS65_LH_BFX4 U8606 ( .A(n9557), .Z(n9556) );
  HS65_LH_NOR2X2 U8622 ( .A(n9351), .B(n9455), .Z(n7677) );
  HS65_LL_CNHLSX7 \clk_gate_u_DataPath/u_fetch/pc1/to_iram_block_reg/latch  ( 
        .CP(clk), .E(\u_DataPath/u_fetch/pc1/N3 ), .TE(1'b0), .Q(net3007) );
  HS65_LH_DFPRQX4 clk_r_REG859_S4 ( .D(n6727), .CP(net3007), .RN(n2814), .Q(
        n9473) );
  HS65_LH_DFPQX4 clk_r_REG948_S6 ( .D(n9431), .CP(clk), .Q(n9430) );
  HS65_LL_DFPRQNX4 clk_r_REG618_S4 ( .D(n7993), .CP(net3007), .RN(n7677), .QN(
        n9565) );
  HS65_LL_DFPRQNX9 clk_r_REG598_S4 ( .D(n8022), .CP(net3007), .RN(n7677), .QN(
        n9564) );
  HS65_LL_DFPQX35 clk_r_REG198_S4 ( .D(\u_DataPath/pc_4_i [30]), .CP(net3007), 
        .Q(n8968) );
  HS65_LL_DFPQX9 clk_r_REG8_S3 ( .D(n6749), .CP(clk), .Q(n9455) );
  HS65_LL_DFPQX9 clk_r_REG626_S6 ( .D(\u_DataPath/jump_i ), .CP(clk), .Q(n9351) );
  HS65_LL_DFPRQX9 clk_r_REG619_S4 ( .D(n7970), .CP(net3007), .RN(n7677), .Q(
        n8601) );
  HS65_LH_DFPQX9 clk_r_REG706_S1 ( .D(n7013), .CP(clk), .Q(n9334) );
  HS65_LH_DFPQX4 clk_r_REG625_S5 ( .D(\u_DataPath/cw_to_ex_i [20]), .CP(clk), 
        .Q(n9446) );
  HS65_LH_DFPQX4 clk_r_REG798_S1 ( .D(n7204), .CP(clk), .Q(n9410) );
  HS65_LH_DFPQX4 clk_r_REG350_S2 ( .D(n5676), .CP(clk), .Q(n9390) );
  HS65_LH_DFPQX4 clk_r_REG41_S3 ( .D(\u_DataPath/jump_address_i [15]), .CP(clk), .Q(n9326) );
  HS65_LH_DFPQX4 clk_r_REG464_S2 ( .D(n5703), .CP(clk), .Q(n9302) );
  HS65_LH_DFPQX4 clk_r_REG612_S2 ( .D(n2930), .CP(clk), .Q(n9282) );
  HS65_LH_DFPQX4 clk_r_REG378_S2 ( .D(n5803), .CP(clk), .Q(n9237) );
  HS65_LH_DFPQX4 clk_r_REG19_S2 ( .D(n7304), .CP(clk), .Q(n9215) );
  HS65_LH_DFPQX4 clk_r_REG529_S2 ( .D(n5638), .CP(clk), .Q(n9126) );
  HS65_LH_DFPQX4 clk_r_REG272_S2 ( .D(n5881), .CP(clk), .Q(n9093) );
  HS65_LH_DFPQX4 clk_r_REG638_S6 ( .D(n8047), .CP(clk), .Q(n9071) );
  HS65_LH_DFPQX4 clk_r_REG528_S2 ( .D(n5922), .CP(clk), .Q(n9036) );
  HS65_LH_DFPQX4 clk_r_REG184_S4 ( .D(\u_DataPath/pc_4_i [28]), .CP(net3007), 
        .Q(n9020) );
  HS65_LH_DFPQX4 clk_r_REG530_S2 ( .D(n5885), .CP(clk), .Q(n9000) );
  HS65_LH_DFPQX4 clk_r_REG270_S2 ( .D(n5629), .CP(clk), .Q(n8980) );
  HS65_LH_DFPQX4 clk_r_REG154_S2 ( .D(\u_DataPath/pc_4_i [20]), .CP(net3007), 
        .Q(n8962) );
  HS65_LH_DFPQX4 clk_r_REG338_S2 ( .D(n5546), .CP(clk), .Q(n8934) );
  HS65_LH_DFPQX4 clk_r_REG486_S2 ( .D(n5659), .CP(clk), .Q(n8917) );
  HS65_LH_DFPQX4 clk_r_REG242_S2 ( .D(n5726), .CP(clk), .Q(n8897) );
  HS65_LH_DFPQX4 clk_r_REG176_S1 ( .D(\u_DataPath/branch_target_i [26]), .CP(
        clk), .Q(n8876) );
  HS65_LH_DFPQX4 clk_r_REG158_S1 ( .D(\u_DataPath/branch_target_i [20]), .CP(
        clk), .Q(n8836) );
  HS65_LH_DFPQX4 clk_r_REG434_S2 ( .D(n5537), .CP(clk), .Q(n8775) );
  HS65_LH_DFPQX4 clk_r_REG63_S3 ( .D(n8354), .CP(clk), .Q(n8756) );
  HS65_LH_DFPQX4 clk_r_REG372_S2 ( .D(n5539), .CP(clk), .Q(n8738) );
  HS65_LH_DFPQX4 clk_r_REG103_S1 ( .D(n8145), .CP(clk), .Q(n8718) );
  HS65_LH_DFPQX4 clk_r_REG67_S1 ( .D(n8237), .CP(clk), .Q(n8699) );
  HS65_LH_DFPQX4 clk_r_REG509_S3 ( .D(\u_DataPath/data_read_ex_2_i [14]), .CP(
        clk), .Q(n8683) );
  HS65_LH_DFPQX4 clk_r_REG501_S3 ( .D(\u_DataPath/data_read_ex_1_i [23]), .CP(
        clk), .Q(n8667) );
  HS65_LH_DFPQX4 clk_r_REG25_S2 ( .D(\u_DataPath/data_read_ex_2_i [28]), .CP(
        clk), .Q(n8651) );
  HS65_LH_DFPQX4 clk_r_REG544_S2 ( .D(\u_DataPath/data_read_ex_1_i [5]), .CP(
        clk), .Q(n8634) );
  HS65_LH_DFPQX4 clk_r_REG219_S3 ( .D(\u_DataPath/jump_address_i [28]), .CP(
        clk), .Q(n8618) );
  HS65_LH_DFPQX4 clk_r_REG230_S3 ( .D(n8206), .CP(clk), .Q(n8599) );
  HS65_LH_DFPQX4 clk_r_REG418_S3 ( .D(\u_DataPath/mem_writedata_out_i [18]), 
        .CP(clk), .Q(n8582) );
  HS65_LH_DFPQX4 clk_r_REG9_S4 ( .D(addr_to_iram_11), .CP(net3007), .Q(n8532)
         );
  HS65_LH_DFPQX4 clk_r_REG26_S3 ( .D(n8333), .CP(clk), .Q(n8757) );
  HS65_LH_DFPSQX18 clk_r_REG729_S4 ( .D(opcode_i[0]), .CP(net3007), .SN(n9553), 
        .Q(n8882) );
  HS65_LH_IVX4 U4667 ( .A(Data_out_fromRAM[29]), .Z(n8318) );
  HS65_LH_IVX4 U4004 ( .A(Data_out_fromRAM[26]), .Z(n8250) );
  HS65_LH_IVX4 U4666 ( .A(Data_out_fromRAM[30]), .Z(n8288) );
  HS65_LH_CNIVX3 U5154 ( .A(n8748), .Z(n3017) );
  HS65_LH_IVX9 U3933 ( .A(n8663), .Z(\u_DataPath/dataOut_exe_i [14]) );
  HS65_LH_IVX9 U3940 ( .A(n8679), .Z(\u_DataPath/dataOut_exe_i [13]) );
  HS65_LL_AOI211X1 U6596 ( .A(n9174), .B(n8600), .C(n8622), .D(n8569), .Z(
        n7972) );
  HS65_LL_NAND2X2 U6642 ( .A(n9314), .B(n9252), .Z(n8279) );
  HS65_LH_AOI21X2 U3536 ( .A(n8714), .B(n9038), .C(n8738), .Z(n5573) );
  HS65_LH_IVX7 U4072 ( .A(n8665), .Z(\u_DataPath/jump_address_i [17]) );
  HS65_LH_OR2X9 U8590 ( .A(n8553), .B(n9012), .Z(n3135) );
  HS65_LH_IVX4 U4608 ( .A(n8713), .Z(n5914) );
  HS65_LH_IVX2 U8380 ( .A(n8697), .Z(n3100) );
  HS65_LL_AOI12X4 U5026 ( .A(n9174), .B(n8706), .C(n8732), .Z(n8362) );
  HS65_LL_IVX9 U4162 ( .A(n2782), .Z(n2800) );
  HS65_LH_IVX4 U3697 ( .A(n5847), .Z(n5908) );
  HS65_LL_NAND2X5 U4979 ( .A(n8279), .B(n8768), .Z(
        \u_DataPath/dataOut_exe_i [0]) );
  HS65_LH_NOR2X3 U4149 ( .A(\u_DataPath/dataOut_exe_i [14]), .B(n9012), .Z(
        n3047) );
  HS65_LH_NOR2X5 U5835 ( .A(n9333), .B(n7629), .Z(n7433) );
  HS65_LH_IVX4 U3668 ( .A(\u_DataPath/dataOut_exe_i [29]), .Z(n3124) );
  HS65_LH_OR2X9 U3423 ( .A(\u_DataPath/dataOut_exe_i [31]), .B(n9012), .Z(
        n3238) );
  HS65_LL_IVX9 U3565 ( .A(n3236), .Z(n2710) );
  HS65_LH_IVX7 U5891 ( .A(n5775), .Z(n5894) );
  HS65_LH_AOI12X2 U4148 ( .A(n9139), .B(n5775), .C(n5746), .Z(n5793) );
  HS65_LH_CNIVX3 U5148 ( .A(\u_DataPath/cw_to_ex_i [1]), .Z(n5015) );
  HS65_LL_IVX9 U4121 ( .A(n3018), .Z(n2798) );
  HS65_LL_IVX13 U3435 ( .A(n3090), .Z(n3184) );
  HS65_LH_NAND2X5 U4906 ( .A(n8769), .B(n2712), .Z(n3013) );
  HS65_LL_OAI21X3 U5609 ( .A(n9425), .B(n8796), .C(n2982), .Z(n7674) );
  HS65_LH_NAND2X4 U4130 ( .A(n8376), .B(n2712), .Z(n2972) );
  HS65_LL_NAND2X2 U5949 ( .A(n3184), .B(n8818), .Z(n2950) );
  HS65_LL_NAND2X4 U4604 ( .A(n3174), .B(n9054), .Z(n2976) );
  HS65_LH_NAND2X5 U5012 ( .A(n9402), .B(n2798), .Z(n8392) );
  HS65_LH_NAND2X4 U7300 ( .A(n7674), .B(n2712), .Z(n2983) );
  HS65_LH_NAND2X4 U5017 ( .A(n8719), .B(n2798), .Z(n8440) );
  HS65_LH_NAND2X4 U5021 ( .A(n8718), .B(n2798), .Z(n8428) );
  HS65_LH_AOI12X3 U4541 ( .A(n7654), .B(n2798), .C(n2919), .Z(n2920) );
  HS65_LL_NAND2AX4 U6612 ( .A(n3123), .B(n3122), .Z(n4533) );
  HS65_LH_AOI22X3 U6721 ( .A(n3124), .B(n2800), .C(n8695), .D(n2798), .Z(n3125) );
  HS65_LL_OAI12X2 U8382 ( .A(\u_DataPath/dataOut_exe_i [25]), .B(n3178), .C(
        n3086), .Z(n3087) );
  HS65_LH_NOR2X3 U5048 ( .A(n3174), .B(n8417), .Z(n3042) );
  HS65_LH_NAND2X4 U4647 ( .A(\u_DataPath/cw_to_ex_i [1]), .B(n5062), .Z(n5365)
         );
  HS65_LL_OAI21X2 U3831 ( .A(n8674), .B(n3181), .C(n2972), .Z(n2973) );
  HS65_LH_OAI21X3 U6703 ( .A(\u_DataPath/dataOut_exe_i [3]), .B(n3178), .C(
        n2983), .Z(n2984) );
  HS65_LL_IVX4 U6594 ( .A(\u_DataPath/u_execute/A_inALU_i[26] ), .Z(n3975) );
  HS65_LL_IVX7 U3551 ( .A(n4918), .Z(\sub_x_51/A[21] ) );
  HS65_LH_NAND2X7 U4492 ( .A(n9354), .B(n7303), .Z(n7633) );
  HS65_LH_NAND2X5 U7152 ( .A(n4032), .B(n5079), .Z(n5356) );
  HS65_LL_NOR2X6 U3818 ( .A(n2974), .B(n2973), .Z(\lte_x_57/B[2] ) );
  HS65_LL_NOR2X2 U8573 ( .A(n2975), .B(n8159), .Z(n2980) );
  HS65_LH_NOR2X5 U4081 ( .A(n2925), .B(n8387), .Z(n4880) );
  HS65_LH_NAND2X5 U8122 ( .A(n3039), .B(n3073), .Z(n5108) );
  HS65_LH_AOI22X1 U4957 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][9] ), .B(n9242), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][9] ), .D(n8861), .Z(n7068) );
  HS65_LH_AOI22X1 U4931 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][26] ), .B(n9242), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][26] ), .D(
        n8861), .Z(n6793) );
  HS65_LH_IVX2 U9374 ( .A(n8219), .Z(n8221) );
  HS65_LL_IVX7 U3377 ( .A(n4794), .Z(n2802) );
  HS65_LH_IVX9 U3783 ( .A(\lte_x_57/B[4] ), .Z(n3948) );
  HS65_LL_NAND2X4 U3414 ( .A(n4533), .B(n5196), .Z(n5445) );
  HS65_LL_IVX4 U5599 ( .A(n4870), .Z(n3222) );
  HS65_LHS_XOR2X3 U8285 ( .A(n4533), .B(n5196), .Z(n4963) );
  HS65_LH_NAND2X5 U5471 ( .A(n5529), .B(n5067), .Z(n5303) );
  HS65_LH_NOR2X5 U5538 ( .A(\lte_x_57/B[15] ), .B(n5084), .Z(n3896) );
  HS65_LH_NAND2X5 U5548 ( .A(\u_DataPath/u_execute/A_inALU_i[26] ), .B(n5190), 
        .Z(n4602) );
  HS65_LH_NAND2X5 U3621 ( .A(\sub_x_51/A[27] ), .B(n3106), .Z(n3355) );
  HS65_LH_NAND2X5 U5555 ( .A(\lte_x_57/B[28] ), .B(n4902), .Z(n4522) );
  HS65_LH_AOI22X1 U6630 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][22] ), .B(n9242), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][22] ), .D(
        n9166), .Z(n7188) );
  HS65_LH_NOR2X5 U3619 ( .A(\sub_x_51/A[8] ), .B(n5201), .Z(n4275) );
  HS65_LH_NOR2X5 U5424 ( .A(n5192), .B(n5067), .Z(n3419) );
  HS65_LL_NOR2X2 U5556 ( .A(\lte_x_57/B[29] ), .B(n5196), .Z(n4519) );
  HS65_LH_NAND2X7 U4171 ( .A(\u_DataPath/cw_to_ex_i [2]), .B(n3292), .Z(n7315)
         );
  HS65_LH_AOI22X1 U5696 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][12] ), .B(n9242), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][12] ), .D(
        n8861), .Z(n7148) );
  HS65_LL_OAI12X5 U3815 ( .A(n2993), .B(n2844), .C(n2992), .Z(n3251) );
  HS65_LH_AOI22X1 U3771 ( .A(n9243), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][0] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][0] ), .D(n9197), 
        .Z(n7287) );
  HS65_LH_AOI22X1 U4968 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][5] ), .B(n9242), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][5] ), .D(n8861), .Z(n7088) );
  HS65_LH_AOI22X1 U5618 ( .A(n9207), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][0] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][0] ), .D(n9095), 
        .Z(n7288) );
  HS65_LH_AOI22X1 U6699 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][4] ), .B(n9242), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][4] ), .D(n8861), .Z(n6032) );
  HS65_LH_AOI22X1 U6698 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][2] ), .B(n9242), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][2] ), .D(n9166), .Z(n6154) );
  HS65_LL_AOI12X6 U5562 ( .A(n2798), .B(n2980), .C(n2979), .Z(n5092) );
  HS65_LL_IVX7 U4443 ( .A(n3241), .Z(n5208) );
  HS65_LL_IVX7 U3386 ( .A(n5508), .Z(n5487) );
  HS65_LH_NOR2X5 U8236 ( .A(n5192), .B(n3200), .Z(n5193) );
  HS65_LH_IVX4 U4036 ( .A(n4718), .Z(n4719) );
  HS65_LH_NOR2X5 U5578 ( .A(n5385), .B(n3338), .Z(n4316) );
  HS65_LH_IVX7 U4027 ( .A(n5304), .Z(n4997) );
  HS65_LL_IVX7 U4893 ( .A(n3247), .Z(n5072) );
  HS65_LH_NAND2X4 U4022 ( .A(n4684), .B(n4687), .Z(n3281) );
  HS65_LH_NAND2X5 U4808 ( .A(n5455), .B(n5450), .Z(n4003) );
  HS65_LH_CNIVX3 U4802 ( .A(n3353), .Z(n3354) );
  HS65_LH_CNIVX3 U4447 ( .A(n4602), .Z(n3359) );
  HS65_LH_CNIVX3 U8265 ( .A(n4258), .Z(n3677) );
  HS65_LH_CNIVX3 U3609 ( .A(n5516), .Z(n4944) );
  HS65_LH_NAND2X5 U8120 ( .A(\lte_x_57/B[11] ), .B(n3075), .Z(n5111) );
  HS65_LH_IVX9 U7131 ( .A(n5187), .Z(n3187) );
  HS65_LHS_XNOR2X3 U8720 ( .A(\lte_x_57/B[2] ), .B(n5092), .Z(n4948) );
  HS65_LH_IVX4 U3601 ( .A(n4681), .Z(n3275) );
  HS65_LH_IVX4 U4464 ( .A(n3861), .Z(n3862) );
  HS65_LL_IVX9 U4685 ( .A(n2995), .Z(n5211) );
  HS65_LH_NAND2X7 U4014 ( .A(n4338), .B(n4337), .Z(n4344) );
  HS65_LH_NOR2X3 U4466 ( .A(n2825), .B(n2829), .Z(n3715) );
  HS65_LHS_XOR2X3 U7699 ( .A(\lte_x_57/B[4] ), .B(n5208), .Z(n4987) );
  HS65_LH_NAND2X5 U4423 ( .A(n5145), .B(n4641), .Z(n3212) );
  HS65_LH_IVX2 U7696 ( .A(n4884), .Z(n4885) );
  HS65_LH_NOR2X2 U4418 ( .A(n5146), .B(n5070), .Z(n5071) );
  HS65_LH_NAND2X5 U3711 ( .A(\lte_x_57/B[4] ), .B(n2792), .Z(n3807) );
  HS65_LL_CNIVX3 U6460 ( .A(n3539), .Z(n3248) );
  HS65_LH_NOR2X2 U4816 ( .A(n4533), .B(n3225), .Z(n3327) );
  HS65_LH_NOR2X5 U4001 ( .A(n5311), .B(n4738), .Z(n3242) );
  HS65_LH_NAND2X4 U3708 ( .A(\sub_x_51/A[27] ), .B(n3826), .Z(n3328) );
  HS65_LH_NOR2X3 U7134 ( .A(n5311), .B(n2829), .Z(n4658) );
  HS65_LH_NOR2X2 U8287 ( .A(n4846), .B(n3204), .Z(n4504) );
  HS65_LH_NAND2X5 U5452 ( .A(n5517), .B(n4985), .Z(n4033) );
  HS65_LL_IVX7 U4468 ( .A(n2829), .Z(n5498) );
  HS65_LH_NAND2X4 U5341 ( .A(n3355), .B(n3354), .Z(n3364) );
  HS65_LH_NAND2X5 U3996 ( .A(n4522), .B(n4412), .Z(n4418) );
  HS65_LH_NOR2X2 U5525 ( .A(n2825), .B(n3225), .Z(n3490) );
  HS65_LL_AOI12X2 U4420 ( .A(n5312), .B(n5311), .C(n5014), .Z(n4011) );
  HS65_LH_NOR2X3 U5508 ( .A(n4630), .B(n4964), .Z(n3303) );
  HS65_LH_IVX7 U4469 ( .A(n3848), .Z(n3849) );
  HS65_LH_NAND2X7 U5512 ( .A(\lte_x_57/B[29] ), .B(n3742), .Z(n3484) );
  HS65_LH_IVX4 U4381 ( .A(n3664), .Z(n3665) );
  HS65_LH_CNIVX3 U8183 ( .A(n5006), .Z(n5000) );
  HS65_LH_IVX2 U7026 ( .A(n4596), .Z(n3311) );
  HS65_LH_CNIVX3 U3655 ( .A(n4431), .Z(n3285) );
  HS65_LL_CNBFX14 U4030 ( .A(n2796), .Z(n5496) );
  HS65_LH_CNIVX3 U8328 ( .A(n3715), .Z(n3346) );
  HS65_LH_OAI21X2 U4408 ( .A(n5286), .B(n5004), .C(n5298), .Z(n5001) );
  HS65_LH_MUX21I1X6 U6415 ( .D0(n3242), .D1(n4431), .S0(n2830), .Z(n3243) );
  HS65_LL_AOI12X2 U8159 ( .A(n5349), .B(n5341), .C(n5334), .Z(n3953) );
  HS65_LH_NAND2X5 U5322 ( .A(n5262), .B(n5194), .Z(n5198) );
  HS65_LH_CNIVX3 U8304 ( .A(n3825), .Z(n3830) );
  HS65_LH_IVX2 U8215 ( .A(n4212), .Z(n4213) );
  HS65_LH_IVX2 U7694 ( .A(n5341), .Z(n4883) );
  HS65_LH_NAND3X3 U4383 ( .A(n4884), .B(n5028), .C(n5024), .Z(n4897) );
  HS65_LH_NAND2X4 U3692 ( .A(n5024), .B(n5023), .Z(n5387) );
  HS65_LH_IVX4 U4409 ( .A(n4216), .Z(n4803) );
  HS65_LH_IVX2 U7039 ( .A(n5373), .Z(n5374) );
  HS65_LH_NAND2X4 U4806 ( .A(n5452), .B(n5303), .Z(n3976) );
  HS65_LH_IVX4 U8661 ( .A(n3536), .Z(n3537) );
  HS65_LL_AOI12X2 U3957 ( .A(n3267), .B(n4376), .C(n3266), .Z(n3455) );
  HS65_LL_NAND3X2 U3822 ( .A(n3864), .B(n3863), .C(n3862), .Z(n5483) );
  HS65_LH_AOI12X6 U3507 ( .A(\sub_x_51/A[13] ), .B(n5496), .C(n3342), .Z(n3916) );
  HS65_LL_OAI12X2 U4511 ( .A(n4367), .B(n3636), .C(n5127), .Z(n3190) );
  HS65_LH_IVX4 U3623 ( .A(n3569), .Z(n3570) );
  HS65_LL_IVX2 U6377 ( .A(n3267), .Z(n3249) );
  HS65_LH_NAND2X4 U4828 ( .A(n3584), .B(n3583), .Z(n3585) );
  HS65_LH_CNIVX3 U4406 ( .A(n4770), .Z(n4185) );
  HS65_LH_NAND2X4 U4829 ( .A(n3582), .B(n3581), .Z(n3586) );
  HS65_LH_CNIVX3 U6376 ( .A(n4458), .Z(n4459) );
  HS65_LH_NAND2X5 U4364 ( .A(n4767), .B(n4766), .Z(n4772) );
  HS65_LH_CNIVX3 U8696 ( .A(n4850), .Z(n3718) );
  HS65_LH_OAI21X3 U6484 ( .A(n3379), .B(n4192), .C(n4191), .Z(n4193) );
  HS65_LH_NOR2X5 U5272 ( .A(n4644), .B(n4638), .Z(n4647) );
  HS65_LH_NAND2X4 U3631 ( .A(n3574), .B(n3572), .Z(n3296) );
  HS65_LH_NAND2X4 U4434 ( .A(\sub_x_51/A[18] ), .B(n5496), .Z(n3644) );
  HS65_LL_OAI21X2 U3823 ( .A(n3993), .B(n3338), .C(n3643), .Z(n3645) );
  HS65_LH_CNIVX3 U4386 ( .A(n4603), .Z(n3357) );
  HS65_LH_IVX4 U4753 ( .A(n4610), .Z(n4753) );
  HS65_LH_NAND3X3 U5346 ( .A(n3408), .B(n3407), .C(n3406), .Z(n4512) );
  HS65_LH_NAND2X2 U3949 ( .A(n5231), .B(n5202), .Z(n5206) );
  HS65_LL_OAI12X2 U8220 ( .A(n4426), .B(n5245), .C(n5244), .Z(n5249) );
  HS65_LH_NAND2X5 U6381 ( .A(n3538), .B(n3537), .Z(n3544) );
  HS65_LH_IVX4 U3939 ( .A(n3883), .Z(n3884) );
  HS65_LH_OAI21X3 U8322 ( .A(n3591), .B(n4738), .C(n3243), .Z(n4392) );
  HS65_LL_IVX7 U3564 ( .A(n5481), .Z(n4294) );
  HS65_LL_OAI12X2 U6254 ( .A(n4541), .B(n4643), .C(n5140), .Z(n4542) );
  HS65_LH_IVX7 U6335 ( .A(n4392), .Z(n4614) );
  HS65_LH_IVX4 U4397 ( .A(n4827), .Z(n4254) );
  HS65_LL_OAI12X2 U5309 ( .A(n3275), .B(n4689), .C(n3274), .Z(n3276) );
  HS65_LH_CNIVX3 U3938 ( .A(n3695), .Z(n3698) );
  HS65_LH_IVX7 U5284 ( .A(n4177), .Z(n4090) );
  HS65_LH_NAND2X5 U3577 ( .A(n5255), .B(n5185), .Z(n5258) );
  HS65_LH_IVX2 U7031 ( .A(n5435), .Z(n5053) );
  HS65_LH_CNIVX3 U4788 ( .A(n3692), .Z(n3693) );
  HS65_LH_OAI21X3 U6320 ( .A(n5258), .B(n5257), .C(n5256), .Z(n5274) );
  HS65_LH_NOR2X3 U3928 ( .A(n4014), .B(n3990), .Z(n4017) );
  HS65_LH_NOR2X5 U3597 ( .A(n5429), .B(n5428), .Z(n5430) );
  HS65_LL_OAI12X5 U3887 ( .A(n2823), .B(n2828), .C(n2860), .Z(n4732) );
  HS65_LH_NOR2X5 U7019 ( .A(n4321), .B(n4614), .Z(n3244) );
  HS65_LH_NOR2X2 U5303 ( .A(n4292), .B(n4068), .Z(n3802) );
  HS65_LH_OAI21X3 U5327 ( .A(n4514), .B(n5499), .C(n4513), .Z(n4515) );
  HS65_LL_NOR2X5 U3630 ( .A(n3454), .B(n3271), .Z(n4683) );
  HS65_LH_IVX7 U4384 ( .A(n4111), .Z(n4615) );
  HS65_LL_AOI12X2 U7714 ( .A(n5465), .B(n5464), .C(n5463), .Z(n5467) );
  HS65_LH_NOR2X5 U5294 ( .A(n4709), .B(n4705), .Z(n4712) );
  HS65_LH_IVX2 U3547 ( .A(n5461), .Z(n5468) );
  HS65_LH_NAND2X5 U4716 ( .A(n4618), .B(n5511), .Z(n4558) );
  HS65_LH_OAI211X3 U6272 ( .A(n4653), .B(n4783), .C(n3546), .D(n3545), .Z(
        n3548) );
  HS65_LH_NOR3X1 U4738 ( .A(n4674), .B(n5211), .C(n4146), .Z(n3479) );
  HS65_LH_IVX7 U4790 ( .A(n3836), .Z(n4562) );
  HS65_LH_IVX7 U4787 ( .A(n4070), .Z(n4478) );
  HS65_LH_NAND2X5 U6221 ( .A(n5484), .B(n4066), .Z(n4030) );
  HS65_LL_OAI12X5 U3525 ( .A(n4105), .B(n3199), .C(n3198), .Z(n4646) );
  HS65_LL_AOI112X1 U6282 ( .A(n4692), .B(n3360), .C(n3359), .D(n3358), .Z(
        n3361) );
  HS65_LH_NAND2X4 U3852 ( .A(n4721), .B(n4723), .Z(n4137) );
  HS65_LH_IVX7 U4748 ( .A(n4480), .Z(n4506) );
  HS65_LH_NAND2X7 U4373 ( .A(n5505), .B(n4334), .Z(n4335) );
  HS65_LH_OAI21X3 U4715 ( .A(n3288), .B(n3287), .C(n5510), .Z(n3289) );
  HS65_LH_NAND2X4 U5251 ( .A(n4490), .B(n4723), .Z(n4492) );
  HS65_LH_NAND2X2 U8272 ( .A(n4667), .B(n4615), .Z(n3298) );
  HS65_LH_NAND2AX4 U4705 ( .A(n4154), .B(n4153), .Z(n4155) );
  HS65_LL_NOR2X5 U3850 ( .A(n4104), .B(n3199), .Z(n4639) );
  HS65_LL_AOI12X2 U6994 ( .A(n3277), .B(n4692), .C(n3276), .Z(n3278) );
  HS65_LH_IVX2 U4362 ( .A(n4039), .Z(n3803) );
  HS65_LH_NAND2X5 U3501 ( .A(n7325), .B(n4051), .Z(n4052) );
  HS65_LL_OAI12X2 U3671 ( .A(n3542), .B(n4695), .C(n3541), .Z(n3543) );
  HS65_LL_NAND2X4 U3418 ( .A(n3649), .B(n3648), .Z(n5485) );
  HS65_LL_AOI12X2 U6991 ( .A(n4551), .B(n4646), .C(n3374), .Z(n3375) );
  HS65_LH_OAI21X3 U3803 ( .A(n4281), .B(n5481), .C(n4160), .Z(n4161) );
  HS65_LL_OAI12X2 U4317 ( .A(n4511), .B(n4744), .C(n4510), .Z(n4516) );
  HS65_LL_AOI12X2 U4348 ( .A(n4596), .B(n4646), .C(n4595), .Z(n4597) );
  HS65_LL_AOI12X2 U3888 ( .A(n5443), .B(n5442), .C(n5441), .Z(n5474) );
  HS65_LL_OAI12X2 U3419 ( .A(n4137), .B(n4695), .C(n4136), .Z(n4138) );
  HS65_LH_OAI22X3 U6247 ( .A(n4659), .B(n4506), .C(n4441), .D(n4665), .Z(n4442) );
  HS65_LL_IVX2 U4315 ( .A(n3600), .Z(n3601) );
  HS65_LL_AOI12X2 U6958 ( .A(n4676), .B(n4675), .C(n4674), .Z(n4677) );
  HS65_LH_NAND2X5 U6150 ( .A(n7325), .B(n3661), .Z(n3662) );
  HS65_LL_OAI112X1 U6178 ( .A(n3320), .B(n3334), .C(n3333), .D(n3332), .Z(
        n3368) );
  HS65_LL_OAI12X3 U3382 ( .A(n3892), .B(n4273), .C(n3891), .Z(n3893) );
  HS65_LH_NOR2X3 U3890 ( .A(n4738), .B(n3868), .Z(n3497) );
  HS65_LL_NAND3X2 U3410 ( .A(n3291), .B(n3290), .C(n3289), .Z(n3305) );
  HS65_LL_OAI12X2 U3388 ( .A(n4107), .B(n4714), .C(n4106), .Z(n4108) );
  HS65_LLS_XOR2X3 U3387 ( .A(n3651), .B(n4714), .Z(n3652) );
  HS65_LL_OAI12X2 U4146 ( .A(n4554), .B(n4714), .C(n4553), .Z(n4555) );
  HS65_LL_OAI12X3 U3391 ( .A(n3376), .B(n4714), .C(n3375), .Z(n3377) );
  HS65_LL_OAI12X2 U4697 ( .A(n4714), .B(n3210), .C(n3209), .Z(n3211) );
  HS65_LL_OAI12X3 U3389 ( .A(n4104), .B(n4714), .C(n4105), .Z(n3499) );
  HS65_LH_NAND2X4 U3643 ( .A(n5492), .B(n4583), .Z(n4584) );
  HS65_LL_IVX2 U3489 ( .A(n4758), .Z(n4759) );
  HS65_LL_OAI12X3 U3390 ( .A(n4402), .B(n4714), .C(n4401), .Z(n4403) );
  HS65_LL_NAND2X2 U3870 ( .A(n5492), .B(n4419), .Z(n4420) );
  HS65_LL_NAND3X2 U4105 ( .A(n4054), .B(n4053), .C(n4052), .Z(n4055) );
  HS65_LL_CNIVX3 U8725 ( .A(n8344), .Z(n4360) );
  HS65_LL_NOR3X1 U4688 ( .A(n4302), .B(n4301), .C(n4300), .Z(n4303) );
  HS65_LL_NAND3X2 U4305 ( .A(n4143), .B(n4142), .C(n4141), .Z(n4144) );
  HS65_LL_NAND3X2 U4680 ( .A(n4586), .B(n4585), .C(n4584), .Z(n4587) );
  HS65_LH_IVX9 U3874 ( .A(n3705), .Z(n3706) );
  HS65_LL_NAND2X2 U3459 ( .A(n7327), .B(n3501), .Z(n3502) );
  HS65_LH_NAND2AX7 U4307 ( .A(n3707), .B(n3706), .Z(n3708) );
  HS65_LL_AOI21X2 U3416 ( .A(n7327), .B(n4457), .C(n4456), .Z(n8332) );
  HS65_LL_CB4I6X4 U3865 ( .A(n5528), .B(n5527), .C(n5526), .D(n5525), .Z(n8356) );
  HS65_LL_NOR3X2 U3380 ( .A(n7445), .B(n8352), .C(n8353), .Z(n4365) );
  HS65_LH_IVX2 U8409 ( .A(Data_out_fromRAM[31]), .Z(n8311) );
  HS65_LH_IVX9 U3962 ( .A(n8662), .Z(\u_DataPath/dataOut_exe_i [12]) );
  HS65_LH_NOR2X2 U4562 ( .A(n8747), .B(n9012), .Z(n2974) );
  HS65_LL_AND2ABX35 U5734 ( .A(n9351), .B(n9455), .Z(n2814) );
  HS65_LHS_XOR2X3 U8792 ( .A(n8917), .B(n9238), .Z(\u_DataPath/toPC2_i [2]) );
  HS65_LH_IVX4 U3968 ( .A(n8732), .Z(n7959) );
  HS65_LL_AOI211X2 U5006 ( .A(n9400), .B(n9211), .C(n8742), .D(n8569), .Z(
        n7977) );
  HS65_LL_OA112X4 U5637 ( .A(n9021), .B(n8723), .C(n8605), .D(n7959), .Z(n8000) );
  HS65_LH_IVX9 U3930 ( .A(\u_DataPath/dataOut_exe_i [1]), .Z(n8045) );
  HS65_LH_NOR2X5 U5882 ( .A(n8639), .B(n2800), .Z(n3215) );
  HS65_LH_NAND2X5 U3569 ( .A(n8296), .B(n2800), .Z(n8380) );
  HS65_LHS_XNOR2X3 U6720 ( .A(n9231), .B(n7429), .Z(
        \u_DataPath/u_execute/link_value_i [15]) );
  HS65_LHS_XNOR2X3 U5024 ( .A(n9380), .B(n7437), .Z(
        \u_DataPath/u_execute/link_value_i [14]) );
  HS65_LH_NOR2X5 U4139 ( .A(\u_DataPath/dataOut_exe_i [26]), .B(n3980), .Z(
        n3113) );
  HS65_LH_IVX9 U6066 ( .A(\u_DataPath/cw_to_ex_i [4]), .Z(n4018) );
  HS65_LH_NOR2X5 U8567 ( .A(n8670), .B(n3181), .Z(n2946) );
  HS65_LH_NAND2X4 U4908 ( .A(n9222), .B(n2797), .Z(n8370) );
  HS65_LH_AOI12X6 U7270 ( .A(n8771), .B(n2712), .C(n2928), .Z(n2929) );
  HS65_LH_NOR2AX13 U3425 ( .A(\u_DataPath/dataOut_exe_i [14]), .B(n3567), .Z(
        n3442) );
  HS65_LH_NOR2AX13 U6687 ( .A(\u_DataPath/dataOut_exe_i [13]), .B(n3567), .Z(
        n3533) );
  HS65_LH_NOR2AX13 U6686 ( .A(n8748), .B(n3567), .Z(n3441) );
  HS65_LH_NOR2AX13 U6684 ( .A(\u_DataPath/dataOut_exe_i [6]), .B(n3567), .Z(
        n3506) );
  HS65_LH_NOR2X5 U4876 ( .A(n8627), .B(n3181), .Z(n3088) );
  HS65_LL_NOR2AX6 U8668 ( .A(n8582), .B(n3450), .Z(n3557) );
  HS65_LL_NOR2AX6 U8657 ( .A(n8575), .B(n3450), .Z(n3525) );
  HS65_LL_NOR2AX6 U8654 ( .A(n8580), .B(n3450), .Z(n3519) );
  HS65_LL_NOR2AX6 U8655 ( .A(n8571), .B(n3450), .Z(n3521) );
  HS65_LL_NOR2AX6 U8653 ( .A(n8570), .B(n3450), .Z(n3517) );
  HS65_LL_NOR2AX6 U8648 ( .A(n8685), .B(n3450), .Z(n3507) );
  HS65_LH_IVX2 U6675 ( .A(n5183), .Z(n8372) );
  HS65_LL_NOR2AX6 U8670 ( .A(n8577), .B(n3450), .Z(n3559) );
  HS65_LL_NOR2AX6 U8667 ( .A(n8583), .B(n3450), .Z(n3555) );
  HS65_LL_NOR2AX6 U8649 ( .A(n8576), .B(n3450), .Z(n3509) );
  HS65_LL_NOR2AX6 U8650 ( .A(n8705), .B(n3450), .Z(n3511) );
  HS65_LL_NOR2AX6 U8652 ( .A(n8566), .B(n3450), .Z(n3515) );
  HS65_LL_NOR2AX6 U8651 ( .A(n8573), .B(n3450), .Z(n3513) );
  HS65_LL_NOR2AX6 U8640 ( .A(n8643), .B(n3450), .Z(n3451) );
  HS65_LHS_XNOR2X3 U6718 ( .A(n8896), .B(n5717), .Z(\u_DataPath/toPC2_i [21])
         );
  HS65_LHS_XNOR2X6 U4845 ( .A(n8918), .B(n5682), .Z(\u_DataPath/toPC2_i [16])
         );
  HS65_LH_NAND2X7 U4219 ( .A(n3174), .B(n9434), .Z(n3050) );
  HS65_LHS_XNOR2X3 U6615 ( .A(n9383), .B(n7425), .Z(
        \u_DataPath/u_execute/link_value_i [17]) );
  HS65_LH_NAND2X5 U3613 ( .A(n3184), .B(n9143), .Z(n2939) );
  HS65_LH_NAND2X4 U4214 ( .A(n3184), .B(n8730), .Z(n3164) );
  HS65_LH_NAND2X4 U4215 ( .A(n3184), .B(n8730), .Z(n3169) );
  HS65_LH_NAND2X4 U6824 ( .A(n3184), .B(n8730), .Z(n3177) );
  HS65_LH_NOR2X3 U4982 ( .A(n6760), .B(n2794), .Z(n8411) );
  HS65_LH_NAND2X5 U4992 ( .A(n3168), .B(n8440), .Z(n3170) );
  HS65_LH_NAND2X5 U5776 ( .A(n3049), .B(n8416), .Z(n3051) );
  HS65_LL_OAI12X6 U3378 ( .A(n3070), .B(n2839), .C(n3069), .Z(n5082) );
  HS65_LH_NOR2AX13 U6713 ( .A(n8762), .B(n3568), .Z(n3445) );
  HS65_LH_NOR2AX13 U6715 ( .A(n9120), .B(n3568), .Z(n3447) );
  HS65_LH_NOR2AX13 U6716 ( .A(n9121), .B(n3568), .Z(n3448) );
  HS65_LHS_XNOR2X3 U8535 ( .A(n8932), .B(n5678), .Z(\u_DataPath/toPC2_i [14])
         );
  HS65_LHS_XNOR2X3 U4981 ( .A(n8897), .B(n5725), .Z(\u_DataPath/toPC2_i [23])
         );
  HS65_LH_IVX7 U4915 ( .A(\lte_x_57/B[25] ), .Z(n5016) );
  HS65_LH_NAND2X7 U3820 ( .A(n3039), .B(n5079), .Z(n4048) );
  HS65_LH_IVX9 U4914 ( .A(\lte_x_57/B[3] ), .Z(n4189) );
  HS65_LH_IVX9 U6582 ( .A(n4902), .Z(n2791) );
  HS65_LH_NAND2X7 U6541 ( .A(\lte_x_57/B[15] ), .B(n5084), .Z(n3898) );
  HS65_LH_NAND2X7 U6486 ( .A(n5192), .B(n5067), .Z(n4578) );
  HS65_LL_IVX7 U3549 ( .A(n5063), .Z(n3188) );
  HS65_LH_NOR2X6 U3998 ( .A(\sub_x_51/A[27] ), .B(n3106), .Z(n3353) );
  HS65_LL_NAND2AX4 U3828 ( .A(n3095), .B(n3094), .Z(n3247) );
  HS65_LH_IVX7 U4010 ( .A(n4046), .Z(n4047) );
  HS65_LH_CNIVX3 U6475 ( .A(n4985), .Z(n4990) );
  HS65_LH_CNIVX3 U8151 ( .A(n4974), .Z(n4977) );
  HS65_LH_CNIVX3 U8152 ( .A(n4975), .Z(n4976) );
  HS65_LH_IVX2 U8149 ( .A(n4963), .Z(n4966) );
  HS65_LH_NOR2X3 U3617 ( .A(n5393), .B(n2830), .Z(n3580) );
  HS65_LH_NOR2X6 U8765 ( .A(\lte_x_57/B[29] ), .B(n3204), .Z(n5070) );
  HS65_LH_NOR2X3 U6565 ( .A(n4283), .B(n3338), .Z(n3335) );
  HS65_LL_IVX7 U4909 ( .A(n2830), .Z(n4796) );
  HS65_LL_NAND2X7 U3562 ( .A(n3222), .B(n9538), .Z(n3225) );
  HS65_LH_NOR2X3 U4040 ( .A(n3054), .B(n3338), .Z(n3342) );
  HS65_LH_IVX9 U5410 ( .A(n3419), .Z(n4577) );
  HS65_LH_NAND2X7 U3763 ( .A(n5284), .B(n5303), .Z(n5299) );
  HS65_LH_NOR2X6 U8134 ( .A(\lte_x_57/B[10] ), .B(n3074), .Z(n5107) );
  HS65_LH_NOR2X6 U6476 ( .A(\lte_x_57/B[4] ), .B(n5208), .Z(n3759) );
  HS65_LH_OAI22X3 U8619 ( .A(n3975), .B(n2829), .C(n2830), .D(n3103), .Z(n3347) );
  HS65_LH_IVX7 U4825 ( .A(n3842), .Z(n3768) );
  HS65_LH_NAND2X7 U8165 ( .A(\lte_x_57/B[11] ), .B(n3075), .Z(n5228) );
  HS65_LH_IVX2 U8361 ( .A(n3372), .Z(n3373) );
  HS65_LH_NOR2X3 U3978 ( .A(n4630), .B(n4970), .Z(n3369) );
  HS65_LH_NOR2X6 U4044 ( .A(n3950), .B(n2829), .Z(n3844) );
  HS65_LH_NAND2X7 U5473 ( .A(n4687), .B(n4681), .Z(n4690) );
  HS65_LH_NOR2X5 U4871 ( .A(n3065), .B(n3322), .Z(n4204) );
  HS65_LH_NOR2X5 U4682 ( .A(n4871), .B(n3322), .Z(n3475) );
  HS65_LH_IVX7 U4780 ( .A(n4552), .Z(n3374) );
  HS65_LH_OAI22X3 U8615 ( .A(n4383), .B(n2829), .C(n2830), .D(n3993), .Z(n3325) );
  HS65_LH_NAND2X7 U4387 ( .A(n4277), .B(n4276), .Z(n4278) );
  HS65_LH_NAND2X4 U3936 ( .A(n4078), .B(n3258), .Z(n4086) );
  HS65_LH_IVX4 U6459 ( .A(n4818), .Z(n4819) );
  HS65_LH_NAND2X7 U5476 ( .A(n4910), .B(n5187), .Z(n5288) );
  HS65_LH_CNIVX3 U7125 ( .A(n5495), .Z(n5501) );
  HS65_LH_NAND3X5 U5319 ( .A(n5350), .B(n5349), .C(n5348), .Z(n5351) );
  HS65_LH_IVX7 U3961 ( .A(n4765), .Z(n4766) );
  HS65_LH_NAND2X4 U6428 ( .A(n3767), .B(n3766), .Z(n3770) );
  HS65_LH_NOR2X3 U8222 ( .A(\add_x_50/A[19] ), .B(n3189), .Z(n5247) );
  HS65_LH_NAND2X7 U5505 ( .A(n3784), .B(n3783), .Z(n3785) );
  HS65_LH_IVX9 U3988 ( .A(n3759), .Z(n3874) );
  HS65_LH_CNIVX3 U8724 ( .A(n4862), .Z(n4350) );
  HS65_LH_NAND2X4 U6361 ( .A(n4237), .B(n4238), .Z(n3669) );
  HS65_LH_NAND2X4 U4596 ( .A(\add_x_50/A[19] ), .B(n3742), .Z(n3569) );
  HS65_LH_CNIVX7 U4414 ( .A(n5010), .Z(n4930) );
  HS65_LH_CNIVX3 U8176 ( .A(n5348), .Z(n5340) );
  HS65_LH_NAND2X5 U3954 ( .A(n4552), .B(n4551), .Z(n4556) );
  HS65_LH_IVX7 U5407 ( .A(n4488), .Z(n4489) );
  HS65_LH_IVX7 U3604 ( .A(n3379), .Z(n4149) );
  HS65_LH_NOR2X5 U3635 ( .A(n4775), .B(n4317), .Z(n3386) );
  HS65_LH_CNIVX3 U5388 ( .A(n4946), .Z(n4947) );
  HS65_LH_CNIVX3 U8153 ( .A(n4952), .Z(n4953) );
  HS65_LH_NAND2X4 U8716 ( .A(n4781), .B(n5251), .Z(n4129) );
  HS65_LH_NAND2X5 U3616 ( .A(\lte_x_57/B[25] ), .B(n3742), .Z(n3488) );
  HS65_LH_AOI12X2 U8331 ( .A(n4641), .B(n4640), .C(n5444), .Z(n4642) );
  HS65_LH_NAND2X4 U4797 ( .A(n5009), .B(n3310), .Z(n3318) );
  HS65_LH_IVX4 U3987 ( .A(n5292), .Z(n5282) );
  HS65_LH_NAND2X7 U4775 ( .A(n5301), .B(n5005), .Z(n5007) );
  HS65_LH_NOR2X5 U3787 ( .A(n3903), .B(n3259), .Z(n3905) );
  HS65_LH_NOR2X6 U4778 ( .A(n3976), .B(n4003), .Z(n3989) );
  HS65_LH_CNIVX3 U4818 ( .A(n3788), .Z(n3789) );
  HS65_LH_NAND2X4 U6386 ( .A(n4487), .B(n3250), .Z(n4494) );
  HS65_LH_CNIVX3 U4781 ( .A(n5245), .Z(n4425) );
  HS65_LH_NAND2X7 U3970 ( .A(n5125), .B(n5051), .Z(n5435) );
  HS65_LH_IVX4 U8277 ( .A(n4823), .Z(n4339) );
  HS65_LH_IVX2 U6384 ( .A(n4912), .Z(n4913) );
  HS65_LH_AOI12X2 U6379 ( .A(n3248), .B(n4376), .C(n3540), .Z(n3541) );
  HS65_LH_IVX9 U3615 ( .A(n3228), .Z(n4115) );
  HS65_LH_NAND2X7 U3625 ( .A(n4448), .B(n3659), .Z(n3660) );
  HS65_LH_NAND3X5 U5338 ( .A(n4991), .B(n4990), .C(n4989), .Z(n4992) );
  HS65_LL_AOI12X2 U4506 ( .A(n4724), .B(n3269), .C(n3268), .Z(n3270) );
  HS65_LH_CNIVX3 U8743 ( .A(n4724), .Z(n4726) );
  HS65_LH_NAND2X7 U3611 ( .A(\sub_x_51/A[5] ), .B(n5496), .Z(n4777) );
  HS65_LH_IVX7 U4000 ( .A(n4468), .Z(n4063) );
  HS65_LH_OA12X4 U4771 ( .A(n3966), .B(n3965), .C(n3964), .Z(n2833) );
  HS65_LH_NOR2X2 U8235 ( .A(n4458), .B(n5184), .Z(n5185) );
  HS65_LH_CNIVX3 U4378 ( .A(n4325), .Z(n4326) );
  HS65_LH_NAND2X4 U4776 ( .A(n5434), .B(n5433), .Z(n5462) );
  HS65_LH_NOR2X6 U5367 ( .A(n5283), .B(n5282), .Z(n5293) );
  HS65_LH_IVX4 U7028 ( .A(n4369), .Z(n4370) );
  HS65_LH_OAI12X3 U6344 ( .A(n5003), .B(n5290), .C(n5292), .Z(n5463) );
  HS65_LH_IVX2 U7606 ( .A(n5038), .Z(n5048) );
  HS65_LH_IVX2 U4502 ( .A(n5413), .Z(n5044) );
  HS65_LH_NOR2X6 U5295 ( .A(n3888), .B(n3884), .Z(n3890) );
  HS65_LH_IVX2 U8244 ( .A(n3989), .Z(n3990) );
  HS65_LH_NOR2X6 U5312 ( .A(n4690), .B(n4682), .Z(n4691) );
  HS65_LH_IVX2 U3989 ( .A(n4514), .Z(n4432) );
  HS65_LH_IVX7 U5285 ( .A(n4829), .Z(n4253) );
  HS65_LH_NOR2X5 U4755 ( .A(n4818), .B(n4339), .Z(n4342) );
  HS65_LH_NAND2X5 U6317 ( .A(n4743), .B(n4609), .Z(n4134) );
  HS65_LH_CNIVX3 U3588 ( .A(n4571), .Z(n4295) );
  HS65_LH_NOR2X3 U5299 ( .A(n5206), .B(n5240), .Z(n5243) );
  HS65_LH_OAI21X3 U6348 ( .A(n3790), .B(n3789), .C(n4673), .Z(n3791) );
  HS65_LH_NAND2AX7 U7075 ( .A(n3645), .B(n3644), .Z(n3647) );
  HS65_LH_NAND2X5 U3950 ( .A(n4366), .B(n4368), .Z(n3635) );
  HS65_LH_IVX9 U4733 ( .A(n4176), .Z(n4092) );
  HS65_LH_IVX9 U4813 ( .A(n3845), .Z(n3846) );
  HS65_LH_IVX7 U3542 ( .A(n3796), .Z(n3797) );
  HS65_LH_IVX9 U3528 ( .A(n4289), .Z(n5504) );
  HS65_LH_OAI12X3 U5301 ( .A(n4709), .B(n4708), .C(n5131), .Z(n4710) );
  HS65_LL_OAI21X2 U6271 ( .A(n4662), .B(n2776), .C(n4327), .Z(n4328) );
  HS65_LH_IVX9 U3892 ( .A(n5323), .Z(n5324) );
  HS65_LL_OAI21X2 U5243 ( .A(n5499), .B(n4196), .C(n4195), .Z(n4200) );
  HS65_LH_NOR3X4 U5286 ( .A(n3992), .B(n4014), .C(n3986), .Z(n3987) );
  HS65_LH_OAI112X4 U3919 ( .A(n5502), .B(n4564), .C(n3642), .D(n3641), .Z(
        n3657) );
  HS65_LH_NAND2X4 U4343 ( .A(n4090), .B(n3890), .Z(n3892) );
  HS65_LH_IVX7 U3914 ( .A(n3890), .Z(n2808) );
  HS65_LH_OAI21X3 U3903 ( .A(n5499), .B(n4308), .C(n3919), .Z(n3920) );
  HS65_LH_AOI12X2 U5298 ( .A(n4823), .B(n4822), .C(n4821), .Z(n4824) );
  HS65_LH_AOI211X2 U5280 ( .A(n4781), .B(n5252), .C(n4750), .D(n4749), .Z(
        n4752) );
  HS65_LH_NAND2X5 U3648 ( .A(n5199), .B(n5275), .Z(n5278) );
  HS65_LH_CBI4I1X3 U3523 ( .A(n3968), .B(n3967), .C(n3969), .D(n2833), .Z(
        n3988) );
  HS65_LH_NAND2X5 U4370 ( .A(n4774), .B(n4773), .Z(n4817) );
  HS65_LH_NAND2X5 U6224 ( .A(\lte_x_57/B[2] ), .B(n4197), .Z(n4198) );
  HS65_LH_NAND2AX7 U5255 ( .A(n5054), .B(n2834), .Z(n5055) );
  HS65_LL_AOI21X2 U3884 ( .A(n5326), .B(n5325), .C(n5324), .Z(n5380) );
  HS65_LH_NAND2X5 U4334 ( .A(n7327), .B(n4355), .Z(n4356) );
  HS65_LH_NAND2X4 U6301 ( .A(n4673), .B(n3835), .Z(n4159) );
  HS65_LL_NOR2X2 U3383 ( .A(n2810), .B(n3889), .Z(n3891) );
  HS65_LH_NAND2X5 U4324 ( .A(n7325), .B(n4174), .Z(n4182) );
  HS65_LH_OAI21X3 U6963 ( .A(n4948), .B(n4630), .C(n4198), .Z(n4199) );
  HS65_LH_NAND2X4 U4366 ( .A(n7325), .B(n3764), .Z(n3773) );
  HS65_LH_NAND2X4 U5224 ( .A(n4712), .B(n4706), .Z(n4715) );
  HS65_LH_NAND3X5 U4341 ( .A(n4320), .B(n4319), .C(n4318), .Z(n4359) );
  HS65_LH_AOI22X4 U4355 ( .A(n4743), .B(n4739), .C(n4830), .D(n4672), .Z(n3550) );
  HS65_LH_NOR3X4 U5209 ( .A(n4504), .B(n4503), .C(n4502), .Z(n4505) );
  HS65_LH_OAI12X3 U6207 ( .A(n3669), .B(n4273), .C(n3668), .Z(n3670) );
  HS65_LH_OAI211X5 U3886 ( .A(n4812), .B(n4737), .C(n2827), .D(n2832), .Z(
        n4358) );
  HS65_LH_NOR3X3 U4301 ( .A(n4124), .B(n4123), .C(n4122), .Z(n4143) );
  HS65_LH_NAND2X7 U5190 ( .A(n7325), .B(n4736), .Z(n4762) );
  HS65_LL_AOI21X2 U4168 ( .A(n5486), .B(n4045), .C(n4044), .Z(n4053) );
  HS65_LH_NAND2X5 U4684 ( .A(n7325), .B(n4495), .Z(n4496) );
  HS65_LH_NAND2X5 U4309 ( .A(n7325), .B(n3282), .Z(n3307) );
  HS65_LH_AOI211X3 U3881 ( .A(n4667), .B(n4567), .C(n4566), .D(n4565), .Z(
        n4588) );
  HS65_LL_OAI21X2 U5216 ( .A(n2776), .B(n4624), .C(n4227), .Z(n4391) );
  HS65_LL_AOI21X3 U5175 ( .A(n4774), .B(n4145), .C(n4144), .Z(n8354) );
  HS65_LH_NAND2X5 U4084 ( .A(n5492), .B(n4532), .Z(n4538) );
  HS65_LH_IVX9 U4310 ( .A(n4234), .Z(n4235) );
  HS65_LH_CNIVX3 U9393 ( .A(Data_out_fromRAM[16]), .Z(n8187) );
  HS65_LH_CNIVX3 U9390 ( .A(Data_out_fromRAM[18]), .Z(n8242) );
  HS65_LH_IVX7 U4669 ( .A(Data_out_fromRAM[27]), .Z(n8216) );
  HS65_LH_IVX7 U4671 ( .A(Data_out_fromRAM[24]), .Z(n8231) );
  HS65_LL_AOI21X2 U6579 ( .A(n8800), .B(n8731), .C(n8621), .Z(n7985) );
  HS65_LH_IVX4 U7580 ( .A(n8692), .Z(n3163) );
  HS65_LH_IVX7 U4173 ( .A(n8699), .Z(n8407) );
  HS65_LH_CNIVX7 U6527 ( .A(n8644), .Z(\u_DataPath/jump_address_i [23]) );
  HS65_LH_IVX7 U5064 ( .A(n8694), .Z(n3131) );
  HS65_LHS_XNOR2X6 U7450 ( .A(n8811), .B(n9061), .Z(n6489) );
  HS65_LH_CNIVX7 U7567 ( .A(\u_DataPath/from_mem_data_out_i [3]), .Z(n2981) );
  HS65_LHS_XNOR2X6 U7455 ( .A(n9464), .B(n9058), .Z(n6487) );
  HS65_LH_IVX4 U5156 ( .A(\u_DataPath/dataOut_exe_i [17]), .Z(n3130) );
  HS65_LH_NAND2X5 U4576 ( .A(n8890), .B(n5613), .Z(n5550) );
  HS65_LHS_XNOR2X3 U6774 ( .A(n8944), .B(n5713), .Z(\u_DataPath/toPC2_i [3])
         );
  HS65_LH_IVX4 U4660 ( .A(\u_DataPath/dataOut_exe_i [23]), .Z(n3161) );
  HS65_LH_IVX7 U3929 ( .A(n8296), .Z(\u_DataPath/dataOut_exe_i [3]) );
  HS65_LH_IVX9 U6049 ( .A(\u_DataPath/from_mem_data_out_i [4]), .Z(n2941) );
  HS65_LH_IVX4 U4588 ( .A(n8245), .Z(n2924) );
  HS65_LH_NOR2X6 U5832 ( .A(n8748), .B(n3178), .Z(n3015) );
  HS65_LH_NOR2X5 U6752 ( .A(\u_DataPath/dataOut_exe_i [28]), .B(n3980), .Z(
        n3119) );
  HS65_LL_IVX27 U3910 ( .A(\u_DataPath/cw_to_ex_i [14]), .Z(n3090) );
  HS65_LHS_XNOR2X3 U6762 ( .A(n8920), .B(n5705), .Z(\u_DataPath/toPC2_i [4])
         );
  HS65_LL_NOR2X3 U5984 ( .A(\u_DataPath/dataOut_exe_i [0]), .B(n8045), .Z(
        n3565) );
  HS65_LH_IVX7 U3880 ( .A(n5793), .Z(n5884) );
  HS65_LL_OAI12X3 U4550 ( .A(n5752), .B(n5793), .C(n5751), .Z(n5924) );
  HS65_LL_NAND2X7 U4891 ( .A(n7961), .B(n8000), .Z(\u_DataPath/cw_to_ex_i [2])
         );
  HS65_LH_NAND2X4 U5033 ( .A(n3090), .B(n8402), .Z(n3019) );
  HS65_LH_CNIVX3 U5013 ( .A(n2712), .Z(n3137) );
  HS65_LH_NOR2X6 U3650 ( .A(n8628), .B(n3181), .Z(n3052) );
  HS65_LH_NAND2X5 U6726 ( .A(n8245), .B(n2712), .Z(n2921) );
  HS65_LHS_XNOR2X3 U8538 ( .A(n8926), .B(n5686), .Z(\u_DataPath/toPC2_i [10])
         );
  HS65_LH_NOR2X6 U7297 ( .A(n3019), .B(n8400), .Z(n3020) );
  HS65_LH_NAND2X4 U5950 ( .A(n3184), .B(n9436), .Z(n3012) );
  HS65_LH_NAND2X7 U5953 ( .A(n3184), .B(n9452), .Z(n3062) );
  HS65_LH_NAND2X5 U4609 ( .A(n3184), .B(n9360), .Z(n3043) );
  HS65_LH_CNIVX3 U8438 ( .A(n7329), .Z(n8397) );
  HS65_LH_NAND2X7 U4991 ( .A(n2932), .B(n8392), .Z(n2934) );
  HS65_LL_IVX9 U5523 ( .A(n4533), .Z(\lte_x_57/B[29] ) );
  HS65_LHS_XOR2X3 U5005 ( .A(n8930), .B(n5587), .Z(\u_DataPath/toPC2_i [12])
         );
  HS65_LH_IVX4 U4601 ( .A(n2976), .Z(n2975) );
  HS65_LH_NOR2X5 U3614 ( .A(n3091), .B(n2794), .Z(n3092) );
  HS65_LL_IVX9 U4843 ( .A(n5082), .Z(n2786) );
  HS65_LH_IVX7 U5638 ( .A(n8436), .Z(n3183) );
  HS65_LH_NOR2X6 U5642 ( .A(n3132), .B(n8423), .Z(n3133) );
  HS65_LH_IVX4 U5643 ( .A(n5934), .Z(n8386) );
  HS65_LL_NOR2X5 U6800 ( .A(n3240), .B(n3245), .Z(n3587) );
  HS65_LL_OAI211X3 U4116 ( .A(n8224), .B(n8456), .C(n7314), .D(n7313), .Z(
        n8219) );
  HS65_LH_IVX9 U3816 ( .A(\lte_x_57/B[6] ), .Z(n3951) );
  HS65_LH_AOI22X3 U7974 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][28] ), .B(n9062), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][28] ), .D(
        n8863), .Z(n7584) );
  HS65_LH_IVX7 U3979 ( .A(n5362), .Z(n5028) );
  HS65_LH_NAND2X7 U7148 ( .A(n5393), .B(n5392), .Z(n5361) );
  HS65_LH_CNIVX3 U8146 ( .A(n4957), .Z(n4960) );
  HS65_LH_IVX7 U3801 ( .A(n3587), .Z(n3589) );
  HS65_LH_CNIVX3 U4435 ( .A(n5424), .Z(n5425) );
  HS65_LH_NAND2X4 U3415 ( .A(\lte_x_57/B[29] ), .B(n5196), .Z(n4521) );
  HS65_LH_AOI22X3 U6600 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][0] ), .B(n9199), 
        .C(n9198), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][0] ), .Z(n7283)
         );
  HS65_LH_IVX9 U4862 ( .A(n5004), .Z(n5301) );
  HS65_LH_CNIVX7 U3755 ( .A(n5036), .Z(n5332) );
  HS65_LH_IVX4 U4442 ( .A(n5295), .Z(n3985) );
  HS65_LH_NAND2X7 U8781 ( .A(\lte_x_57/B[29] ), .B(n3204), .Z(n5263) );
  HS65_LH_IVX18 U3373 ( .A(n4591), .Z(n7327) );
  HS65_LH_IVX7 U3736 ( .A(n5284), .Z(n3978) );
  HS65_LH_IVX7 U4035 ( .A(n5298), .Z(n3977) );
  HS65_LH_NAND2X7 U6470 ( .A(n3054), .B(n5203), .Z(n5388) );
  HS65_LH_IVX4 U4452 ( .A(n5334), .Z(n5039) );
  HS65_LH_IVX9 U4794 ( .A(n5337), .Z(n5408) );
  HS65_LL_CNBFX14 U3758 ( .A(n3338), .Z(n3322) );
  HS65_LH_IVX4 U4451 ( .A(n4519), .Z(n4520) );
  HS65_LH_NOR3X1 U4412 ( .A(n4794), .B(n5529), .C(n3200), .Z(n4568) );
  HS65_LH_CNIVX3 U8177 ( .A(n5309), .Z(n5310) );
  HS65_LL_NAND2X4 U4453 ( .A(\lte_x_57/B[7] ), .B(n5207), .Z(n5219) );
  HS65_LH_IVX7 U3603 ( .A(n4684), .Z(n4685) );
  HS65_LH_IVX4 U4803 ( .A(n4983), .Z(n4994) );
  HS65_LH_NAND2X7 U8123 ( .A(\lte_x_57/B[15] ), .B(n2788), .Z(n5115) );
  HS65_LH_CNIVX3 U4415 ( .A(n4970), .Z(n4979) );
  HS65_LH_IVX7 U8306 ( .A(n4523), .Z(n4412) );
  HS65_LL_AOI12X2 U4702 ( .A(n8981), .B(n5920), .C(n9299), .Z(n5768) );
  HS65_LH_NAND2X7 U5493 ( .A(\lte_x_57/B[25] ), .B(n5072), .Z(n3418) );
  HS65_LH_IVX7 U4824 ( .A(n5396), .Z(n5030) );
  HS65_LH_OAI22X3 U5454 ( .A(n5312), .B(n5311), .C(n5310), .D(n5437), .Z(n5314) );
  HS65_LH_IVX9 U5441 ( .A(n5097), .Z(n3841) );
  HS65_LH_IVX7 U4379 ( .A(n5281), .Z(n5315) );
  HS65_LH_NAND2X7 U4440 ( .A(n3138), .B(n5186), .Z(n5367) );
  HS65_LH_NOR2X3 U5336 ( .A(n3372), .B(n5193), .Z(n5194) );
  HS65_LH_NAND2X5 U3699 ( .A(n2824), .B(n5064), .Z(n5292) );
  HS65_LH_NAND2X7 U6448 ( .A(\add_x_50/A[19] ), .B(n5246), .Z(n3538) );
  HS65_LH_NAND2X4 U4428 ( .A(n5449), .B(n4636), .Z(n4651) );
  HS65_LH_CNIVX3 U4437 ( .A(n5333), .Z(n5405) );
  HS65_LH_IVX4 U5426 ( .A(n4686), .Z(n3274) );
  HS65_LL_NOR2X2 U6438 ( .A(\lte_x_57/B[11] ), .B(n3075), .Z(n3664) );
  HS65_LH_CNIVX3 U8339 ( .A(n5191), .Z(n3310) );
  HS65_LH_NOR2X6 U4779 ( .A(n5332), .B(n5408), .Z(n5348) );
  HS65_LH_IVX7 U4398 ( .A(n4169), .Z(n4081) );
  HS65_LH_NOR2X6 U3730 ( .A(n4910), .B(n5187), .Z(n5296) );
  HS65_LH_IVX7 U4018 ( .A(n4347), .Z(n4348) );
  HS65_LH_OAI21X3 U4826 ( .A(n4902), .B(n4901), .C(n5437), .Z(n4903) );
  HS65_LH_IVX18 U3375 ( .A(n4846), .Z(n4781) );
  HS65_LH_NOR2X5 U5542 ( .A(n4283), .B(n2829), .Z(n4317) );
  HS65_LH_IVX9 U5356 ( .A(n5426), .Z(n3667) );
  HS65_LH_NOR2X3 U4375 ( .A(n5408), .B(n5407), .Z(n5409) );
  HS65_LH_IVX9 U3599 ( .A(n5003), .Z(n5283) );
  HS65_LH_IVX4 U8279 ( .A(n4864), .Z(n4349) );
  HS65_LH_IVX9 U3594 ( .A(n5027), .Z(n5364) );
  HS65_LH_CBI4I1X5 U5329 ( .A(n5316), .B(n5450), .C(n5451), .D(n5315), .Z(
        n5320) );
  HS65_LH_CNIVX3 U7705 ( .A(n4313), .Z(n4314) );
  HS65_LH_IVX9 U4814 ( .A(n4447), .Z(n3659) );
  HS65_LH_NAND2X5 U8142 ( .A(\add_x_50/A[19] ), .B(n3189), .Z(n5127) );
  HS65_LH_OAI21X3 U7153 ( .A(n4203), .B(n2830), .C(n3682), .Z(n3685) );
  HS65_LH_NAND2X7 U4792 ( .A(n4641), .B(n4637), .Z(n4644) );
  HS65_LH_IVX9 U4405 ( .A(n5297), .Z(n5005) );
  HS65_LH_IVX7 U4457 ( .A(n3741), .Z(n3323) );
  HS65_LH_IVX7 U4025 ( .A(n4662), .Z(n3911) );
  HS65_LH_AOI21X6 U4850 ( .A(n3742), .B(\sub_x_51/A[27] ), .C(n3594), .Z(n4118) );
  HS65_LH_CNIVX3 U6145 ( .A(n4951), .Z(n4955) );
  HS65_LH_IVX7 U4805 ( .A(n4950), .Z(n5164) );
  HS65_LH_NOR3X3 U3993 ( .A(n4988), .B(n4987), .C(n4986), .Z(n4989) );
  HS65_LH_CNIVX3 U8164 ( .A(n4204), .Z(n4205) );
  HS65_LH_NAND2X4 U4034 ( .A(n3239), .B(n3742), .Z(n3591) );
  HS65_LH_AOI21X6 U4661 ( .A(\lte_x_57/B[10] ), .B(n3826), .C(n4209), .Z(n4126) );
  HS65_LH_IVX4 U4449 ( .A(n3682), .Z(n3403) );
  HS65_LH_IVX9 U3629 ( .A(n4750), .Z(n4621) );
  HS65_LH_NAND2X5 U6494 ( .A(n5509), .B(n5508), .Z(n5513) );
  HS65_LHS_XNOR2X3 U4038 ( .A(n8986), .B(n5928), .Z(
        \u_DataPath/u_execute/resAdd1_i [28]) );
  HS65_LH_OAI21X2 U4800 ( .A(n5452), .B(n5451), .C(n5450), .Z(n5460) );
  HS65_LH_OAI12X3 U5354 ( .A(n3972), .B(n3971), .C(n3970), .Z(n3973) );
  HS65_LH_NAND3X5 U4769 ( .A(n5039), .B(n5403), .C(n5405), .Z(n5421) );
  HS65_LH_NAND2X5 U3606 ( .A(n7327), .B(n5488), .Z(n5494) );
  HS65_LH_NOR2X6 U4846 ( .A(n3716), .B(n3715), .Z(n3788) );
  HS65_LH_IVX9 U4801 ( .A(n5296), .Z(n5051) );
  HS65_LH_IVX7 U3627 ( .A(n3860), .Z(n3863) );
  HS65_LH_NOR2X5 U4367 ( .A(n3466), .B(n4284), .Z(n3467) );
  HS65_LH_AOI21X2 U8199 ( .A(n4918), .B(n5066), .C(n5433), .Z(n3991) );
  HS65_LH_NAND2X7 U4426 ( .A(n3286), .B(n3584), .Z(n4113) );
  HS65_LH_CNIVX3 U4376 ( .A(n5017), .Z(n5018) );
  HS65_LL_NAND3X5 U5343 ( .A(n4949), .B(n4948), .C(n4947), .Z(n5162) );
  HS65_LH_NOR2X5 U4786 ( .A(n5154), .B(n5075), .Z(n5156) );
  HS65_LH_NOR2X5 U5405 ( .A(n3322), .B(n4621), .Z(n3795) );
  HS65_LH_IVX9 U5328 ( .A(n4171), .Z(n4080) );
  HS65_LH_NAND2X7 U5355 ( .A(n5494), .B(n5493), .Z(n5520) );
  HS65_LH_CNIVX3 U8257 ( .A(n3885), .Z(n3887) );
  HS65_LH_NAND2X5 U6479 ( .A(\u_DataPath/u_execute/A_inALU_i[26] ), .B(n5496), 
        .Z(n3486) );
  HS65_LH_NOR2X6 U6389 ( .A(n5395), .B(n5396), .Z(n5363) );
  HS65_LH_CNIVX3 U4389 ( .A(n4604), .Z(n3356) );
  HS65_LH_IVX9 U4011 ( .A(n3915), .Z(n3344) );
  HS65_LH_IVX7 U4436 ( .A(n3924), .Z(n4322) );
  HS65_LH_IVX9 U4357 ( .A(n4638), .Z(n4400) );
  HS65_LH_AOI22X3 U4752 ( .A(n4781), .B(n5077), .C(n3911), .D(n4850), .Z(n3701) );
  HS65_LH_OAI12X3 U4756 ( .A(n5411), .B(n5410), .C(n5409), .Z(n5432) );
  HS65_LH_CNIVX3 U8787 ( .A(n5394), .Z(n5398) );
  HS65_LH_CNIVX3 U4368 ( .A(n4972), .Z(n4786) );
  HS65_LH_NOR2X6 U5360 ( .A(n2994), .B(n4284), .Z(n3719) );
  HS65_LH_NOR2X5 U4353 ( .A(n4592), .B(n3311), .Z(n3314) );
  HS65_LH_CBI4I1X5 U4773 ( .A(n5460), .B(n5459), .C(n5458), .D(n5457), .Z(
        n5472) );
  HS65_LH_NAND2X7 U4799 ( .A(n3418), .B(n3417), .Z(n3424) );
  HS65_LH_AOI12X3 U7127 ( .A(\lte_x_57/B[10] ), .B(n5496), .C(n4212), .Z(n3459) );
  HS65_LH_AOI112X3 U3608 ( .A(n5367), .B(n5366), .C(n5365), .D(n5364), .Z(
        n5368) );
  HS65_LH_AOI21X2 U8224 ( .A(n5269), .B(n5268), .C(n5267), .Z(n5270) );
  HS65_LL_AOI21X2 U3955 ( .A(n3000), .B(n4862), .C(n2999), .Z(n3001) );
  HS65_LH_OAI21X3 U4815 ( .A(n5420), .B(n5345), .C(n5344), .Z(n5346) );
  HS65_LH_NOR2X6 U4745 ( .A(n4541), .B(n4638), .Z(n4543) );
  HS65_LH_CNIVX3 U3844 ( .A(n3730), .Z(n3731) );
  HS65_LL_OAI21X2 U4720 ( .A(n4644), .B(n4643), .C(n4642), .Z(n4645) );
  HS65_LH_IVX7 U3995 ( .A(n4290), .Z(n4291) );
  HS65_LH_IVX4 U4493 ( .A(n3719), .Z(n4783) );
  HS65_LH_IVX4 U7602 ( .A(n4721), .Z(n4722) );
  HS65_LH_NOR2X6 U5402 ( .A(n4207), .B(n4206), .Z(n4840) );
  HS65_LH_NAND2X7 U5317 ( .A(n5126), .B(n4425), .Z(n4429) );
  HS65_LH_NOR2X3 U3953 ( .A(n4591), .B(n9542), .Z(n3819) );
  HS65_LH_OAI21X3 U4347 ( .A(n5420), .B(n5419), .C(n5418), .Z(n5422) );
  HS65_LH_NAND2X5 U4783 ( .A(n4435), .B(n4434), .Z(n4436) );
  HS65_LH_IVX7 U3922 ( .A(n3326), .Z(n4119) );
  HS65_LH_NOR2X5 U3935 ( .A(n5462), .B(n5435), .Z(n5440) );
  HS65_LH_IVX7 U3578 ( .A(n5293), .Z(n5287) );
  HS65_LH_OAI12X3 U3585 ( .A(n4747), .B(n4468), .C(n3727), .Z(n3728) );
  HS65_LH_IVX7 U4796 ( .A(n4473), .Z(n4511) );
  HS65_LH_CNIVX3 U8155 ( .A(n4914), .Z(n4915) );
  HS65_LH_NAND2X5 U4374 ( .A(n4768), .B(n4185), .Z(n4186) );
  HS65_LH_IVX4 U8296 ( .A(n4477), .Z(n4034) );
  HS65_LH_IVX9 U4399 ( .A(n3916), .Z(n3343) );
  HS65_LH_IVX7 U4499 ( .A(n4038), .Z(n4068) );
  HS65_LH_OAI22X6 U8614 ( .A(n3379), .B(n3103), .C(n4662), .D(n5481), .Z(n3321) );
  HS65_LH_AOI211X3 U3945 ( .A(n5304), .B(n5303), .C(n3374), .D(n5302), .Z(
        n5305) );
  HS65_LH_CNIVX3 U3942 ( .A(n4704), .Z(n4705) );
  HS65_LH_NAND2X5 U5348 ( .A(n4426), .B(n3650), .Z(n3651) );
  HS65_LH_NOR2X5 U5326 ( .A(n4601), .B(n3356), .Z(n3360) );
  HS65_LH_IVX9 U3983 ( .A(n3923), .Z(n4323) );
  HS65_LH_IVX7 U3572 ( .A(n3733), .Z(n3387) );
  HS65_LHS_XOR2X3 U6837 ( .A(n9136), .B(n5668), .Z(\u_DataPath/toPC2_i [30])
         );
  HS65_LH_OAI12X3 U4336 ( .A(n3482), .B(n4619), .C(n4119), .Z(n4031) );
  HS65_LH_IVX2 U3913 ( .A(n3959), .Z(n3967) );
  HS65_LH_CBI4I1X5 U7006 ( .A(n4936), .B(n4935), .C(n4934), .D(n4933), .Z(
        n4937) );
  HS65_LH_AOI12X2 U4737 ( .A(n4342), .B(n4822), .C(n4341), .Z(n4343) );
  HS65_LL_AOI12X3 U3500 ( .A(n3191), .B(n4369), .C(n3190), .Z(n4105) );
  HS65_LH_OAI12X3 U4736 ( .A(n3997), .B(n3996), .C(n3995), .Z(n3998) );
  HS65_LL_NAND2X2 U6259 ( .A(n4294), .B(n4038), .Z(n4042) );
  HS65_LH_IVX9 U3602 ( .A(n4150), .Z(n4057) );
  HS65_LH_OAI22X6 U6263 ( .A(n4747), .B(n4254), .C(n4624), .D(n4253), .Z(n4255) );
  HS65_LH_IVX9 U4765 ( .A(n4831), .Z(n4386) );
  HS65_LH_NAND2X7 U7135 ( .A(n4830), .B(n4567), .Z(n3472) );
  HS65_LH_IVX9 U7018 ( .A(n3454), .Z(n4723) );
  HS65_LH_AOI31X2 U5236 ( .A(n4778), .B(n4777), .C(n4776), .D(n5499), .Z(n4779) );
  HS65_LH_NOR2X5 U4430 ( .A(n4292), .B(n4291), .Z(n4293) );
  HS65_LH_NAND2X7 U3544 ( .A(n4830), .B(n4789), .Z(n4320) );
  HS65_LH_IVX4 U4388 ( .A(n4657), .Z(n4664) );
  HS65_LH_NAND2X5 U6385 ( .A(n3847), .B(n3846), .Z(n3850) );
  HS65_LH_CNIVX3 U4346 ( .A(n5428), .Z(n5402) );
  HS65_LH_NAND2X5 U6339 ( .A(n4610), .B(n4831), .Z(n4117) );
  HS65_LH_IVX2 U8340 ( .A(n4618), .Z(n3334) );
  HS65_LH_NAND2X4 U4731 ( .A(n3999), .B(n3998), .Z(n4000) );
  HS65_LH_NAND2AX7 U5258 ( .A(n3608), .B(n3607), .Z(n3609) );
  HS65_LL_OAI21X2 U5256 ( .A(n5499), .B(n4222), .C(n3597), .Z(n3598) );
  HS65_LH_NOR2X6 U4713 ( .A(n2808), .B(n2809), .Z(n2810) );
  HS65_LL_AOI21X2 U3429 ( .A(n4842), .B(n4478), .C(n3793), .Z(n4430) );
  HS65_LH_OAI112X4 U4717 ( .A(n4564), .B(n4386), .C(n4385), .D(n4384), .Z(
        n4387) );
  HS65_LH_CNIVX3 U4728 ( .A(n4148), .Z(n4156) );
  HS65_LH_NAND2X7 U4377 ( .A(n4740), .B(n4827), .Z(n4133) );
  HS65_LH_IVX9 U3904 ( .A(n4104), .Z(n4706) );
  HS65_LH_OAI21X3 U3900 ( .A(n5499), .B(n4068), .C(n4067), .Z(n4072) );
  HS65_LH_AOI21X2 U5259 ( .A(n5466), .B(n5013), .C(n5054), .Z(n5060) );
  HS65_LH_OAI12X3 U5217 ( .A(n5226), .B(n5225), .C(n5224), .Z(n5242) );
  HS65_LH_AOI12X2 U6984 ( .A(n5505), .B(n5504), .C(n5503), .Z(n5519) );
  HS65_LL_OAI211X1 U5210 ( .A(n4614), .B(n4613), .C(n4612), .D(n4611), .Z(
        n4632) );
  HS65_LH_NAND2X5 U5227 ( .A(n7325), .B(n4265), .Z(n4266) );
  HS65_LH_OAI21X3 U4319 ( .A(n4031), .B(n4784), .C(n4030), .Z(n4036) );
  HS65_LL_IVX4 U6216 ( .A(n3666), .Z(n4273) );
  HS65_LH_NAND2X5 U5218 ( .A(n7327), .B(n4867), .Z(n4868) );
  HS65_LH_AOI12X2 U6989 ( .A(n4704), .B(n4711), .C(n4707), .Z(n4106) );
  HS65_LH_AOI12X2 U4704 ( .A(n3314), .B(n4646), .C(n3313), .Z(n3315) );
  HS65_LL_AOI12X2 U5219 ( .A(n4646), .B(n3208), .C(n3207), .Z(n3209) );
  HS65_LL_NAND2X2 U5228 ( .A(n3666), .B(n3071), .Z(n3085) );
  HS65_LL_AOI12X2 U3762 ( .A(n5484), .B(n3803), .C(n3802), .Z(n3814) );
  HS65_LH_IVX7 U4709 ( .A(n4646), .Z(n4553) );
  HS65_LH_IVX4 U4710 ( .A(n4639), .Z(n4554) );
  HS65_LH_NAND2X5 U5220 ( .A(n7327), .B(n3771), .Z(n3772) );
  HS65_LH_AOI21X4 U3490 ( .A(n4400), .B(n4646), .C(n4399), .Z(n4401) );
  HS65_LH_NAND2X5 U4333 ( .A(n4543), .B(n4639), .Z(n4545) );
  HS65_LH_CNIVX3 U4727 ( .A(n4159), .Z(n4162) );
  HS65_LL_OAI21X2 U7077 ( .A(n4506), .B(n4665), .C(n4505), .Z(n4507) );
  HS65_LH_NAND2X4 U4312 ( .A(n7325), .B(n4451), .Z(n4452) );
  HS65_LL_OAI21X2 U4692 ( .A(n4649), .B(n4714), .C(n4648), .Z(n4650) );
  HS65_LH_IVX9 U5203 ( .A(n4529), .Z(n4530) );
  HS65_LL_OAI21X2 U6947 ( .A(n4545), .B(n4714), .C(n4544), .Z(n4546) );
  HS65_LH_NAND2X7 U3682 ( .A(n5492), .B(n7320), .Z(n4698) );
  HS65_LH_NAND2X7 U4693 ( .A(n7325), .B(n3613), .Z(n3622) );
  HS65_LH_NAND2X7 U3670 ( .A(n7327), .B(n3672), .Z(n3711) );
  HS65_LH_NAND2X5 U4690 ( .A(n4774), .B(n4097), .Z(n4098) );
  HS65_LH_NAND2X5 U3669 ( .A(n7327), .B(n3620), .Z(n3621) );
  HS65_LH_NAND2X7 U6152 ( .A(n4774), .B(n3639), .Z(n3640) );
  HS65_LH_IVX7 U3859 ( .A(n8354), .Z(n4363) );
  HS65_LL_NAND3X2 U7340 ( .A(n8333), .B(n8332), .C(n8331), .Z(n5179) );
  HS65_LH_AOI12X6 U6133 ( .A(n4774), .B(n4397), .C(n4396), .Z(n8335) );
  HS65_LH_CNIVX3 U3862 ( .A(n8356), .Z(n5530) );
  HS65_LH_IVX9 U5544 ( .A(n3160), .Z(\add_x_50/A[23] ) );
  HS65_LH_IVX9 U6622 ( .A(n3128), .Z(n4910) );
  HS65_LH_CNIVX7 U5350 ( .A(n5433), .Z(n5290) );
  HS65_LH_AOI21X2 U3829 ( .A(\lte_x_57/B[10] ), .B(n3742), .C(n3335), .Z(n3926) );
  HS65_LH_AOI21X2 U6474 ( .A(\lte_x_57/B[14] ), .B(n5496), .C(n4204), .Z(n3471) );
  HS65_LH_AOI21X2 U3509 ( .A(\lte_x_57/B[15] ), .B(n3826), .C(n3341), .Z(n3915) );
  HS65_LH_AOI21X2 U4859 ( .A(n4796), .B(\lte_x_57/B[6] ), .C(n3844), .Z(n4127)
         );
  HS65_LH_AOI21X2 U6293 ( .A(n5001), .B(n5000), .C(n4999), .Z(n5466) );
  HS65_LH_AOI21X2 U5276 ( .A(n3841), .B(n4863), .C(n3768), .Z(n3769) );
  HS65_LH_DFPSQX4 clk_r_REG732_S4 ( .D(n5935), .CP(net3007), .SN(n9553), .Q(
        n9343) );
  HS65_LH_AOI21X2 U8366 ( .A(n5507), .B(n4902), .C(n5506), .Z(n4408) );
  HS65_LH_AOI21X2 U6313 ( .A(n4864), .B(n4863), .C(n4862), .Z(n4865) );
  HS65_LH_DFPSQX9 clk_r_REG885_S4 ( .D(n2815), .CP(net3007), .SN(n9553), .Q(
        n9169) );
  HS65_LH_DFPSQX9 clk_r_REG875_S4 ( .D(n8015), .CP(net3007), .SN(n9553), .Q(
        n9221) );
  HS65_LH_DFPSQX9 clk_r_REG872_S4 ( .D(n2817), .CP(net3007), .SN(n9553), .Q(
        n9168) );
  HS65_LH_DFPSQX9 clk_r_REG802_S4 ( .D(n2811), .CP(net3007), .SN(n9553), .Q(
        n9167) );
  HS65_LL_AOI21X2 U5177 ( .A(n7327), .B(n3309), .C(n3308), .Z(n8328) );
  HS65_LH_AOI21X2 U5557 ( .A(n8892), .B(n5721), .C(n9309), .Z(n5560) );
  HS65_LH_DFPRQX9 clk_r_REG788_S4 ( .D(n6015), .CP(net3007), .RN(n9553), .Q(
        n8946) );
  HS65_LH_DFPRQX9 clk_r_REG735_S4 ( .D(n6016), .CP(net3007), .RN(n9553), .Q(
        n8948) );
  HS65_LH_DFPRQX9 clk_r_REG821_S4 ( .D(n6530), .CP(net3007), .RN(n9553), .Q(
        n8939) );
  HS65_LH_DFPRQX9 clk_r_REG854_S4 ( .D(n6499), .CP(net3007), .RN(n9553), .Q(
        n8857) );
  HS65_LH_DFPRQX9 clk_r_REG858_S4 ( .D(n6977), .CP(net3007), .RN(n9553), .Q(
        n8885) );
  HS65_LH_DFPRQX9 clk_r_REG804_S4 ( .D(n6347), .CP(net3007), .RN(n9553), .Q(
        n8933) );
  HS65_LL_NAND3X5 U3449 ( .A(n6486), .B(n6485), .C(n6484), .Z(n7302) );
  HS65_LH_DFPSQX9 clk_r_REG782_S4 ( .D(n6122), .CP(net3007), .SN(n9553), .Q(
        n8863) );
  HS65_LH_DFPSQX9 clk_r_REG783_S4 ( .D(n7500), .CP(net3007), .SN(n9553), .Q(
        n9227) );
  HS65_LH_DFPSQX9 clk_r_REG846_S4 ( .D(n7003), .CP(net3007), .SN(n9553), .Q(
        n8884) );
  HS65_LH_DFPSQX9 clk_r_REG627_S4 ( .D(n7955), .CP(net3007), .SN(n9553), .Q(
        n9063) );
  HS65_LH_BFX9 U3399 ( .A(n6861), .Z(n7719) );
  HS65_LH_DFPSQX9 clk_r_REG728_S4 ( .D(n7967), .CP(net3007), .SN(n9553), .Q(
        n9069) );
  HS65_LL_DFPSQX4 clk_r_REG613_S4 ( .D(n7979), .CP(net3007), .SN(n7677), .Q(
        n9317) );
  HS65_LH_DFPSQX9 clk_r_REG723_S4 ( .D(n8021), .CP(net3007), .SN(n9553), .Q(
        n9076) );
  HS65_LH_AOI21X2 U3370 ( .A(n9036), .B(n5924), .C(n9306), .Z(n5842) );
  HS65_LL_NAND2X2 U3374 ( .A(n3081), .B(n3883), .Z(n3083) );
  HS65_LH_OAI21X2 U3393 ( .A(n4281), .B(n4792), .C(n4280), .Z(n4302) );
  HS65_LH_OAI21X2 U3395 ( .A(n4792), .B(n4791), .C(n4790), .Z(n4810) );
  HS65_LH_OAI22X1 U3396 ( .A(n5481), .B(n4308), .C(n4333), .D(n4792), .Z(n3704) );
  HS65_LH_OAI21X2 U3397 ( .A(n4792), .B(n4840), .C(n4215), .Z(n4231) );
  HS65_LH_NOR2X2 U3400 ( .A(n4792), .B(n4289), .Z(n3855) );
  HS65_LL_OAI21X2 U3401 ( .A(n4820), .B(n4336), .C(n4338), .Z(n3254) );
  HS65_LH_IVX2 U3403 ( .A(n4336), .Z(n4337) );
  HS65_LL_AOI12X2 U3404 ( .A(n5507), .B(n4346), .C(n5506), .Z(n4311) );
  HS65_LL_AOI12X2 U3406 ( .A(n4781), .B(n4346), .C(n4309), .Z(n4310) );
  HS65_LL_OR2X9 U3409 ( .A(n3174), .B(n8373), .Z(n2857) );
  HS65_LL_NAND2X2 U3412 ( .A(n3174), .B(n9135), .Z(n2962) );
  HS65_LL_OAI21X2 U3421 ( .A(n2824), .B(n2829), .C(n3624), .Z(n3691) );
  HS65_LL_NAND2X2 U3422 ( .A(\lte_x_57/B[7] ), .B(n5496), .Z(n3733) );
  HS65_LL_AOI21X2 U3424 ( .A(n2792), .B(\sub_x_51/A[8] ), .C(n3731), .Z(n3732)
         );
  HS65_LL_IVX9 U3426 ( .A(n4203), .Z(\lte_x_57/B[11] ) );
  HS65_LH_OAI21X2 U3430 ( .A(n4171), .B(n2823), .C(n4170), .Z(n4172) );
  HS65_LL_AOI12X2 U3431 ( .A(\sub_x_51/A[20] ), .B(n4208), .C(n3490), .Z(n3491) );
  HS65_LH_AOI22X1 U3433 ( .A(n3128), .B(n4208), .C(\sub_x_51/A[16] ), .D(n5498), .Z(n3404) );
  HS65_LH_NAND2X2 U3434 ( .A(\lte_x_57/B[2] ), .B(n4208), .Z(n4116) );
  HS65_LH_NAND2X2 U3440 ( .A(\sub_x_51/A[22] ), .B(n4208), .Z(n3574) );
  HS65_LH_NAND2X2 U3443 ( .A(\sub_x_51/A[8] ), .B(n4208), .Z(n3463) );
  HS65_LL_NAND2X4 U3450 ( .A(\lte_x_57/B[28] ), .B(n4208), .Z(n3823) );
  HS65_LH_NAND2X2 U3464 ( .A(\lte_x_57/B[15] ), .B(n4208), .Z(n3686) );
  HS65_LH_NAND2X2 U3482 ( .A(\add_x_50/A[23] ), .B(n4208), .Z(n3627) );
  HS65_LH_NAND2X2 U3508 ( .A(\sub_x_51/A[18] ), .B(n4208), .Z(n3573) );
  HS65_LH_NAND2X2 U3521 ( .A(\add_x_50/A[19] ), .B(n4208), .Z(n3624) );
  HS65_LL_AOI21X2 U3529 ( .A(n4260), .B(n3261), .C(n3260), .Z(n4170) );
  HS65_LL_NOR2X2 U3543 ( .A(n5481), .B(n4039), .Z(n3739) );
  HS65_LL_NOR2X5 U3571 ( .A(n3738), .B(n3737), .Z(n4039) );
  HS65_LL_OAI12X6 U3580 ( .A(n8427), .B(n3156), .C(n3155), .Z(n5063) );
  HS65_LL_NAND2X7 U3581 ( .A(n3154), .B(n8428), .Z(n3156) );
  HS65_LH_NOR2X3 U3582 ( .A(\lte_x_57/B[2] ), .B(n2994), .Z(n4770) );
  HS65_LL_NOR2X3 U3583 ( .A(\lte_x_57/B[2] ), .B(n5092), .Z(n4804) );
  HS65_LL_IVX7 U3587 ( .A(\lte_x_57/B[2] ), .Z(n4192) );
  HS65_LH_NAND2X2 U3589 ( .A(n2994), .B(\lte_x_57/B[2] ), .Z(n5214) );
  HS65_LL_NOR2X6 U3605 ( .A(n3138), .B(n3322), .Z(n3741) );
  HS65_LL_NAND2X7 U3618 ( .A(n2918), .B(n9103), .Z(n3018) );
  HS65_LL_NAND2X7 U3637 ( .A(n3033), .B(n3032), .Z(n5201) );
  HS65_LL_NAND2X7 U3653 ( .A(n8394), .B(n3031), .Z(n3032) );
  HS65_LL_NAND2X7 U3666 ( .A(n2981), .B(n9425), .Z(n2982) );
  HS65_LL_NAND2X2 U3683 ( .A(n3899), .B(n4080), .Z(n3608) );
  HS65_LL_IVX9 U3684 ( .A(n3899), .Z(n3259) );
  HS65_LL_NOR2X5 U3694 ( .A(n8343), .B(n3882), .Z(n3939) );
  HS65_LL_OAI21X2 U3701 ( .A(n4270), .B(n4273), .C(n4272), .Z(n4025) );
  HS65_LH_AOI22X1 U3721 ( .A(\sub_x_51/A[21] ), .B(n3826), .C(n2796), .D(
        \add_x_50/A[19] ), .Z(n3384) );
  HS65_LH_NAND2X2 U3764 ( .A(\lte_x_57/B[25] ), .B(n2796), .Z(n3629) );
  HS65_LH_NAND2X2 U3767 ( .A(\sub_x_51/A[16] ), .B(n2796), .Z(n3584) );
  HS65_LL_NAND2X2 U3784 ( .A(\lte_x_57/B[3] ), .B(n2796), .Z(n3806) );
  HS65_LH_NAND2X2 U3792 ( .A(n5192), .B(n2796), .Z(n3575) );
  HS65_LH_NAND2X2 U3799 ( .A(n2780), .B(n2796), .Z(n4114) );
  HS65_LL_NAND2X2 U3810 ( .A(\lte_x_57/B[14] ), .B(n2796), .Z(n3852) );
  HS65_LH_NAND2X2 U3821 ( .A(\sub_x_51/A[20] ), .B(n2796), .Z(n3572) );
  HS65_LL_NAND2X5 U3825 ( .A(\sub_x_51/A[21] ), .B(n2796), .Z(n3625) );
  HS65_LH_NAND3X2 U3827 ( .A(n4225), .B(n5486), .C(n4572), .Z(n4280) );
  HS65_LH_NAND2X2 U3843 ( .A(n4225), .B(n4828), .Z(n4120) );
  HS65_LH_NAND3X2 U3869 ( .A(n5486), .B(n4225), .C(n4477), .Z(n3717) );
  HS65_LH_AOI22X1 U3873 ( .A(n4843), .B(n4225), .C(n5505), .D(n3596), .Z(n3597) );
  HS65_LH_AOI22X1 U3876 ( .A(n4225), .B(n3865), .C(n4671), .D(n4573), .Z(n3648) );
  HS65_LH_NAND2X2 U3889 ( .A(n4225), .B(n3836), .Z(n4148) );
  HS65_LH_OAI21X2 U3891 ( .A(n3713), .B(n3712), .C(n4225), .Z(n3399) );
  HS65_LH_NAND3X2 U3893 ( .A(n4225), .B(n5486), .C(n4573), .Z(n4160) );
  HS65_LH_OAI21X2 U3901 ( .A(n3691), .B(n3690), .C(n4225), .Z(n3626) );
  HS65_LL_AOI22X1 U3907 ( .A(n4225), .B(n4479), .C(n4673), .D(n4466), .Z(n4064) );
  HS65_LL_NAND2X2 U3908 ( .A(n4225), .B(n4066), .Z(n3792) );
  HS65_LL_NAND2X2 U3915 ( .A(n4536), .B(n4225), .Z(n4564) );
  HS65_LH_NAND2X2 U3920 ( .A(\sub_x_51/A[13] ), .B(n5082), .Z(n4078) );
  HS65_LH_NOR2X2 U3921 ( .A(n3065), .B(n5082), .Z(n5362) );
  HS65_LH_NAND2X2 U3923 ( .A(n3065), .B(n5082), .Z(n3961) );
  HS65_LL_AOI21X2 U3926 ( .A(n5082), .B(n4781), .C(n4057), .Z(n4059) );
  HS65_LH_AOI22X1 U3951 ( .A(n4671), .B(n4789), .C(n4842), .D(n4739), .Z(n4676) );
  HS65_LL_AOI21X2 U3952 ( .A(n4842), .B(n4392), .C(n4135), .Z(n4142) );
  HS65_LH_AOI21X2 U3963 ( .A(n4842), .B(n3795), .C(n3721), .Z(n3722) );
  HS65_LH_NAND2X2 U3964 ( .A(n4842), .B(n3696), .Z(n3630) );
  HS65_LH_AOI22X1 U3965 ( .A(n4673), .B(n4290), .C(n4842), .D(n4572), .Z(n3649) );
  HS65_LL_NAND2X2 U3967 ( .A(n4842), .B(n4573), .Z(n3496) );
  HS65_LL_IVX2 U3971 ( .A(n4842), .Z(n2776) );
  HS65_LH_OAI22X1 U3981 ( .A(n3103), .B(n3225), .C(n4901), .D(n2829), .Z(n4509) );
  HS65_LH_OAI21X2 U3982 ( .A(n3065), .B(n3225), .C(n3683), .Z(n3684) );
  HS65_LH_OAI21X2 U3985 ( .A(n3054), .B(n3225), .C(n4205), .Z(n4206) );
  HS65_LH_OAI21X2 U4015 ( .A(n3225), .B(n4910), .C(n3323), .Z(n3324) );
  HS65_LH_OAI21X2 U4020 ( .A(n4910), .B(n3225), .C(n3686), .Z(n3689) );
  HS65_LH_OAI21X2 U4023 ( .A(n5148), .B(n3225), .C(n3396), .Z(n3397) );
  HS65_LH_NOR2X2 U4026 ( .A(n3948), .B(n3225), .Z(n4187) );
  HS65_LH_NOR2X2 U4031 ( .A(n4192), .B(n3225), .Z(n3476) );
  HS65_LL_OAI21X2 U4037 ( .A(n3103), .B(n3225), .C(n3407), .Z(n3713) );
  HS65_LH_NOR2X2 U4045 ( .A(n5385), .B(n3225), .Z(n3859) );
  HS65_LH_NOR2X2 U4077 ( .A(n4283), .B(n3225), .Z(n4209) );
  HS65_LH_NOR2X2 U4091 ( .A(n4032), .B(n3225), .Z(n4313) );
  HS65_LH_NOR2X2 U4100 ( .A(n4871), .B(n3225), .Z(n3319) );
  HS65_LH_NOR2X2 U4101 ( .A(n3160), .B(n3225), .Z(n3714) );
  HS65_LL_NOR2X2 U4117 ( .A(n3993), .B(n3225), .Z(n3724) );
  HS65_LL_NOR2X2 U4129 ( .A(n3962), .B(n3225), .Z(n3740) );
  HS65_LL_OAI21X3 U4145 ( .A(n4444), .B(n4448), .C(n4446), .Z(n4376) );
  HS65_LL_NAND2X2 U4158 ( .A(n3128), .B(n5187), .Z(n4446) );
  HS65_LL_NOR2X5 U4170 ( .A(n5187), .B(n3128), .Z(n4444) );
  HS65_LL_NAND2X14 U4221 ( .A(n4870), .B(n9538), .Z(n3338) );
  HS65_LL_NAND2X7 U4297 ( .A(n3221), .B(n3220), .Z(n4870) );
  HS65_LL_OAI12X12 U4321 ( .A(n2963), .B(n2857), .C(n2962), .Z(n9538) );
  HS65_LH_NAND2AX4 U4339 ( .A(n4170), .B(n3899), .Z(n3610) );
  HS65_LL_OA12X9 U4344 ( .A(n4170), .B(n3265), .C(n3264), .Z(n2860) );
  HS65_LH_NAND2X2 U4345 ( .A(n4691), .B(n4683), .Z(n4694) );
  HS65_LH_IVX2 U4349 ( .A(n4683), .Z(n4580) );
  HS65_LL_NAND2X2 U4352 ( .A(n4577), .B(n4683), .Z(n3422) );
  HS65_LL_NAND2X2 U4359 ( .A(n4525), .B(n4683), .Z(n4526) );
  HS65_LL_NAND2X2 U4410 ( .A(n3277), .B(n4683), .Z(n3279) );
  HS65_LL_NAND2X2 U4421 ( .A(n3360), .B(n4683), .Z(n3362) );
  HS65_LL_NAND2X7 U4422 ( .A(n4414), .B(n4683), .Z(n4416) );
  HS65_LH_IVX7 U4424 ( .A(n7445), .Z(n8196) );
  HS65_LL_OAI21X3 U4427 ( .A(n4813), .B(n4738), .C(n3640), .Z(n7445) );
  HS65_LH_NOR2X6 U4438 ( .A(n5481), .B(n5480), .Z(n5482) );
  HS65_LH_IVX4 U4448 ( .A(n4500), .Z(n4501) );
  HS65_LH_IVX7 U4456 ( .A(n4832), .Z(n4224) );
  HS65_LH_AOI12X4 U4467 ( .A(n4414), .B(n4692), .C(n4413), .Z(n4415) );
  HS65_LL_AOI21X2 U4498 ( .A(n5517), .B(n3579), .C(n3578), .Z(n3599) );
  HS65_LH_NAND2X4 U4510 ( .A(n5076), .B(n5156), .Z(n5160) );
  HS65_LH_AOI12X2 U4516 ( .A(n4175), .B(n4092), .C(n4091), .Z(n4093) );
  HS65_LH_IVX7 U4520 ( .A(n4863), .Z(n3002) );
  HS65_LH_IVX7 U4583 ( .A(n4092), .Z(n2809) );
  HS65_LH_NAND2X7 U4657 ( .A(n5434), .B(n3157), .Z(n3637) );
  HS65_LHS_XNOR2X6 U4672 ( .A(n9108), .B(n5674), .Z(\u_DataPath/toPC2_i [29])
         );
  HS65_LH_IVX7 U4683 ( .A(n4689), .Z(n4413) );
  HS65_LH_IVX7 U4686 ( .A(n3455), .Z(n4729) );
  HS65_LH_NAND2X4 U4687 ( .A(n3886), .B(n5394), .Z(n5029) );
  HS65_LH_NOR2X6 U4706 ( .A(n3985), .B(n5283), .Z(n5250) );
  HS65_LH_OAI12X6 U4712 ( .A(n8979), .B(n5560), .C(n9037), .Z(n5674) );
  HS65_LH_IVX7 U4718 ( .A(n5502), .Z(n5511) );
  HS65_LH_NAND2X7 U4719 ( .A(n3128), .B(n3187), .Z(n5244) );
  HS65_LH_NOR3X4 U4721 ( .A(n5316), .B(n4998), .C(n4931), .Z(n4904) );
  HS65_LH_NAND2X7 U4723 ( .A(n3777), .B(n3776), .Z(n3778) );
  HS65_LH_IVX7 U4726 ( .A(n3875), .Z(n3761) );
  HS65_LH_NAND2X7 U4732 ( .A(n5452), .B(n5450), .Z(n5280) );
  HS65_LH_IVX7 U4747 ( .A(n5299), .Z(n5285) );
  HS65_LH_NAND2X7 U4757 ( .A(n4997), .B(n4552), .Z(n5006) );
  HS65_LH_IVX7 U4772 ( .A(n4846), .Z(n5509) );
  HS65_LH_IVX7 U4774 ( .A(n5449), .Z(n5313) );
  HS65_LH_NAND2X7 U4817 ( .A(n2793), .B(n5203), .Z(n4169) );
  HS65_LH_IVX9 U4822 ( .A(n5077), .Z(n3075) );
  HS65_LH_NOR2X5 U4831 ( .A(\lte_x_57/B[15] ), .B(n2788), .Z(n5085) );
  HS65_LH_CNIVX7 U4832 ( .A(n5089), .Z(n2998) );
  HS65_LH_IVX7 U4833 ( .A(n3963), .Z(n3960) );
  HS65_LH_AO22X9 U4836 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][0] ), .B(n9206), 
        .C(n9205), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][0] ), .Z(n7282)
         );
  HS65_LH_IVX7 U4837 ( .A(n4774), .Z(n4591) );
  HS65_LH_NAND2X7 U4838 ( .A(n3975), .B(n5190), .Z(n5450) );
  HS65_LH_AOI22X3 U4857 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][31] ), .B(n9204), 
        .C(n9203), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][31] ), .Z(n7498)
         );
  HS65_LH_NOR2X6 U4867 ( .A(n9293), .B(n7633), .Z(n7307) );
  HS65_LH_NOR2X6 U4869 ( .A(n5079), .B(n3039), .Z(n4046) );
  HS65_LH_NAND2X7 U4880 ( .A(n9043), .B(n7311), .Z(n8037) );
  HS65_LH_NAND2X7 U4890 ( .A(n9043), .B(n7311), .Z(n2820) );
  HS65_LH_IVX7 U4903 ( .A(n3150), .Z(n3151) );
  HS65_LH_IVX7 U4910 ( .A(n8379), .Z(n2993) );
  HS65_LH_IVX7 U4918 ( .A(n2813), .Z(n8165) );
  HS65_LH_NOR3X4 U4936 ( .A(n6495), .B(n6494), .C(n6493), .Z(n6496) );
  HS65_LH_NAND2X7 U4941 ( .A(n9294), .B(n2797), .Z(n8388) );
  HS65_LH_NAND2X7 U4943 ( .A(n9407), .B(n2797), .Z(n8424) );
  HS65_LH_IVX7 U4945 ( .A(n5611), .Z(n5682) );
  HS65_LH_NAND2X7 U4947 ( .A(n9353), .B(n6758), .Z(n7635) );
  HS65_LH_BFX18 U4948 ( .A(n8528), .Z(Address_toRAM[16]) );
  HS65_LH_BFX18 U4958 ( .A(n8527), .Z(Address_toRAM[17]) );
  HS65_LH_BFX18 U4969 ( .A(n8529), .Z(Address_toRAM[0]) );
  HS65_LH_BFX18 U5002 ( .A(n9566), .Z(Address_toRAM[27]) );
  HS65_LH_BFX18 U5034 ( .A(n3534), .Z(Address_toRAM[29]) );
  HS65_LL_NAND2X14 U5049 ( .A(n3564), .B(n9456), .Z(n3450) );
  HS65_LH_IVX7 U5061 ( .A(n3028), .Z(n2961) );
  HS65_LL_NAND2X5 U5172 ( .A(\u_DataPath/dataOut_exe_i [0]), .B(n9115), .Z(
        n8164) );
  HS65_LH_IVX7 U5181 ( .A(n7973), .Z(n7994) );
  HS65_LH_NAND2X7 U5188 ( .A(n9416), .B(n7437), .Z(n7641) );
  HS65_LH_NAND2X7 U5213 ( .A(n6492), .B(n6491), .Z(n6493) );
  HS65_LHS_XNOR2X3 U5235 ( .A(n9213), .B(n7433), .Z(
        \u_DataPath/u_execute/link_value_i [13]) );
  HS65_LL_BFX27 U5239 ( .A(n3439), .Z(n3567) );
  HS65_LH_IVX2 U5241 ( .A(n9565), .Z(n8688) );
  HS65_LH_NOR2X6 U5244 ( .A(n9295), .B(n9075), .Z(n7305) );
  HS65_LH_IVX7 U5247 ( .A(n8684), .Z(\u_DataPath/jump_address_i [18]) );
  HS65_LH_NOR2X6 U5265 ( .A(n8980), .B(n9005), .Z(n5613) );
  HS65_LH_IVX7 U5267 ( .A(n8664), .Z(\u_DataPath/dataOut_exe_i [6]) );
  HS65_LH_CNIVX3 U5288 ( .A(Data_out_fromRAM[20]), .Z(n8291) );
  HS65_LH_AOI21X6 U5291 ( .A(n4774), .B(n4635), .C(n4634), .Z(n8334) );
  HS65_LH_NAND2X7 U5307 ( .A(n4762), .B(n4761), .Z(n4763) );
  HS65_LH_NAND2X7 U5311 ( .A(n4817), .B(n4816), .Z(n8323) );
  HS65_LH_NAND2X5 U5314 ( .A(n7327), .B(n4180), .Z(n4181) );
  HS65_LL_NAND3AX3 U5315 ( .A(n3704), .B(n3703), .C(n3702), .Z(n3705) );
  HS65_LH_NAND3X5 U5316 ( .A(n4159), .B(n4148), .C(n3838), .Z(n3839) );
  HS65_LH_NOR3X4 U5351 ( .A(n3922), .B(n3921), .C(n3920), .Z(n3933) );
  HS65_LH_AOI22X4 U5366 ( .A(n4610), .B(n4827), .C(n4740), .D(n4609), .Z(n4611) );
  HS65_LH_CNIVX3 U5377 ( .A(n4466), .Z(n3392) );
  HS65_LH_NAND2X5 U5392 ( .A(n4667), .B(n4382), .Z(n4110) );
  HS65_LH_IVX4 U5406 ( .A(n4382), .Z(n4623) );
  HS65_LH_OAI12X3 U5408 ( .A(n4917), .B(n4916), .C(n4915), .Z(n4925) );
  HS65_LH_AOI12X6 U5409 ( .A(n8893), .B(n5674), .C(n9304), .Z(n5668) );
  HS65_LH_NAND2X5 U5438 ( .A(n3384), .B(n3383), .Z(n4473) );
  HS65_LH_NAND2X7 U5442 ( .A(n4126), .B(n4125), .Z(n4609) );
  HS65_LH_NAND3X5 U5443 ( .A(n3830), .B(n3829), .C(n3828), .Z(n4569) );
  HS65_LH_NOR2X5 U5447 ( .A(n5011), .B(n5010), .Z(n5017) );
  HS65_LH_NOR2X6 U5448 ( .A(\lte_x_57/B[25] ), .B(n5072), .Z(n3416) );
  HS65_LH_NAND2X5 U5470 ( .A(n4720), .B(n4719), .Z(n4735) );
  HS65_LH_NAND2X5 U5474 ( .A(n4521), .B(n4520), .Z(n4531) );
  HS65_LH_CNIVX3 U5480 ( .A(n4945), .Z(n4949) );
  HS65_LH_NOR2X5 U5482 ( .A(n4533), .B(n5196), .Z(n5011) );
  HS65_LH_NOR2X6 U5494 ( .A(\sub_x_51/A[13] ), .B(n2786), .Z(n5391) );
  HS65_LH_NAND2X5 U5515 ( .A(\lte_x_57/B[30] ), .B(n5312), .Z(n4684) );
  HS65_LH_NAND2X7 U5517 ( .A(\lte_x_57/B[14] ), .B(n5392), .Z(n3901) );
  HS65_LH_OAI22X4 U5528 ( .A(n3163), .B(n2794), .C(n8650), .D(n2772), .Z(n8442) );
  HS65_LL_CBI4I6X5 U5551 ( .A(n7214), .B(n7213), .C(n7212), .D(n8778), .Z(
        n7311) );
  HS65_LH_IVX4 U5554 ( .A(n5279), .Z(n5527) );
  HS65_LL_BFX9 U5577 ( .A(n3450), .Z(n3568) );
  HS65_LH_NAND2X5 U5586 ( .A(n8700), .B(n2712), .Z(n3045) );
  HS65_LH_CNIVX27 U5590 ( .A(n8164), .Z(nibble[0]) );
  HS65_LH_NAND3X5 U5598 ( .A(n8806), .B(n7414), .C(n9052), .Z(n7978) );
  HS65_LH_NOR2X5 U5606 ( .A(\u_DataPath/dataOut_exe_i [22]), .B(n3178), .Z(
        n3167) );
  HS65_LH_NOR2X5 U5611 ( .A(\u_DataPath/dataOut_exe_i [21]), .B(n3980), .Z(
        n8435) );
  HS65_LH_NOR2X5 U5616 ( .A(n8646), .B(n2772), .Z(n8385) );
  HS65_LH_NOR2X5 U5619 ( .A(\u_DataPath/dataOut_exe_i [19]), .B(n3178), .Z(
        n3147) );
  HS65_LH_IVX4 U5621 ( .A(n7414), .Z(n7963) );
  HS65_LH_NOR2X5 U5627 ( .A(n8553), .B(n3980), .Z(n8420) );
  HS65_LH_NAND3X5 U5647 ( .A(n7348), .B(n8845), .C(n7346), .Z(n7349) );
  HS65_LH_IVX4 U5648 ( .A(n9564), .Z(n8707) );
  HS65_LL_AND2ABX18 U5652 ( .A(n9115), .B(n8454), .Z(n3439) );
  HS65_LH_OAI12X3 U5654 ( .A(n8911), .B(n5847), .C(n8776), .Z(n5775) );
  HS65_LH_IVX4 U5657 ( .A(n8691), .Z(n3173) );
  HS65_LH_IVX4 U5667 ( .A(n8717), .Z(n3142) );
  HS65_LH_NOR2X5 U5668 ( .A(n8747), .B(n2782), .Z(n8375) );
  HS65_LH_NOR2X5 U5671 ( .A(n9084), .B(n9403), .Z(n7441) );
  HS65_LH_IVX4 U5672 ( .A(Data_out_fromRAM[25]), .Z(n8260) );
  HS65_LH_AOI21X6 U5673 ( .A(n7327), .B(n4424), .C(n4423), .Z(n8333) );
  HS65_LH_NAND2X4 U5676 ( .A(n4774), .B(n3895), .Z(n3938) );
  HS65_LL_OAI21X2 U5679 ( .A(n4967), .B(n4630), .C(n4629), .Z(n4631) );
  HS65_LH_AOI22X3 U5680 ( .A(n5510), .B(n4741), .C(n4740), .D(n4739), .Z(n4757) );
  HS65_LH_NAND2X4 U5681 ( .A(n5492), .B(n4087), .Z(n4088) );
  HS65_LH_OA12X9 U5686 ( .A(n5481), .B(n4791), .C(n4335), .Z(n2832) );
  HS65_LH_NAND2X4 U5687 ( .A(n4704), .B(n4706), .Z(n4107) );
  HS65_LH_AOI22X3 U5690 ( .A(n4743), .B(n4827), .C(n4667), .D(n4609), .Z(n4390) );
  HS65_LH_AO22X9 U5692 ( .A(n4830), .B(n4479), .C(n4667), .D(n4466), .Z(n4443)
         );
  HS65_LH_NAND2X4 U5693 ( .A(n5511), .B(n4667), .Z(n4286) );
  HS65_LHS_XOR2X6 U5699 ( .A(n4866), .B(n4865), .Z(n4867) );
  HS65_LHS_XNOR2X6 U5701 ( .A(n4278), .B(n2823), .Z(n9544) );
  HS65_LH_NAND2X4 U5702 ( .A(n4830), .B(n3390), .Z(n4043) );
  HS65_LH_OAI12X3 U5704 ( .A(n4659), .B(n4468), .C(n3799), .Z(n3800) );
  HS65_LH_NOR2X3 U5708 ( .A(n4468), .B(n4564), .Z(n4437) );
  HS65_LH_NAND2X4 U5710 ( .A(n5505), .B(n4572), .Z(n4153) );
  HS65_LH_NAND2AX7 U5711 ( .A(n3405), .B(n3404), .Z(n4480) );
  HS65_LH_OAI22X3 U5716 ( .A(n4747), .B(n3349), .C(n4657), .D(n4659), .Z(n3350) );
  HS65_LH_NAND3X3 U5723 ( .A(n5367), .B(n5288), .C(n5250), .Z(n3986) );
  HS65_LH_NOR2X5 U5727 ( .A(n3275), .B(n4682), .Z(n3277) );
  HS65_LH_NAND2X4 U5730 ( .A(n3736), .B(n3735), .Z(n3737) );
  HS65_LH_CNIVX3 U5731 ( .A(n5363), .Z(n5369) );
  HS65_LH_OAI21X3 U5733 ( .A(n3962), .B(n3322), .C(n3852), .Z(n3853) );
  HS65_LH_OAI21X3 U5735 ( .A(n4192), .B(n3322), .C(n3806), .Z(n3389) );
  HS65_LL_NOR2AX3 U5743 ( .A(n3203), .B(n3202), .Z(n4643) );
  HS65_LL_NOR2X6 U5746 ( .A(n4147), .B(n4613), .Z(n4830) );
  HS65_LH_CNIVX3 U5747 ( .A(n4239), .Z(n4240) );
  HS65_LH_NAND2X4 U5755 ( .A(n4801), .B(n4800), .Z(n4806) );
  HS65_LH_OAI21X3 U5757 ( .A(n3962), .B(n3322), .C(n3573), .Z(n4112) );
  HS65_LH_AO22X9 U5775 ( .A(n2780), .B(n2792), .C(\lte_x_57/B[3] ), .D(n4796), 
        .Z(n2855) );
  HS65_LH_NAND2X4 U5778 ( .A(n4578), .B(n4577), .Z(n4582) );
  HS65_LH_OAI21X3 U5788 ( .A(n5455), .B(n5454), .C(n5453), .Z(n5458) );
  HS65_LH_NAND2X4 U5790 ( .A(\lte_x_57/B[30] ), .B(n2790), .Z(n5145) );
  HS65_LL_NOR2X6 U5809 ( .A(n2946), .B(n2945), .Z(\lte_x_57/B[4] ) );
  HS65_LH_NAND3X3 U5820 ( .A(n5329), .B(n5328), .C(n5327), .Z(n5330) );
  HS65_LH_IVX9 U5828 ( .A(n2824), .Z(\sub_x_51/A[20] ) );
  HS65_LL_NOR2X6 U5830 ( .A(n4879), .B(n4877), .Z(\lte_x_57/B[6] ) );
  HS65_LH_AOI12X2 U5837 ( .A(n9087), .B(n5682), .C(n8711), .Z(n5627) );
  HS65_LHS_XNOR2X6 U5840 ( .A(n9088), .B(n5701), .Z(\u_DataPath/toPC2_i [7])
         );
  HS65_LHS_XNOR2X6 U5852 ( .A(n9007), .B(n5896), .Z(
        \u_DataPath/u_execute/resAdd1_i [9]) );
  HS65_LH_IVX9 U5867 ( .A(n3065), .Z(\sub_x_51/A[13] ) );
  HS65_LH_OAI21X3 U5920 ( .A(n8635), .B(n3181), .C(n3013), .Z(n3014) );
  HS65_LH_AOI12X2 U5968 ( .A(n9342), .B(n5813), .C(n9271), .Z(n5815) );
  HS65_LH_NOR2X3 U6134 ( .A(\u_DataPath/cw_to_ex_i [0]), .B(
        \u_DataPath/cw_to_ex_i [1]), .Z(n5279) );
  HS65_LH_CNIVX3 U6151 ( .A(n2797), .Z(n7646) );
  HS65_LH_NAND2X4 U6179 ( .A(n8721), .B(n2712), .Z(n3086) );
  HS65_LH_AOI211X4 U6214 ( .A(n8816), .B(n8585), .C(n7953), .D(n8743), .Z(
        n7961) );
  HS65_LH_AOI12X2 U6220 ( .A(n8890), .B(n5612), .C(n9300), .Z(n5549) );
  HS65_LHS_XOR2X6 U6223 ( .A(n9212), .B(n7622), .Z(
        \u_DataPath/u_execute/link_value_i [9]) );
  HS65_LH_NOR2X3 U6241 ( .A(n8817), .B(n8802), .Z(n7414) );
  HS65_LHS_XOR2X6 U6246 ( .A(n9343), .B(n9410), .Z(n7205) );
  HS65_LHS_XNOR2X6 U6248 ( .A(n9410), .B(n9169), .Z(n7201) );
  HS65_LH_NAND2X4 U6258 ( .A(n9412), .B(n2782), .Z(n2959) );
  HS65_LH_AOI22X4 U6276 ( .A(n8687), .B(n9053), .C(n9252), .D(n9117), .Z(n8241) );
  HS65_LH_NAND3X6 U6290 ( .A(n9209), .B(n9225), .C(n9334), .Z(n3532) );
  HS65_LH_IVX2 U6302 ( .A(n5042), .Z(n5416) );
  HS65_LH_NAND2X4 U6307 ( .A(n3090), .B(n8413), .Z(n3068) );
  HS65_LH_NAND2X2 U6372 ( .A(\lte_x_57/B[6] ), .B(n4208), .Z(n4211) );
  HS65_LH_IVX2 U6418 ( .A(n5403), .Z(n5411) );
  HS65_LH_OAI21X2 U6423 ( .A(n5115), .B(n4427), .C(n4426), .Z(n5116) );
  HS65_LH_NOR2X2 U6440 ( .A(n5141), .B(n5191), .Z(n5143) );
  HS65_LH_NAND2X2 U6444 ( .A(n4871), .B(n9538), .Z(n5417) );
  HS65_LH_NOR2X3 U6451 ( .A(n5392), .B(n5393), .Z(n5360) );
  HS65_LH_AOI21X2 U6456 ( .A(n5135), .B(n5134), .C(n5133), .Z(n5136) );
  HS65_LH_NOR2X2 U6462 ( .A(n5294), .B(n5002), .Z(n4912) );
  HS65_LH_IVX2 U6492 ( .A(n5336), .Z(n4894) );
  HS65_LHS_XNOR2X3 U6495 ( .A(n4032), .B(n5079), .Z(n4985) );
  HS65_LH_IVX2 U6498 ( .A(n4658), .Z(n4661) );
  HS65_LHS_XNOR2X3 U6499 ( .A(n5508), .B(n2774), .Z(n5516) );
  HS65_LH_AOI21X2 U6511 ( .A(n5402), .B(n5401), .C(n5400), .Z(n5443) );
  HS65_LH_NOR2X2 U6513 ( .A(n4347), .B(n4859), .Z(n5223) );
  HS65_LH_NAND4ABX6 U6532 ( .A(n4979), .B(n4978), .C(n4977), .D(n4976), .Z(
        n4980) );
  HS65_LH_AOI21X2 U6535 ( .A(n5231), .B(n5230), .C(n5229), .Z(n5239) );
  HS65_LH_AO22X4 U6544 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][8] ), .B(n9470), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][8] ), .D(n9267), .Z(n6658) );
  HS65_LH_AOI22X1 U6584 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][8] ), .B(n9191), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][8] ), .D(
        n9471), .Z(n6651) );
  HS65_LH_AOI21X2 U6599 ( .A(n4411), .B(n4156), .C(n4155), .Z(n4165) );
  HS65_LH_AOI21X2 U6604 ( .A(n4830), .B(n4664), .C(n4663), .Z(n4669) );
  HS65_LH_CBI4I1X3 U6610 ( .A(n5507), .B(n5246), .C(n5506), .D(
        \add_x_50/A[19] ), .Z(n3545) );
  HS65_LH_AOI21X2 U6638 ( .A(n5517), .B(n4786), .C(n4785), .Z(n4787) );
  HS65_LH_AO22X4 U6644 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][7] ), .B(n9470), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][7] ), .D(n9267), .Z(n6472) );
  HS65_LH_AOI22X1 U6656 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][13] ), .B(n9250), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][13] ), .D(
        n9265), .Z(n7029) );
  HS65_LH_AOI22X1 U6661 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][3] ), .B(n9242), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][3] ), .D(n9166), .Z(n6134) );
  HS65_LH_AOI22X1 U6666 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][11] ), .B(n9242), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][11] ), .D(
        n8861), .Z(n6813) );
  HS65_LH_AOI22X1 U6668 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][26] ), .B(n8938), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][26] ), .D(
        n9264), .Z(n6940) );
  HS65_LH_AOI22X1 U6673 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][26] ), .B(n9191), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][26] ), .D(
        n9471), .Z(n6938) );
  HS65_LH_AO22X4 U6685 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][19] ), .B(n9251), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][19] ), .D(
        n9155), .Z(n6297) );
  HS65_LH_AO22X4 U6714 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][12] ), .B(n9363), 
        .C(n9257), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][12] ), .Z(n7151)
         );
  HS65_LH_AO22X4 U6743 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][24] ), .B(n9249), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][24] ), .D(
        n9185), .Z(n6276) );
  HS65_LH_AO22X4 U6756 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][17] ), .B(n9364), 
        .C(n9068), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][17] ), .Z(n5946)
         );
  HS65_LH_AOI22X1 U6767 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][1] ), .B(n9250), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][1] ), .D(n9265), .Z(n7251) );
  HS65_LH_AOI22X1 U6775 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][1] ), .B(n9247), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][1] ), .D(n9227), .Z(n7246) );
  HS65_LH_AO22X4 U6812 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][14] ), .B(n9470), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][14] ), .D(
        n9164), .Z(n6876) );
  HS65_LH_AO22X4 U6856 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][30] ), .B(n9249), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][30] ), .D(
        n9185), .Z(n6574) );
  HS65_LH_AOI22X1 U6913 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][31] ), .B(n9259), 
        .C(n9256), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][31] ), .Z(n7519)
         );
  HS65_LH_AO22X4 U6932 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][27] ), .B(n9472), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][27] ), .D(
        n8857), .Z(n6309) );
  HS65_LH_AO22X4 U6978 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][29] ), .B(n9470), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][29] ), .D(
        n9267), .Z(n6925) );
  HS65_LH_AOI22X1 U6987 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][29] ), .B(n8950), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][29] ), .D(
        n9471), .Z(n6915) );
  HS65_LH_AOI22X1 U6996 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][25] ), .B(n9188), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][25] ), .D(
        n9190), .Z(n6958) );
  HS65_LH_AOI22X1 U7021 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][12] ), .B(n9188), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][12] ), .D(
        n9190), .Z(n6690) );
  HS65_LH_AO22X4 U7044 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][15] ), .B(n9469), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][15] ), .D(
        n9475), .Z(n6887) );
  HS65_LH_AO22X4 U7067 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][21] ), .B(n9261), 
        .C(n9263), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][21] ), .Z(n6005)
         );
  HS65_LH_AO22X4 U7084 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][9] ), .B(n8939), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][9] ), .D(
        n9186), .Z(n6996) );
  HS65_LH_AO22X4 U7107 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][20] ), .B(n9251), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][20] ), .D(
        n9186), .Z(n6593) );
  HS65_LH_AO22X4 U7137 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][20] ), .B(n9364), 
        .C(n9253), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][20] ), .Z(n7101)
         );
  HS65_LH_AO22X4 U7144 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][5] ), .B(n9251), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][5] ), .D(
        n9155), .Z(n6633) );
  HS65_LH_AO22X4 U7155 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][10] ), .B(n9470), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][10] ), .D(
        n9267), .Z(n6718) );
  HS65_LH_AO22X4 U7164 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][6] ), .B(n9470), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][6] ), .D(n9267), .Z(n6742) );
  HS65_LH_AO22X4 U7167 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][22] ), .B(n9251), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][22] ), .D(
        n9155), .Z(n6553) );
  HS65_LH_AOI22X1 U7183 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][15] ), .B(n9242), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][15] ), .D(
        n9166), .Z(n7270) );
  HS65_LH_AOI22X1 U7225 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][0] ), .B(n9242), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][0] ), .D(n9166), .Z(n7294) );
  HS65_LH_AO22X4 U7227 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][28] ), .B(n8858), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][28] ), .D(
        n9468), .Z(n6521) );
  HS65_LH_AO22X4 U7228 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][31] ), .B(n8858), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][31] ), .D(
        n9468), .Z(n6604) );
  HS65_LH_AOI22X1 U7241 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][5] ), .B(n9247), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][5] ), .D(n9227), .Z(n7084) );
  HS65_LH_AO22X4 U7293 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][9] ), .B(n9363), 
        .C(n9257), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][9] ), .Z(n7071) );
  HS65_LH_AO22X4 U7294 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][29] ), .B(n9254), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][29] ), .D(
        n9244), .Z(n7551) );
  HS65_LH_AO22X4 U7305 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][27] ), .B(n9254), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][27] ), .D(
        n9244), .Z(n7170) );
  HS65_LH_AOI22X1 U7425 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][23] ), .B(n9242), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][23] ), .D(
        n8861), .Z(n7128) );
  HS65_LH_AO22X4 U7566 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][28] ), .B(n9254), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][28] ), .D(
        n9244), .Z(n7581) );
  HS65_LH_AOI22X1 U7572 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][28] ), .B(n9204), 
        .C(n9203), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][28] ), .Z(n7575)
         );
  HS65_LH_AO22X4 U7579 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][30] ), .B(n9208), 
        .C(n9200), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][30] ), .Z(n7528)
         );
  HS65_LH_AO22X4 U7588 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][13] ), .B(n9472), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][13] ), .D(
        n8857), .Z(n6398) );
  HS65_LH_AO22X4 U7603 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][21] ), .B(n9473), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][21] ), .D(
        n9474), .Z(n6377) );
  HS65_LH_AOI22X1 U7613 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][24] ), .B(n9247), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][24] ), .D(
        n9227), .Z(n5982) );
  HS65_LH_AOI22X1 U7622 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][16] ), .B(n9250), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][16] ), .D(
        n9265), .Z(n6073) );
  HS65_LH_AO22X4 U7706 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][16] ), .B(n9364), 
        .C(n9253), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][16] ), .Z(n6065)
         );
  HS65_LH_AOI22X1 U7716 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][17] ), .B(n8950), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][17] ), .D(
        n9471), .Z(n6364) );
  HS65_LH_AOI22X1 U8118 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][23] ), .B(n9188), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][23] ), .D(
        n9190), .Z(n6336) );
  HS65_LH_AOI22X1 U8124 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][11] ), .B(n9188), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][11] ), .D(
        n9190), .Z(n6506) );
  HS65_LH_AO22X4 U8208 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][1] ), .B(n9154), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][1] ), .D(
        n9194), .Z(n6241) );
  HS65_LH_AO22X4 U8210 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][4] ), .B(n9249), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][4] ), .D(
        n8949), .Z(n6428) );
  HS65_LH_AO22X4 U8216 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][16] ), .B(n9251), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][16] ), .D(
        n9186), .Z(n6179) );
  HS65_LH_AO22X4 U8221 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][4] ), .B(n9364), 
        .C(n9253), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][4] ), .Z(n6023)
         );
  HS65_LH_AOI22X1 U8280 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][2] ), .B(n9246), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][2] ), .D(n9262), .Z(n6225) );
  HS65_LH_AO22X4 U8294 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][3] ), .B(n9472), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][3] ), .D(
        n8857), .Z(n6438) );
  HS65_LH_AO22X4 U8344 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][0] ), .B(n9473), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][0] ), .D(
        n9474), .Z(n6197) );
  HS65_LH_AOI22X1 U8354 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][18] ), .B(n9255), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][18] ), .D(
        n9116), .Z(n6666) );
  HS65_LH_AOI22X1 U8358 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][25] ), .B(n9247), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][25] ), .D(
        n9227), .Z(n7484) );
  HS65_LH_AOI22X1 U8392 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][14] ), .B(n9250), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][14] ), .D(
        n9265), .Z(n6093) );
  HS65_LH_NOR2X6 U8412 ( .A(n3817), .B(n2852), .Z(n3818) );
  HS65_LH_HA1X4 U8609 ( .A0(n7638), .B0(n9356), .CO(n7637), .S0(
        \u_DataPath/u_execute/link_value_i [30]) );
  HS65_LH_AND2X4 U8631 ( .A(n7325), .B(n3425), .Z(n3426) );
  HS65_LL_NAND3X2 U8656 ( .A(n4183), .B(n4182), .C(n4181), .Z(n8349) );
  HS65_LH_NAND2X2 U8690 ( .A(\u_DataPath/dataOut_exe_i [1]), .B(nibble[0]), 
        .Z(n8456) );
  HS65_LL_NAND3X2 U8694 ( .A(n3774), .B(n3773), .C(n3772), .Z(n8343) );
  HS65_LH_AOI21X2 U8700 ( .A(n5492), .B(n3552), .C(n3551), .Z(n8324) );
  HS65_LH_BFX35 U8703 ( .A(n8874), .Z(n9536) );
  HS65_LH_BFX35 U8708 ( .A(n8557), .Z(n9530) );
  HS65_LH_BFX35 U8730 ( .A(n8559), .Z(n9532) );
  HS65_LH_BFX35 U8734 ( .A(n8560), .Z(n9533) );
  HS65_LH_BFX35 U8735 ( .A(n8561), .Z(n9534) );
  HS65_LH_BFX35 U8736 ( .A(n8562), .Z(n9535) );
  HS65_LH_BFX35 U8738 ( .A(n8534), .Z(n9510) );
  HS65_LH_BFX35 U8739 ( .A(n8533), .Z(n9509) );
  HS65_LH_BFX35 U8744 ( .A(n8554), .Z(n9527) );
  HS65_LH_BFX35 U8746 ( .A(n8558), .Z(n9531) );
  HS65_LH_BFX35 U8758 ( .A(n8531), .Z(n9507) );
  HS65_LH_BFX35 U8764 ( .A(n8552), .Z(n9526) );
  HS65_LH_BFX35 U8775 ( .A(n8538), .Z(n9514) );
  HS65_LH_BFX35 U8779 ( .A(n8536), .Z(n9512) );
  HS65_LH_BFX35 U8785 ( .A(n8532), .Z(n9508) );
  HS65_LH_BFX35 U8802 ( .A(n8543), .Z(n9519) );
  HS65_LH_BFX35 U8817 ( .A(n8542), .Z(n9518) );
  HS65_LH_BFX35 U8855 ( .A(n8540), .Z(n9516) );
  HS65_LH_BFX35 U8859 ( .A(n8545), .Z(n9521) );
  HS65_LH_BFX35 U8873 ( .A(n8544), .Z(n9520) );
  HS65_LH_BFX35 U8909 ( .A(n8548), .Z(n9522) );
  HS65_LH_BFX35 U8922 ( .A(n8549), .Z(n9523) );
  HS65_LH_BFX35 U8935 ( .A(n8551), .Z(n9525) );
  HS65_LH_BFX35 U8949 ( .A(n8555), .Z(n9528) );
  HS65_LH_BFX35 U8966 ( .A(n8550), .Z(n9524) );
  HS65_LH_BFX35 U8976 ( .A(n8535), .Z(n9511) );
  HS65_LH_BFX35 U8982 ( .A(n8530), .Z(n9506) );
  HS65_LH_BFX35 U8983 ( .A(n8539), .Z(n9515) );
  HS65_LH_BFX35 U8988 ( .A(n8537), .Z(n9513) );
  HS65_LH_BFX35 U8992 ( .A(n8556), .Z(n9529) );
  HS65_LH_BFX35 U8993 ( .A(n8541), .Z(n9517) );
  HS65_LH_NOR2AX3 U8999 ( .A(\u_DataPath/dataOut_exe_i [19]), .B(n3439), .Z(
        n8527) );
  HS65_LH_NOR2AX3 U9028 ( .A(\u_DataPath/dataOut_exe_i [18]), .B(n3439), .Z(
        n8528) );
  HS65_LH_NOR2AX3 U9036 ( .A(\u_DataPath/dataOut_exe_i [31]), .B(n3439), .Z(
        n3534) );
  HS65_LH_NOR2AX3 U9044 ( .A(n8747), .B(n3439), .Z(n8529) );
  HS65_LH_NOR2AX3 U9050 ( .A(\u_DataPath/dataOut_exe_i [29]), .B(n3439), .Z(
        n9566) );
  HS65_LL_NOR2AX25 U9053 ( .A(n8581), .B(n3450), .Z(n3523) );
  HS65_LL_NOR2AX25 U9060 ( .A(n8764), .B(n3567), .Z(n3554) );
  HS65_LL_NOR2AX25 U9063 ( .A(n9119), .B(n3568), .Z(n3446) );
  HS65_LL_NOR2AX25 U9064 ( .A(\u_DataPath/dataOut_exe_i [26]), .B(n3439), .Z(
        n3535) );
endmodule

