
module DLX ( clk, rst, iram_data, Data_out_fromRAM, addr_to_iram, read_op, 
        write_op, nibble, write_byte, Address_toRAM, Data_in );
  input [31:0] iram_data;
  input [31:0] Data_out_fromRAM;
  output [31:0] addr_to_iram;
  output [1:0] nibble;
  output [31:0] Address_toRAM;
  output [31:0] Data_in;
  input clk, rst;
  output read_op, write_op, write_byte;
  wire   n17215, n17216, n17217, n17218, n17219, n17220, n17221, n17222,
         n17223, n17224, n17225, n17226, n17227, n17228, n17229, n17230,
         n17231, n17232, n17233, n17234, n17235, n17236, n17237, n17238,
         n17239, n17240, n17241, n17242, n17243, n17244, write_op_snps_wire,
         \nibble[1]_snps_wire , Address_toRAM_20, Address_toRAM_19,
         Address_toRAM_18, Address_toRAM_17, Address_toRAM_16,
         Address_toRAM_15, Address_toRAM_14, Address_toRAM_13,
         Address_toRAM_12, Address_toRAM_1, Address_toRAM_0, Data_in_26,
         Data_in_25, Data_in_24, Data_in_23, Data_in_6, Data_in_5, Data_in_4,
         Data_in_3, Data_in_2, Data_in_1, Data_in_0,
         \u_DataPath/takeBranch_out_i , \u_DataPath/reg_write_i ,
         \u_DataPath/jump_i , \u_DataPath/u_fetch/pc1/N3 ,
         \u_DataPath/u_ifidreg/N67 , \u_DataPath/u_ifidreg/N66 ,
         \u_DataPath/u_ifidreg/N65 , \u_DataPath/u_ifidreg/N64 ,
         \u_DataPath/u_ifidreg/N63 , \u_DataPath/u_ifidreg/N62 ,
         \u_DataPath/u_ifidreg/N61 , \u_DataPath/u_ifidreg/N60 ,
         \u_DataPath/u_ifidreg/N59 , \u_DataPath/u_ifidreg/N58 ,
         \u_DataPath/u_ifidreg/N57 , \u_DataPath/u_ifidreg/N56 ,
         \u_DataPath/u_ifidreg/N55 , \u_DataPath/u_ifidreg/N54 ,
         \u_DataPath/u_ifidreg/N53 , \u_DataPath/u_ifidreg/N52 ,
         \u_DataPath/u_ifidreg/N51 , \u_DataPath/u_ifidreg/N50 ,
         \u_DataPath/u_ifidreg/N49 , \u_DataPath/u_ifidreg/N48 ,
         \u_DataPath/u_ifidreg/N47 , \u_DataPath/u_ifidreg/N46 ,
         \u_DataPath/u_ifidreg/N45 , \u_DataPath/u_ifidreg/N44 ,
         \u_DataPath/u_ifidreg/N43 , \u_DataPath/u_ifidreg/N42 ,
         \u_DataPath/u_ifidreg/N41 , \u_DataPath/u_ifidreg/N40 ,
         \u_DataPath/u_ifidreg/N39 , \u_DataPath/u_ifidreg/N38 ,
         \u_DataPath/u_ifidreg/N37 , \u_DataPath/u_ifidreg/N36 ,
         \u_DataPath/u_ifidreg/N35 , \u_DataPath/u_ifidreg/N34 ,
         \u_DataPath/u_ifidreg/N33 , \u_DataPath/u_ifidreg/N32 ,
         \u_DataPath/u_ifidreg/N31 , \u_DataPath/u_ifidreg/N30 ,
         \u_DataPath/u_ifidreg/N29 , \u_DataPath/u_ifidreg/N28 ,
         \u_DataPath/u_ifidreg/N27 , \u_DataPath/u_ifidreg/N26 ,
         \u_DataPath/u_ifidreg/N25 , \u_DataPath/u_ifidreg/N24 ,
         \u_DataPath/u_ifidreg/N23 , \u_DataPath/u_ifidreg/N22 ,
         \u_DataPath/u_ifidreg/N21 , \u_DataPath/u_ifidreg/N20 ,
         \u_DataPath/u_ifidreg/N19 , \u_DataPath/u_ifidreg/N18 ,
         \u_DataPath/u_ifidreg/N17 , \u_DataPath/u_ifidreg/N16 ,
         \u_DataPath/u_ifidreg/N15 , \u_DataPath/u_ifidreg/N14 ,
         \u_DataPath/u_ifidreg/N13 , \u_DataPath/u_ifidreg/N12 ,
         \u_DataPath/u_ifidreg/N11 , \u_DataPath/u_ifidreg/N10 ,
         \u_DataPath/u_ifidreg/N9 , \u_DataPath/u_ifidreg/N8 ,
         \u_DataPath/u_ifidreg/N7 , \u_DataPath/u_ifidreg/N6 ,
         \u_DataPath/u_ifidreg/N5 , \u_DataPath/u_ifidreg/N4 ,
         \u_DataPath/u_decode_unit/reg_file0/N154 ,
         \u_DataPath/u_decode_unit/reg_file0/N153 ,
         \u_DataPath/u_decode_unit/reg_file0/N152 ,
         \u_DataPath/u_decode_unit/reg_file0/N151 ,
         \u_DataPath/u_decode_unit/reg_file0/N150 ,
         \u_DataPath/u_decode_unit/reg_file0/N149 ,
         \u_DataPath/u_decode_unit/reg_file0/N148 ,
         \u_DataPath/u_decode_unit/reg_file0/N147 ,
         \u_DataPath/u_decode_unit/reg_file0/N146 ,
         \u_DataPath/u_decode_unit/reg_file0/N145 ,
         \u_DataPath/u_decode_unit/reg_file0/N144 ,
         \u_DataPath/u_decode_unit/reg_file0/N143 ,
         \u_DataPath/u_decode_unit/reg_file0/N142 ,
         \u_DataPath/u_decode_unit/reg_file0/N141 ,
         \u_DataPath/u_decode_unit/reg_file0/N140 ,
         \u_DataPath/u_decode_unit/reg_file0/N139 ,
         \u_DataPath/u_decode_unit/reg_file0/N138 ,
         \u_DataPath/u_decode_unit/reg_file0/N137 ,
         \u_DataPath/u_decode_unit/reg_file0/N136 ,
         \u_DataPath/u_decode_unit/reg_file0/N135 ,
         \u_DataPath/u_decode_unit/reg_file0/N134 ,
         \u_DataPath/u_decode_unit/reg_file0/N133 ,
         \u_DataPath/u_decode_unit/reg_file0/N132 ,
         \u_DataPath/u_decode_unit/reg_file0/N131 ,
         \u_DataPath/u_decode_unit/reg_file0/N130 ,
         \u_DataPath/u_decode_unit/reg_file0/N129 ,
         \u_DataPath/u_decode_unit/reg_file0/N128 ,
         \u_DataPath/u_decode_unit/reg_file0/N127 ,
         \u_DataPath/u_decode_unit/reg_file0/N126 ,
         \u_DataPath/u_decode_unit/reg_file0/N125 ,
         \u_DataPath/u_decode_unit/reg_file0/N124 ,
         \u_DataPath/u_decode_unit/reg_file0/N123 ,
         \u_DataPath/u_decode_unit/reg_file0/N122 ,
         \u_DataPath/u_decode_unit/reg_file0/N121 ,
         \u_DataPath/u_decode_unit/reg_file0/N120 ,
         \u_DataPath/u_decode_unit/reg_file0/N119 ,
         \u_DataPath/u_decode_unit/reg_file0/N118 ,
         \u_DataPath/u_decode_unit/reg_file0/N117 ,
         \u_DataPath/u_decode_unit/reg_file0/N116 ,
         \u_DataPath/u_decode_unit/reg_file0/N115 ,
         \u_DataPath/u_decode_unit/reg_file0/N114 ,
         \u_DataPath/u_decode_unit/reg_file0/N113 ,
         \u_DataPath/u_decode_unit/reg_file0/N112 ,
         \u_DataPath/u_decode_unit/reg_file0/N111 ,
         \u_DataPath/u_decode_unit/reg_file0/N110 ,
         \u_DataPath/u_decode_unit/reg_file0/N109 ,
         \u_DataPath/u_decode_unit/reg_file0/N108 ,
         \u_DataPath/u_decode_unit/reg_file0/N107 ,
         \u_DataPath/u_decode_unit/reg_file0/N106 ,
         \u_DataPath/u_decode_unit/reg_file0/N105 ,
         \u_DataPath/u_decode_unit/reg_file0/N104 ,
         \u_DataPath/u_decode_unit/reg_file0/N103 ,
         \u_DataPath/u_decode_unit/reg_file0/N102 ,
         \u_DataPath/u_decode_unit/reg_file0/N101 ,
         \u_DataPath/u_decode_unit/reg_file0/N100 ,
         \u_DataPath/u_decode_unit/reg_file0/N99 ,
         \u_DataPath/u_decode_unit/reg_file0/N98 ,
         \u_DataPath/u_decode_unit/reg_file0/N97 ,
         \u_DataPath/u_decode_unit/reg_file0/N96 ,
         \u_DataPath/u_decode_unit/reg_file0/N95 ,
         \u_DataPath/u_decode_unit/reg_file0/N94 ,
         \u_DataPath/u_decode_unit/reg_file0/N93 ,
         \u_DataPath/u_decode_unit/reg_file0/N92 ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][0] ,
         \u_DataPath/u_idexreg/N184 , \u_DataPath/u_idexreg/N56 ,
         \u_DataPath/u_idexreg/N44 , \u_DataPath/u_idexreg/N42 ,
         \u_DataPath/u_idexreg/N40 , \u_DataPath/u_idexreg/N39 ,
         \u_DataPath/u_idexreg/N38 , \u_DataPath/u_idexreg/N37 ,
         \u_DataPath/u_idexreg/N36 , \u_DataPath/u_idexreg/N35 ,
         \u_DataPath/u_idexreg/N34 , \u_DataPath/u_idexreg/N33 ,
         \u_DataPath/u_idexreg/N32 , \u_DataPath/u_idexreg/N31 ,
         \u_DataPath/u_idexreg/N30 , \u_DataPath/u_idexreg/N29 ,
         \u_DataPath/u_idexreg/N28 , \u_DataPath/u_idexreg/N27 ,
         \u_DataPath/u_idexreg/N26 , \u_DataPath/u_idexreg/N25 ,
         \u_DataPath/u_idexreg/N21 , \u_DataPath/u_idexreg/N20 ,
         \u_DataPath/u_idexreg/N19 , \u_DataPath/u_idexreg/N16 ,
         \u_DataPath/u_idexreg/N15 , \u_DataPath/u_idexreg/N13 ,
         \u_DataPath/u_idexreg/N11 , \u_DataPath/u_idexreg/N10 ,
         \u_DataPath/u_idexreg/N8 , \u_DataPath/u_execute/ovf_i ,
         \u_DataPath/u_execute/EXALU/N811 , \u_DataPath/u_execute/EXALU/N810 ,
         \u_DataPath/u_exmemreg/N12 , n68, n69, n70, n73, n74, n99, n100, n101,
         n102, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n137, n178, n179, n180, n189, n190, n191, n192, n193, n195,
         n196, n197, n198, n200, n201, n209, n213, n214, n215, n216, n217,
         n218, n224, n225, n226, n227, n228, n229, n230, n236, n237, n239,
         n240, n241, n242, n243, n244, n245, n246, n251, n253, n254, n255,
         n257, n258, n270, n272, n273, n274, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n288, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n323, n324, n325, n326, n327, n328, n329, n330, n335, n336,
         n337, n338, n347, n348, n1017, n1019, n1020, n1027, n1029, n1033,
         n1036, n1040, n1041, n1043, n1046, n1048, n1054, n1056, n1058, n1059,
         n1065, n1066, n1067, n1101, n1103, n1106, n1113, n1150, n1151, n1152,
         n1173, n1174, n1175, n1196, n1197, n1198, n1219, n1220, n1221, n1242,
         n1243, n1244, n1265, n1266, n1267, n1288, n1289, n1290, n1311, n1312,
         n1313, n1334, n1335, n1336, n1357, n1358, n1359, n1380, n1381, n1382,
         n1403, n1404, n1405, n1426, n1427, n1428, n1449, n1450, n1451, n1472,
         n1473, n1474, n1495, n1496, n1497, n1518, n1519, n1520, n1541, n1542,
         n1543, n1564, n1565, n1566, n1587, n1588, n1589, n1610, n1611, n1612,
         n1633, n1634, n1635, n1656, n1657, n1658, n1679, n1680, n1681, n1702,
         n1703, n1704, n1725, n1726, n1727, n1748, n1749, n1750, n1771, n1772,
         n1773, n1794, n1795, n1796, n1817, n1818, n1819, n1840, n1841, n1842,
         n1895, n1896, n1897, n1898, n1907, n1912, n1913, n1928, n1949, n1950,
         n1951, n1952, n1973, n1974, n1975, n1976, n1997, n1998, n1999, n2000,
         n2021, n2022, n2023, n2024, n2045, n2046, n2047, n2048, n2069, n2070,
         n2071, n2072, n2093, n2094, n2095, n2096, n2117, n2118, n2119, n2120,
         n2141, n2142, n2143, n2144, n2165, n2166, n2167, n2168, n2189, n2190,
         n2191, n2192, n2213, n2214, n2215, n2216, n2237, n2238, n2239, n2240,
         n2261, n2262, n2263, n2264, n2285, n2286, n2287, n2288, n2309, n2310,
         n2311, n2312, n2333, n2334, n2335, n2336, n2357, n2358, n2359, n2360,
         n2381, n2382, n2383, n2384, n2405, n2406, n2407, n2408, n2429, n2430,
         n2431, n2432, n2453, n2454, n2455, n2456, n2477, n2478, n2479, n2480,
         n2501, n2502, n2503, n2504, n2525, n2526, n2527, n2528, n2549, n2550,
         n2551, n2552, n2573, n2574, n2575, n2576, n2597, n2598, n2599, n2600,
         n2621, n2622, n2623, n2624, n2645, n2646, n2647, n2648, n2669, n2670,
         n2671, n2672, n2725, n2726, n2727, n2728, n2729, n2731, n2733, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3542, n3543, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3645, n3646, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3748, n3749,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3851,
         n3852, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3954, n3955, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4057, n4058, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4160, n4161, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4374, n4376, n4393, n4395, n4397, n4399, n4401,
         n4403, n4405, n4407, n4409, n4411, n4413, n4414, n4477, n4543, n4610,
         n4736, n4737, n4738, n4739, n4740, n4741, n4804, n4868, n4935, n5001,
         n5003, n5004, n5067, n5116, n5118, n5120, n5122, n5124, n5126, n5128,
         n5130, n5132, n5133, n5134, n5135, n5136, n5175, n5233, n5234, n5308,
         n5367, n5369, n5371, n5373, n5374, n5375, n5376, n5377, n5507, n5571,
         n5703, n5769, n5835, n5901, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5950, n5953, n5956, n5958, n5959, n5962,
         n5965, n5968, n5971, n5974, n5977, n5980, n5983, n5986, n5989, n5992,
         n5995, n5998, n6001, n6004, n6007, n6009, n6011, n6012, n6013, n6014,
         n6041, n6099, n6100, n6101, n6102, n6103, n6131, n6133, n6135, n6137,
         n6139, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6189, n6217, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6305, n6307, n6309, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6369, n6371, n6373, n6375, n6377, n6379, n6382, n6384, n6386,
         n6388, n6390, n6393, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6446, n6449, n6452, n6455, n6458, n6461, n6464, n6467, n6470,
         n6473, n6476, n6479, n6482, n6485, n6488, n6491, n6496, n6498, n6500,
         n6502, n6504, n6505, n6506, n6507, n6543, n6545, n6547, n6549, n6551,
         n6553, n6555, n6557, n6559, n6561, n6563, n6565, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6618, n6620, n6622,
         n6624, n6626, n6628, n6630, n6632, n6634, n6637, n6639, n6641, n6643,
         n6645, n6647, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6708, n6710, n6712,
         n6714, n6716, n6718, n6720, n6722, n6724, n6726, n6728, n6730, n6732,
         n6734, n6736, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6787, n6788, n6789, n6791,
         n6794, n6797, n6800, n6803, n6806, n6809, n6812, n6815, n6818, n6821,
         n6824, n6827, n6830, n6833, n6836, n6839, n6842, n6845, n6847, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6898, n6901, n6904, n6907, n6910, n6913, n6916,
         n6919, n6922, n6925, n6928, n6931, n6934, n6937, n6940, n6943, n6946,
         n6949, n6952, n6954, n6956, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n7008, n7011,
         n7014, n7017, n7020, n7023, n7026, n7029, n7032, n7035, n7038, n7041,
         n7044, n7047, n7050, n7053, n7056, n7059, n7061, n7063, n7065, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7132, n7134,
         n7136, n7138, n7140, n7142, n7144, n7146, n7148, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7201, n7203, n7205,
         n7207, n7209, n7211, n7213, n7215, n7217, n7219, n7221, n7223, n7225,
         n7227, n7229, n7231, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7302, n7304, n7306, n7308, n7310, n7312, n7314, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7365, n7368, n7371, n7374, n7377, n7380, n7383,
         n7386, n7389, n7392, n7395, n7398, n7401, n7404, n7407, n7410, n7413,
         n7416, n7418, n7420, n7422, n7424, n7425, n7426, n7427, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7499, n7502,
         n7505, n7508, n7511, n7514, n7517, n7519, n7522, n7525, n7528, n7531,
         n7534, n7537, n7540, n7543, n7546, n7549, n7551, n7553, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7606, n7608,
         n7610, n7612, n7614, n7616, n7618, n7620, n7622, n7624, n7626, n7628,
         n7630, n7632, n7634, n7636, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7689, n7692,
         n7695, n7698, n7701, n7704, n7706, n7709, n7712, n7715, n7718, n7721,
         n7724, n7727, n7730, n7733, n7736, n7739, n7742, n7744, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7796, n7798, n7800,
         n7802, n7804, n7806, n7808, n7810, n7812, n7814, n7816, n7818, n7820,
         n7822, n7824, n7826, n7828, n7830, n7832, n7833, n7834, n7835, n7836,
         n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
         n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7882, n7885,
         n7888, n7891, n7894, n7897, n7900, n7903, n7906, n7909, n7912, n7915,
         n7918, n7921, n7924, n7926, n7929, n7932, n7934, n7936, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7987, n7988, n7989, n7991, n7994, n7997, n8000, n8003,
         n8006, n8009, n8012, n8015, n8018, n8021, n8024, n8027, n8030, n8033,
         n8036, n8039, n8041, n8043, n8045, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8093,
         n8094, n8095, n8096, n8097, n8098, n8100, n8103, n8106, n8109, n8112,
         n8115, n8118, n8121, n8124, n8127, n8130, n8133, n8136, n8139, n8142,
         n8145, n8147, n8149, n8151, n8153, n8155, n8156, n8157, n8158, n8198,
         n8200, n8202, n8204, n8206, n8208, n8210, n8212, n8214, n8216, n8218,
         n8219, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230,
         n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240,
         n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250,
         n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260,
         n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270,
         n8272, n8274, n8276, n8278, n8280, n8282, n8284, n8286, n8288, n8290,
         n8292, n8294, n8296, n8298, n8300, n8302, n8304, n8305, n8306, n8307,
         n8308, n8311, n8313, n8315, n8316, n8318, n8320, n8322, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8366, n8368,
         n8370, n8372, n8374, n8376, n8378, n8380, n8382, n8384, n8386, n8388,
         n8390, n8392, n8394, n8396, n8398, n8399, n8400, n8401, n8402, n8403,
         n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
         n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8439, n8440,
         n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8451,
         n8454, n8457, n8460, n8463, n8466, n8469, n8472, n8475, n8478, n8481,
         n8484, n8487, n8490, n8493, n8496, n8499, n8501, n8503, n8505, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8558, n8561,
         n8564, n8567, n8570, n8573, n8576, n8579, n8582, n8585, n8588, n8591,
         n8594, n8597, n8600, n8603, n8606, n8609, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8641, n8642, n8643, n8644, n8645, n8646,
         n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656,
         n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8665, n8668, n8671,
         n8674, n8677, n8680, n8683, n8686, n8689, n8692, n8695, n8698, n8701,
         n8704, n8707, n8710, n8713, n8715, n8717, n8719, n8721, n8723, n8724,
         n8725, n8726, n8756, n8758, n8760, n8762, n8764, n8766, n8768, n8770,
         n8772, n8774, n8776, n8778, n8780, n8782, n8784, n8786, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8840,
         n8842, n8844, n8846, n8848, n8850, n8852, n8854, n8855, n8858, n8859,
         n8860, n8862, n8864, n8866, n8868, n8870, n8872, n8874, n8875, n8876,
         n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886,
         n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896,
         n8897, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8926, n8928, n8931, n8934, n8936, n8939, n8942, n8945, n8948, n8951,
         n8954, n8957, n8960, n8963, n8966, n8969, n8972, n8975, n8978, n8980,
         n8982, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9014, n9016, n9017, n9019, n9020, n9022, n9024, n9026, n9028, n9030,
         n9032, n9034, n9036, n9038, n9040, n9042, n9044, n9046, n9048, n9050,
         n9051, n9052, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9122, n9124, n9126, n9128, n9130, n9132, n9134, n9136, n9138,
         n9140, n9142, n9144, n9146, n9148, n9150, n9152, n9154, n9156, n9158,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9202, n9203, n9204, n9205, n9206, n9208, n9210,
         n9212, n9214, n9216, n9218, n9220, n9222, n9224, n9226, n9228, n9230,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9252, n9254,
         n9256, n9258, n9260, n9262, n9264, n9266, n9270, n9272, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9322, n9323, n9325, n9326, n9328,
         n9329, n9331, n9332, n9334, n9335, n9337, n9338, n9340, n9341, n9343,
         n9344, n9346, n9347, n9349, n9350, n9352, n9353, n9355, n9356, n9358,
         n9359, n9361, n9362, n9364, n9365, n9367, n9368, n9370, n9371, n9373,
         n9374, n9375, n9377, n9380, n9381, n9382, n9383, n9384, n9385, n9386,
         n9387, n9388, n9389, n9417, n9420, n9423, n9426, n9429, n9432, n9435,
         n9438, n9441, n9444, n9447, n9450, n9452, n9455, n9458, n9461, n9464,
         n9466, n9468, n9470, n9472, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9524,
         n9526, n9528, n9532, n9533, n9535, n9538, n9539, n9540, n9541, n9543,
         n9544, n9545, n9548, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10153, n10154, n10155, n10156, n10158, n10159,
         n10160, n10162, n10163, n10164, n10166, n10167, n10168, n10170,
         n10171, n10172, n10174, n10175, n10176, n10178, n10179, n10180,
         n10182, n10183, n10184, n10186, n10187, n10188, n10190, n10191,
         n10192, n10194, n10195, n10196, n10198, n10199, n10200, n10202,
         n10203, n10204, n10206, n10207, n10208, n10210, n10211, n10212,
         n10214, n10215, n10216, n10218, n10219, n10220, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10373, n10376, n10379, n10382,
         n10385, n10387, n10390, n10393, n10396, n10400, n10404, n10408,
         n10412, n10416, n10420, n10424, n10428, n10432, n10437, n10438,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10456, n10457, n10459, n10460,
         n10462, n10463, n10465, n10466, n10468, n10469, n10471, n10472,
         n10474, n10476, n10478, n10480, n10481, n10482, n10483, n10485,
         n10486, n10488, n10490, n10492, n10494, n10496, n10498, n10500,
         n10502, n10504, n10506, n10508, n10510, n10512, n10514, n10516,
         n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
         n10526, n10551, n10553, n10554, n10555, n10556, n10557, n10558,
         n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566,
         n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574,
         n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582,
         n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590,
         n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598,
         n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606,
         n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614,
         n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622,
         n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630,
         n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638,
         n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646,
         n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654,
         n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662,
         n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670,
         n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678,
         n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686,
         n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694,
         n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702,
         n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710,
         n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718,
         n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726,
         n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734,
         n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742,
         n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750,
         n10751, n10753, n10754, n10755, n10756, n10757, n10759, n10760,
         n10761, n10762, n10763, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10773, n10774, n10775, n10776, n10778, n10779,
         n10780, n10781, n10782, n10783, n10784, n10786, n10787, n10788,
         n10789, n10790, n10791, n10793, n10794, n10795, n10796, n10797,
         n10798, n10800, n10801, n10802, n10803, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10813, n10814, n10815, n10816,
         n10817, n10818, n10820, n10821, n10822, n10823, n10824, n10825,
         n10827, n10828, n10829, n10830, n10832, n10833, n10834, n10835,
         n10836, n10837, n10838, n10840, n10841, n10842, n10843, n10844,
         n10845, n10847, n10848, n10849, n10850, n10852, n10853, n10854,
         n10855, n10856, n10857, n10858, n10860, n10861, n10862, n10863,
         n10864, n10865, n10867, n10868, n10869, n10870, n10871, n10872,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n11417, n11418,
         n11436, n11437, n11438, n11439, n11440, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11475, n11476, n11477, n11478,
         n11479, n11480, n11481, n11482, n11483, n11484, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11534, n11535, n11536, n11537, n11538, n11539, n11540,
         n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548,
         n11549, n11550, n11553, n11554, n11555, n11556, n11557, n11558,
         n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566,
         n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574,
         n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582,
         n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590,
         n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598,
         n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606,
         n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614,
         n11615, n11616, n11618, n11619, n11620, n11622, n11624, n11625,
         n11626, n11628, n11629, n11630, n11632, n11633, n11634, n11636,
         n11637, n11638, n11640, n11641, n11642, n11643, n11644, n11645,
         n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653,
         n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661,
         n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669,
         n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677,
         n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685,
         n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693,
         n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701,
         n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709,
         n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717,
         n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725,
         n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733,
         n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741,
         n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749,
         n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757,
         n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765,
         n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773,
         n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781,
         n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789,
         n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797,
         n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805,
         n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813,
         n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821,
         n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829,
         n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837,
         n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845,
         n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853,
         n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861,
         n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869,
         n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877,
         n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885,
         n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893,
         n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901,
         n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909,
         n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917,
         n11918, n11919, n11920, n11921, n11923, n11925, n11927, n11929,
         n11931, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
         n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
         n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
         n11964, n11966, n11968, n11970, n11972, n11974, n11976, n11978,
         n11980, n11982, n11984, n11986, n11987, n11988, n11989, n11990,
         n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998,
         n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006,
         n12007, n12008, n12009, n12010, n12011, n12013, n12015, n12017,
         n12019, n12021, n12023, n12025, n12027, n12029, n12031, n12033,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12056, n12058, n12060, n12062,
         n12064, n12066, n12068, n12070, n12072, n12074, n12076, n12078,
         n12080, n12082, n12084, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12103, n12105, n12107, n12109, n12111,
         n12113, n12115, n12117, n12119, n12121, n12123, n12125, n12127,
         n12129, n12131, n12133, n12135, n12137, n12138, n12139, n12140,
         n12141, n12142, n12143, n12144, n12146, n12148, n12150, n12152,
         n12154, n12156, n12158, n12160, n12162, n12164, n12166, n12168,
         n12170, n12172, n12174, n12176, n12178, n12180, n12182, n12184,
         n12186, n12187, n12188, n12189, n12190, n12191, n12193, n12195,
         n12197, n12199, n12201, n12203, n12205, n12207, n12209, n12211,
         n12213, n12215, n12217, n12219, n12221, n12223, n12225, n12227,
         n12229, n12231, n12232, n12233, n12234, n12236, n12238, n12240,
         n12242, n12244, n12246, n12248, n12250, n12252, n12254, n12256,
         n12258, n12260, n12262, n12264, n12266, n12268, n12270, n12272,
         n12274, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
         n12483, n12484, n12485, n12486, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
         n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
         n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
         n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
         n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731,
         n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
         n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747,
         n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
         n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
         n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771,
         n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
         n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
         n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
         n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803,
         n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
         n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819,
         n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
         n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
         n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843,
         n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
         n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
         n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
         n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
         n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931,
         n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939,
         n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947,
         n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955,
         n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963,
         n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971,
         n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979,
         n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987,
         n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995,
         n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003,
         n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011,
         n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019,
         n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027,
         n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035,
         n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
         n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051,
         n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
         n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067,
         n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075,
         n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083,
         n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091,
         n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099,
         n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107,
         n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
         n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123,
         n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131,
         n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139,
         n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147,
         n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155,
         n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163,
         n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171,
         n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179,
         n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187,
         n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195,
         n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203,
         n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211,
         n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219,
         n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227,
         n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235,
         n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243,
         n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
         n13252, n13253, n13254, n13255, n13256, n13257, n13259, n13260,
         n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268,
         n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276,
         n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284,
         n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292,
         n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300,
         n13302, n13304, n13306, n13308, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13349, n13351, n13353, n13355, n13357, n13359,
         n13361, n13363, n13365, n13367, n13369, n13371, n13373, n13375,
         n13377, n13379, n13381, n13383, n13385, n13387, n13388, n13389,
         n13390, n13392, n13394, n13396, n13398, n13400, n13402, n13404,
         n13406, n13408, n13410, n13412, n13414, n13416, n13418, n13420,
         n13422, n13424, n13426, n13428, n13430, n13432, n13433, n13434,
         n13435, n13436, n13437, n13439, n13441, n13443, n13445, n13447,
         n13449, n13451, n13453, n13455, n13457, n13459, n13461, n13463,
         n13465, n13467, n13469, n13471, n13473, n13475, n13477, n13478,
         n13479, n13480, n13482, n13484, n13486, n13488, n13490, n13492,
         n13494, n13496, n13498, n13500, n13502, n13504, n13506, n13508,
         n13510, n13512, n13514, n13516, n13518, n13520, n13522, n13523,
         n13524, n13525, n13526, n13527, n13528, n13530, n13531, n13532,
         n13533, n13536, n13537, n13538, n13539, n13540, n13541, n13542,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13556,
         n13557, n13558, n13559, n13560, n13561, n13565, n13566, n13567,
         n13568, n13569, n13570, n13574, n13575, n13576, n13577, n13578,
         n13579, n13582, n13583, n13584, n13585, n13586, n13587, n13589,
         n13590, n13591, n13592, n13593, n13594, n13596, n13597, n13599,
         n13600, n13601, n13603, n13604, n13605, n13606, n13607, n13609,
         n13610, n13612, n13613, n13614, n13616, n13618, n13619, n13621,
         n13622, n13624, n13626, n13628, n13630, n13632, n13633, n13635,
         n13636, n13637, n13639, n13640, n13641, n13642, n13643, n13644,
         n13645, n13646, n13647, n13648, n13649, n13650, n13652, n13653,
         n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661,
         n13662, n13663, n13665, n13666, n13667, n13668, n13669, n13670,
         n13671, n13672, n13673, n13674, n13675, n13676, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13730, n13731,
         n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739,
         n13740, n13741, n13743, n13744, n13745, n13746, n13747, n13748,
         n13749, n13750, n13751, n13752, n13753, n13755, n13756, n13757,
         n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13766,
         n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774,
         n13775, n13776, n13777, n13779, n13780, n13781, n13782, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13830, n13831, n13832, n13833, n13834, n13835,
         n13836, n13837, n13838, n13839, n13841, n13842, n13843, n13844,
         n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852,
         n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861,
         n13862, n13863, n13864, n13865, n13867, n13868, n13869, n13870,
         n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878,
         n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886,
         n13887, n13888, n13889, n13890, n13892, n13893, \nibble[0]_snps_wire ,
         n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902,
         n13903, n13904, n13905, \Data_in[15]_snps_wire , n13907,
         \Data_in[14]_snps_wire , n13909, \Data_in[9]_snps_wire , n13911,
         \Data_in[11]_snps_wire , n13913, \Data_in[10]_snps_wire , n13915,
         \Data_in[8]_snps_wire , n13917, \Data_in[13]_snps_wire , n13919,
         \Data_in[12]_snps_wire , n13921, \Data_in[30]_snps_wire , n13923,
         \Data_in[29]_snps_wire , n13925, \Address_toRAM[10]_snps_wire ,
         n13927, \Address_toRAM[7]_snps_wire , n13929,
         \Address_toRAM[11]_snps_wire , n13931, \Address_toRAM[9]_snps_wire ,
         n13933, \Address_toRAM[4]_snps_wire , n13935,
         \Address_toRAM[6]_snps_wire , n13937, \Address_toRAM[2]_snps_wire ,
         n13939, \Address_toRAM[5]_snps_wire , n13941,
         \Address_toRAM[3]_snps_wire , n13943, n13944, n13945, addr_to_iram_29,
         addr_to_iram_28, addr_to_iram_27, addr_to_iram_26, addr_to_iram_25,
         addr_to_iram_24, addr_to_iram_23, addr_to_iram_22, addr_to_iram_21,
         addr_to_iram_20, addr_to_iram_19, addr_to_iram_18, addr_to_iram_17,
         addr_to_iram_16, addr_to_iram_15, addr_to_iram_14, addr_to_iram_13,
         addr_to_iram_12, addr_to_iram_11, addr_to_iram_10, addr_to_iram_9,
         addr_to_iram_8, addr_to_iram_7, addr_to_iram_6, addr_to_iram_5,
         addr_to_iram_4, addr_to_iram_3, addr_to_iram_2, addr_to_iram_1,
         addr_to_iram_0, n13947, n13949, n13951, n13953, n13955, n13957,
         n13959, n13961, n13963, n13965, n13967, n13969, n13971, n13973,
         n13975, n13977, n13979, n13981, n13983, n13985, n13987, n13989,
         n13991, n13993, n13995, n13997, n13999, n14001, n14002, n14004,
         n14005, n14006, n14008, \Data_in[7]_snps_wire , n14010,
         read_op_snps_wire, n14012, \Data_in[22]_snps_wire , n14014,
         \Data_in[21]_snps_wire , n14016, \Data_in[20]_snps_wire , n14018,
         \Data_in[19]_snps_wire , n14020, \Data_in[18]_snps_wire , n14022,
         \Data_in[17]_snps_wire , n14024, \Data_in[16]_snps_wire , n14026,
         n14027, n14029, n14030, n14031, n14032, n14033, n14034, n14035,
         n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043,
         n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051,
         n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059,
         n14060, n14064, n14065, write_byte_snps_wire, n14067, n14068, n14069,
         n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
         n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085,
         n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093,
         n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101,
         n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109,
         n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117,
         n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
         n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133,
         n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141,
         n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
         n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157,
         n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
         n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
         n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181,
         n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189,
         n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197,
         n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205,
         n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213,
         n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221,
         n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14230,
         n14231, n14232, n14233, n14234, n14235, n14236, n14238, n14239,
         n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
         n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
         n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271,
         n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
         n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
         n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
         n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
         n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
         n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
         n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399,
         n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14510, n14511, n14513, n14514, n14515,
         n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523,
         n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531,
         n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539,
         n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547,
         n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555,
         n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563,
         n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571,
         n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
         n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
         n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595,
         n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603,
         n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611,
         n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619,
         n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627,
         n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635,
         n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643,
         n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
         n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
         n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667,
         n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
         n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683,
         n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691,
         n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699,
         n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
         n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715,
         n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
         n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
         n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739,
         n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
         n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
         n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14842, n14843, n14844,
         n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852,
         n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860,
         n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868,
         n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876,
         n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884,
         n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892,
         n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900,
         n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908,
         n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916,
         n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924,
         n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932,
         n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940,
         n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948,
         n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956,
         n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964,
         n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972,
         n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980,
         n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988,
         n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996,
         n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004,
         n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012,
         n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020,
         n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028,
         n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036,
         n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044,
         n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052,
         n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060,
         n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068,
         n15069, n15070, n15071, n15073, n15074, n15075, n15076, n15077,
         n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085,
         n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093,
         n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101,
         n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109,
         n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117,
         n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125,
         n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133,
         n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141,
         n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149,
         n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157,
         n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165,
         n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173,
         n15174, n15175, n15177, n15178, n15179, n15180, n15181, n15182,
         n15183, n15185, n15186, n15187, n15188, n15189, n15190, n15191,
         n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199,
         n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207,
         n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215,
         n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223,
         n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231,
         n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239,
         n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247,
         n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255,
         n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263,
         n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271,
         n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279,
         n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287,
         n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295,
         n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303,
         n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311,
         n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319,
         n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327,
         n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335,
         n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343,
         n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351,
         n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359,
         n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367,
         n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375,
         n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383,
         n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391,
         n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399,
         n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407,
         n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415,
         n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423,
         n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431,
         n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439,
         n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447,
         n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455,
         n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463,
         n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471,
         n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479,
         n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487,
         n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495,
         n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503,
         n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511,
         n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15520,
         n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,
         n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,
         n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
         n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552,
         n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, \Address_toRAM[8]_snps_wire ,
         n15664, n15665, \Data_in[27]_snps_wire , \Data_in[28]_snps_wire ,
         \Data_in[31]_snps_wire , n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15717, n15718, n15719, n15720, n15721, n15722,
         n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730,
         n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738,
         n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746,
         n15747, n15748, n15749, n15750, n15751, n15753, n15754, n15755,
         n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763,
         n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771,
         n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779,
         n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787,
         n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795,
         n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803,
         n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811,
         n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819,
         n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827,
         n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835,
         n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843,
         n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851,
         n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859,
         n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867,
         n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875,
         n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883,
         n15884, n15885, n15886, n15887, n15888, n15889, n15890, n15891,
         n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899,
         n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907,
         n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915,
         n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923,
         n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931,
         n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939,
         n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947,
         n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955,
         n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963,
         n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971,
         n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979,
         n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987,
         n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995,
         n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003,
         n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011,
         n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019,
         n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027,
         n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035,
         n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043,
         n16044, n16046, n16047, n16048, n16049, n16050, n16051, n16052,
         n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16060,
         n16061, n16062, n16063, n16064, n16065, n16066, n16067, n16068,
         n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076,
         n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084,
         n16085, n16086, n16087, n16088, n16089, n16090, n16091, n16092,
         n16093, n16094, n16095, n16096, n16097, n16098, n16099, n16100,
         n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108,
         n16109, n16110, n16111, n16112, n16113, n16114, n16115, n16116,
         n16117, n16118, n16119, n16120, n16121, n16122, n16123, n16124,
         n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132,
         n16133, n16134, n16135, n16136, n16137, n16138, n16139, n16140,
         n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148,
         n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156,
         n16157, n16158, n16159, n16160, n16161, n16162, n16163, n16164,
         n16165, n16166, n16167, n16168, n16169, n16170, n16171, n16172,
         n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180,
         n16181, n16182, n16183, n16184, n16185, n16186, n16187, n16188,
         n16189, n16190, n16191, n16192, n16193, n16194, n16195, n16196,
         n16197, n16198, n16199, n16200, n16201, n16202, n16203, n16204,
         n16205, n16206, n16207, n16208, n16209, n16210, n16211, n16212,
         n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220,
         n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228,
         n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236,
         n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244,
         n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252,
         n16253, n16254, n16255, n16256, n16257, n16258, n16259, n16260,
         n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268,
         n16269, n16270, n16271, n16272, n16273, n16274, n16275, n16276,
         n16277, n16278, n16279, n16280, n16281, n16282, n16283, n16284,
         n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292,
         n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300,
         n16301, n16302, n16304, n16305, n16306, n16307, n16309, n16310,
         n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318,
         n16319, n16320, n16321, n16322, n16323, n16325, n16326, n16327,
         n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335,
         n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343,
         n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351,
         n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359,
         n16360, n16361, n16362, n16363, n16364, n16365, n16367, n16368,
         n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376,
         n16377, n16379, n16380, n16381, n16383, n16384, n16385, n16386,
         n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394,
         n16395, n16396, n16397, n16399, n16400, n16401, n16402, n16403,
         n16404, n16405, n16406, n16408, n16409, n16410, n16411, n16412,
         n16413, n16414, n16415, n16417, n16418, n16419, n16420, n16421,
         n16424, n16425, n16426, n16427, n16429, n16432, n16433, n16436,
         n16437, n16439, n16442, n16443, n16444, n16445, n16446, n16447,
         n16450, n16452, n16453, n16455, n16456, n16457, n16458, n16459,
         n16460, n16461, n16464, n16466, n16468, n16469, n16470, n16471,
         n16473, n16474, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690,
         n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698,
         n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706,
         n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714,
         n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722,
         n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730,
         n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738,
         n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746,
         n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754,
         n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762,
         n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770,
         n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778,
         n16779, n16780, n16781, n16782, n16783, n16784, n16785, n16786,
         n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794,
         n16795, n16796, n16797, n16798, n16799, n16800, n16801, n16802,
         n16803, n16804, n16805, n16806, n16807, n16808, n16809, n16810,
         n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818,
         n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826,
         n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834,
         n16835, n16836, n16837, n16838, n16839, n16841, n16842, n16843,
         n16844, n16845, n16846, n16847, n16848, n16849, n16850, n16851,
         n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859,
         n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867,
         n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875,
         n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883,
         n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16891,
         n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899,
         n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907,
         n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915,
         n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923,
         n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931,
         n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939,
         n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947,
         n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955,
         n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963,
         n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971,
         n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979,
         n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987,
         n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995,
         n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003,
         n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011,
         n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019,
         n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027,
         n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035,
         n17036, n17037, n17038, n17039, n17040, n17041, n17043, n17044,
         n17045, n17046, n17047, n17048, n17049, n17050, n17051, n17052,
         n17053, n17054, n17055, n17056, n17057, n17058, n17059, n17060,
         n17061, n17062, n17063, n17064, n17065, n17066, n17067, n17068,
         n17069, n17070, n17071, n17072, n17073, n17074, n17075, n17076,
         n17077, n17078, n17079, n17080, n17081, n17082, n17083, n17084,
         n17085, n17086, n17087, n17088, n17089, n17090, n17091, n17092,
         n17093, n17094, n17095, n17096, n17097, n17098, n17099, n17100,
         n17101, n17102, n17103, n17104, n17105, n17106, n17107, n17108,
         n17109, n17110, n17111, n17112, n17113, n17114, n17116, n17117,
         n17118, n17119, n17120, n17121, n17122, n17123, n17124, n17125,
         n17126, n17127, n17128, n17129, n17130, n17131, n17132, n17133,
         n17134, n17135, n17136, n17137, n17138, n17139, n17140, n17141,
         n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149,
         n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17157,
         n17158, n17159, n17160, n17161, n17162, n17164, n17165, n17166,
         n17167, n17168, n17169, n17170, n17171, n17172, n17173, n17174,
         n17175, n17176, n17177, n17178, n17179, n17180, n17181, n17182,
         n17183, n17184, n17185, n17186, n17187, n17188, n17189, n17190,
         n17191, n17192, n17193, n17194, n17195, n17196, n17197, n17198,
         n17199, n17200, n17201, n17202, n17203, n17204, n17205, n17206,
         n17207, n17208, n17209, n17210, n17211, n17213, n17214, n17245,
         n17246, n17247, n17248, n17249, n17250, n17251, n17252, n17253,
         n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261,
         n17262, n17263, n17264, n17265, n17266, n17267, n17268, n17269,
         n17270, n17271, n17272, n17273, n17274, n17275, n17276, n17277,
         n17278, n17279, n17280, n17281, n17282, n17283, n17284, n17285,
         n17286, n17287, n17288, n17289, n17290, n17291, n17292, n17293,
         n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301,
         n17302, n17303, n17304, n17305, n17306, n17307, n17308, n17309,
         n17310, n17311, n17312, n17313, n17314, n17315, n17316, n17317,
         n17318, n17319, n17320, n17321, n17322, n17323, n17324, n17325,
         n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333,
         n17334, n17335, n17336, n17337, n17338, n17339, n17340, n17341,
         n17342, n17343, n17344, n17345, n17346, n17347, n17348, n17349,
         n17350, n17351, n17352, n17353, n17354, n17355, n17356, n17357,
         n17358, n17359, n17360, n17361, n17362, n17363, n17364, n17365,
         n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373,
         n17374, n17375, n17376, n17377, n17378, n17379, n17380, n17381,
         n17382, n17383, n17384, n17385, n17386, n17387, n17388, n17389,
         n17390, n17391, n17392, n17393, n17394, n17395, n17396, n17397,
         n17398, n17399, n17400, n17401, n17402, n17403, n17404, n17405,
         n17406, n17407, n17408, n17409, n17410, n17411, n17412, n17413,
         n17414, n17415, n17416, n17417, n17418, n17419, n17420, n17421,
         n17422, n17423, n17424, n17425, n17426, n17427, n17428, n17429,
         n17430, n17431, n17432, n17433, n17434, n17435, n17436, n17437,
         n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445,
         n17446, n17447, n17448, n17449, n17450, n17451, n17452, n17453,
         n17454, n17455, n17456, n17457, n17458, n17459, n17460, n17461,
         n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469,
         n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477,
         n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485,
         n17486, n17487, n17488, n17489, n17490, n17491, n17492, n17493,
         n17494, n17495, n17496, n17497, n17498, n17499, n17500, n17501,
         n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509,
         n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517,
         n17518, n17519, n17520, n17521, n17522, n17523, n17524, n17525,
         n17526, n17527, n17528, n17529, n17530, n17531, n17532, n17533,
         n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541,
         n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549,
         n17550, n17551, n17552, n17553, n17554, n17555, n17556, n17557,
         n17558, n17559, n17560, n17561, n17562, n17563, n17564, n17565,
         n17566, n17567, n17568, n17569, n17570, n17571, n17572, n17573,
         n17574, n17575, n17576, n17577, n17578, n17579, n17580, n17581,
         n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589,
         n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597,
         n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605,
         n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613,
         n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621,
         n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629,
         n17630, n17631, n17632, n17633, n17634, n17635, n17636, n17637,
         n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645,
         n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653,
         n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661,
         n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669,
         n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677,
         n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685,
         n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693,
         n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701,
         n17702, n17703, n17704, n17705, n17706, n17707, n17708, n17709,
         n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717,
         n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725,
         n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733,
         n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741,
         n17742, n17743, n17744, n17745, n17746, n17747, n17748, n17749,
         n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757,
         n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765,
         n17766, n17767, n17768, n17769, n17770, n17771, n17772, n17773,
         n17774, n17775, n17776, n17777, n17778, n17779, n17780, n17781,
         n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789,
         n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797,
         n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805,
         n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813,
         n17814, n17815, n17816, n17817, n17818, n17819, n17820, n17821,
         n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829,
         n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837,
         n17838, n17839, n17840, n17841, n17842, n17843, n17844, n17845,
         n17846, n17847, n17848, n17849, n17850, n17851, n17852, n17853,
         n17854, n17855, n17856, n17857, n17858, n17859, n17860, n17861,
         n17862, n17863, n17864, n17865, n17866, n17867, n17868, n17869,
         n17870, n17871, n17872, n17873, n17874, n17875, n17876, n17877,
         n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17885,
         n17886, n17887, n17888, n17889, n17890, n17891, n17892, n17893,
         n17894, n17895, n17896, n17897, n17898, n17899, n17900, n17901,
         n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909,
         n17910, n17911, n17912, n17913, n17914, n17915, n17916, n17917,
         n17918, n17919, n17920, n17921, n17922, n17923, n17924, n17925,
         n17926, n17927, n17928, n17929, n17930, n17931, n17932, n17933,
         n17934, n17935, n17936, n17937, n17938, n17939, n17940, n17941,
         n17942, n17943, n17944, n17945, n17946, n17947, n17948, n17949,
         n17950, n17951, n17952, n17953, n17954, n17955, n17956, n17957,
         n17958, n17959, n17960, n17961, n17962, n17963, n17964, n17965,
         n17966, n17967, n17968, n17969, n17970, n17971, n17972, n17973,
         n17974, n17975, n17976, n17977, n17978, n17979, n17980, n17981,
         n17982, n17983, n17984, n17985, n17986, n17987, n17988, n17989,
         n17990, n17991, n17992, n17993, n17994, n17995, n17996, n17997,
         n17998, n17999, n18000, n18001, n18002, n18003, n18004, n18005,
         n18006, n18007, n18008, n18009, n18010, n18011, n18012, n18013,
         n18014, n18015, n18016, n18017, n18018, n18019, n18020, n18021,
         n18022, n18023, n18024, n18025, n18026, n18027, n18028, n18029,
         n18030, n18031, n18032, n18033, n18034, n18035, n18036, n18037,
         n18038, n18039, n18040, n18041, n18042, n18043, n18044, n18045,
         n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053,
         n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061,
         n18062, n18063, n18064, n18065, n18066, n18067, n18068, n18069,
         n18070, n18071, n18072, n18073, n18074, n18075, n18076, n18077,
         n18078, n18079, n18080, n18081, n18082, n18083, n18084, n18085,
         n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093,
         n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101,
         n18102, n18103, n18104, n18105, n18106, n18107, n18108, n18109,
         n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117,
         n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125,
         n18126, n18127, n18128, n18129, n18130, n18131, n18132, n18133,
         n18134, n18135, n18136, n18137, n18138, n18139, n18140, n18141,
         n18142, n18143, n18144, n18145, n18146, n18147, n18148, n18149,
         n18150, n18151, n18152, n18153, n18154, n18155, n18156, n18157,
         n18158, n18159, n18160, n18348, n19087, n19088, n19089, n19090,
         n20341, n20342, n20433, n20916, n21117, n21638, n21749, n21994,
         n22001, n22006, n24656, n25850, n25851, n25922, n26240, n26241,
         n26257, n26258, n26577, n26759, n27019, n27066, n27100, n27442,
         n27462, n27481, n27498, n27516, n27534, n27555, n27573, n27591,
         n27609, n27626, n27639, n27652, n27665, n27787, n27790, n29426,
         n29434, n29440, n29442, n29443, n29451, n29534, n29535, n29536,
         n29538, n29540, n29542, n29543, n29547, n29548, n29549, n29551,
         n29552, n29553, n29554, n29559, n29560, n29561, n29562, n29563,
         n29564, n29565, n29566, n29567, n29568, n29569, n29570, n29571,
         n29572, n29573, n29574, n29575, n29576, n29577, n29578, n29579,
         n29580, n29581, n29582, n29583, n29584, n29585, n29586, n29587,
         n29588, n29589, n29590, n29591, n29592, n29593, n29594, n29595,
         n29596, n29597, n29598, n29599, n29600, n29602, n29603, n29604,
         n29605, n29606, n29609, n29610, n29615, n29616, n29617, n29618,
         n29619, n29620, n29622, n29623, n29624, n29635, n29643, n29644,
         n29645, n29646, n29647, n29648, n29649, n29650, n29651, n29652,
         n29653, n29654, n29655, n29656, n29657, n29658, n29659, n29660,
         n29661, n29662, n29663, n29664, n29665, n29666, n29667, n29668,
         n29669, n29670, n29671, n29672, n29673, n29674, n29675, n29676,
         n29677, n29678, n29679, n29680, n29681, n29682, n29683, n29684,
         n29685, n29686, n29687, n29688, n29689, n29690, n29691, n29692,
         n29693, n29694, n29697, n29698, n29699, n29700, n29701, n29702,
         n29703, n29704, n29705, n29706, n29707, n29708, n29709, n29710,
         n29711, n29712, n29713, n29714, n29715, n29716, n29717, n29718,
         n29719, n29720, n29721, n29722, n29723, n29724, n29725, n29726,
         n29727, n29728, n29729, n29730, n29731, n29732, n29733, n29734,
         n29735, n29736, n29737, n29738, n29739, n29740, n29741, n29742,
         n29743, n29744, n29745, n29746, n29747, n29748, n29749, n29750,
         n29751, n29752, n29753, n29754, n29755, n29756, n29757, n29758,
         n29759, n29760, n29761, n29762, n29763, n29764, n29765, n29766,
         n29767, n29768, n29769, n29770, n29771, n29772, n29773, n29774,
         n29775, n29776, n29777, n29778, n29779, n29780, n29781, n29782,
         n29783, n29784, n29785, n29786, n29787, n29788, n29789, n29790,
         n29791, n29792, n29793, n29794, n29795, n29796, n29797, n29798,
         n29799, n29800, n29801, n29802, n29803, n29804, n29805, n29806,
         n29807, n29808, n29809, n29810, n29811, n29812, n29813, n29814,
         n29815, n29816, n29817, n29818, n29819, n29820, n29821, n29822,
         n29823, n29824, n29825, n29826, n29827, n29828, n29829, n29830,
         n29831, n29832, n29833, n29834, n29835, n29836, n29837, n29838,
         n29839, n29840, n29841, n29842, n29843, n29844, n29845, n29846,
         n29847, n29848, n29849, n29850, n29851, n29852, n29853, n29854,
         n29855, n29856, n29857, n29858, n29859, n29860, n29861, n29862,
         n29863, n29864, n29865, n29866, n29867, n29868, n29869, n29870,
         n29871, n29872, n29873, n29874, n29875, n29876, n29877, n29878,
         n29879, n29880, n29881, n29882, n29883, n29884, n29885, n29886,
         n29887, n29888, n29889, n29890, n29891, n29892, n29893, n29894,
         n29895, n29896, n29897, n29898, n29899, n29900, n29901, n29902,
         n29903, n29904, n29905, n29906, n29907, n29908, n29909, n29910,
         n29911, n29912, n29913, n29914, n29915, n29916, n29917, n29918,
         n29919, n29920, n29921, n29922, n29923, n29924, n29925, n29926,
         n29927, n29928, n29929, n29930, n29931, n29932, n29933, n29934,
         n29935, n29936, n29937, n29938, n29939, n29940, n29941, n29942,
         n29943, n29944, n29945, n29946, n29947, n29948, n29949, n29950,
         n29951, n29952, n29953, n29954, n29955, n29956, n29957, n29958,
         n29959, n29960, n29961, n29962, n29963, n29964, n29965, n29966,
         n29967, n29968, n29969, n29970, n29971, n29972, n29973, n29974,
         n29975, n29976, n29977, n29978, n29979, n29980, n29981, n29982,
         n29983, n29984, n29985, n29986, n29987, n29988, n29989, n29990,
         n29991, n29992, n29993, n29994, n29995, n29996, n29997, n29998,
         n29999, n30000, n30001, n30002, n30003, n30004, n30005, n30006,
         n30007, n30008, n30009, n30010, n30011, n30012, n30013, n30014,
         n30015, n30016, n30017, n30018, n30019, n30020, n30021, n30022,
         n30023, n30024, n30025, n30026, n30027, n30028, n30029, n30030,
         n30031, n30032, n30033, n30034, n30035, n30036, n30037, n30038,
         n30039, n30040, n30041, n30042, n30043, n30044, n30045, n30046,
         n30047, n30048, n30049, n30050, n30051, n30052, n30053, n30054,
         n30055, n30056, n30057, n30058, n30059, n30060, n30061, n30062,
         n30063, n30064, n30065, n30066, n30067, n30068, n30069, n30070,
         n30071, n30072, n30073, n30074, n30075, n30076, n30077, n30078,
         n30079, n30080, n30081, n30082, n30083, n30084, n30085, n30086,
         n30087, n30088, n30089, n30090, n30091, n30092, n30093, n30094,
         n30095, n30096, n30097, n30098, n30099, n30100, n30101, n30102,
         n30103, n30104, n30105, n30106, n30107, n30108, n30109, n30110,
         n30111, n30112, n30113, n30114, n30115, n30116, n30117, n30118,
         n30119, n30120, n30121, n30122, n30123, n30124, n30125, n30126,
         n30127, n30128, n30129, n30130, n30131, n30132, n30133, n30134,
         n30135, n30136, n30137, n30138, n30139, n30140, n30141, n30142,
         n30143, n30144, n30145, n30146, n30147, n30148, n30149, n30150,
         n30151, n30152, n30153, n30154, n30155, n30156, n30157, n30158,
         n30159, n30160, n30161, n30162, n30163, n30164, n30165, n30166,
         n30167, n30168, n30169, n30170, n30171, n30172, n30173, n30174,
         n30175, n30176, n30177, n30178, n30179, n30180, n30181, n30182,
         n30183, n30184, n30185, n30186, n30187, n30188, n30189, n30190,
         n30191, n30192, n30193, n30194, n30195, n30196, n30197, n30198,
         n30199, n30200, n30201, n30202, n30203, n30204, n30205, n30206,
         n30207, n30208, n30209, n30210, n30211, n30212, n30213, n30214,
         n30215, n30216, n30217, n30218, n30219, n30220, n30221, n30222,
         n30223, n30224, n30225, n30226, n30227, n30228, n30229, n30230,
         n30231, n30232, n30233, n30234, n30235, n30236, n30237, n30238,
         n30239, n30240, n30241, n30242, n30243, n30244, n30245, n30246,
         n30247, n30248, n30249, n30250, n30251, n30252, n30253, n30254,
         n30255, n30256, n30257, n30258, n30259, n30260, n30261, n30262,
         n30263, n30264, n30265, n30266, n30267, n30268, n30269, n30270,
         n30271, n30272, n30273, n30274, n30275, n30276, n30277, n30278,
         n30279, n30280, n30281, n30282, n30283, n30284, n30285, n30286,
         n30287, n30288, n30289, n30290, n30291, n30292, n30293, n30294,
         n30295, n30296, n30297, n30298, n30299, n30300, n30301, n30302,
         n30303, n30304, n30305, n30306, n30307, n30308, n30309, n30310,
         n30311, n30312, n30313, n30314, n30315, n30316, n30317, n30318,
         n30319, n30320, n30321, n30322, n30323, n30324, n30325, n30326,
         n30327, n30328, n30329, n30330, n30331, n30332, n30333, n30334,
         n30335, n30336, n30337, n30338, n30339, n30340, n30341, n30342,
         n30343, n30344, n30345, n30346, n30347, n30348, n30349, n30350,
         n30351, n30352, n30353, n30354, n30355, n30356, n30357, n30358,
         n30359, n30360, n30361, n30362, n30363, n30364, n30365, n30366,
         n30367, n30368, n30369, n30370, n30371, n30372, n30373, n30374,
         n30375, n30376, n30377, n30378, n30379, n30380, n30381, n30382,
         n30383, n30384, n30385, n30386, n30387, n30388, n30389, n30390,
         n30391, n30392, n30393, n30394, n30395, n30396, n30397, n30398,
         n30399, n30400, n30401, n30402, n30403, n30404, n30405, n30406,
         n30407, n30408, n30409, n30410, n30411, n30412, n30413, n30414,
         n30415, n30416, n30417, n30418, n30419, n30420, n30421, n30422,
         n30423, n30424, n30425, n30426, n30427, n30428, n30429, n30430,
         n30431, n30432, n30433, n30434, n30435, n30436, n30437, n30438,
         n30439, n30440, n30441, n30442, n30443, n30444, n30445, n30446,
         n30447, n30448, n30449, n30450, n30451, n30452, n30453, n30454,
         n30455, n30456, n30457, n30458, n30459, n30460, n30461, n30462,
         n30463, n30464, n30465, n30466, n30467, n30468, n30469, n30470,
         n30471, n30472, n30473, n30474, n30475, n30476, n30477, n30478,
         n30479, n30480, n30481, n30482, n30483, n30484, n30485, n30486,
         n30487, n30488, n30489, n30490, n30491, n30492, n30493, n30494,
         n30495, n30496, n30497, n30498, n30499, n30500, n30501, n30502,
         n30503, n30504, n30505, n30506, n30507, n30508, n30509, n30510,
         n30511, n30512, n30513, n30514, n30515, n30516, n30517, n30518,
         n30519, n30520, n30521, n30522, n30523, n30524, n30525, n30526,
         n30527, n30528, n30529, n30530, n30531, n30532, n30533, n30534,
         n30535, n30536, n30537, n30538, n30539, n30540, n30541, n30542,
         n30543, n30544, n30545, n30546, n30547, n30548, n30549, n30550,
         n30551, n30552, n30553, n30554, n30555, n30556, n30557, n30558,
         n30559, n30560, n30561, n30562, n30563, n30564, n30565, n30566,
         n30567, n30568, n30569, n30570, n30571, n30572, n30573, n30574,
         n30575, n30576, n30577, n30578, n30579, n30580, n30581, n30582,
         n30583, n30584, n30585, n30586, n30587, n30588, n30589, n30590,
         n30591, n30592, n30593, n30594, n30595, n30596, n30597, n30598,
         n30599, n30600, n30601, n30602, n30603, n30604, n30605, n30606,
         n30607, n30608, n30609, n30610, n30611, n30612, n30613, n30614,
         n30615, n30616, n30617, n30618, n30619, n30620, n30621, n30622,
         n30623, n30624, n30625, n30626, n30627, n30628, n30629, n30630,
         n30631, n30632, n30633, n30634, n30635, n30636, n30637, n30638,
         n30639, n30640, n30641, n30642, n30643, n30644, n30645, n30646,
         n30647, n30648, n30649, n30650, n30651, n30652, n30653, n30654,
         n30655, n30656, n30657, n30658, n30659, n30660, n30661, n30662,
         n30663, n30664, n30665, n30666, n30667, n30668, n30669, n30670,
         n30671, n30672, n30673, n30674, n30675, n30676, n30677, n30678,
         n30679, n30680, n30681, n30682, n30683, n30684, n30685, n30686,
         n30687, n30688, n30689, n30690, n30691, n30692, n30693, n30694,
         n30695, n30696, n30697, n30698, n30699, n30700, n30701, n30702,
         n30703, n30704, n30705, n30706, n30707, n30708, n30709, n30710,
         n30711, n30712, n30713, n30714, n30715, n30716, n30717, n30718,
         n30719, n30720, n30721, n30722, n30723, n30724, n30725, n30726,
         n30727, n30728, n30729, n30730, n30731, n30732, n30733, n30734,
         n30735, n30736, n30737, n30738, n30739, n30740, n30741, n30742,
         n30743, n30744, n30745, n30746, n30747, n30748, n30749, n30750,
         n30751, n30752, n30753, n30754, n30755, n30756, n30757, n30758,
         n30759, n30760, n30761, n30762, n30763, n30764, n30765, n30766,
         n30767, n30768, n30769, n30770, n30771, n30772, n30773, n30774,
         n30775, n30776, n30777, n30778, n30779, n30780, n30781, n30782,
         n30783, n30784, n30785, n30786, n30787, n30788, n30789, n30790,
         n30791, n30792, n30793, n30794, n30795, n30796, n30797, n30798,
         n30799, n30800, n30801, n30802, n30803, n30804, n30805, n30806,
         n30807, n30808, n30809, n30810, n30811, n30812, n30813, n30814,
         n30815, n30816, n30817, n30818, n30819, n30820, n30821, n30822,
         n30823, n30824, n30825, n30826, n30827, n30828, n30829, n30830,
         n30831, n30832, n30833, n30834, n30835, n30836, n30837, n30838,
         n30839, n30840, n30841, n30842, n30843, n30844, n30845, n30846,
         n30847, n30848, n30849, n30850, n30851, n30852, n30853, n30854,
         n30855, n30856, n30857, n30858, n30859, n30860, n30861, n30862,
         n30863, n30864, n30865, n30866, n30867, n30868, n30869, n30870,
         n30871, n30872, n30873, n30874, n30875, n30876, n30877, n30878,
         n30879, n30880, n30881, n30882, n30883, n30884, n30885, n30886,
         n30887, n30888, n30889, n30890, n30891, n30892, n30893, n30894,
         n30895, n30896, n30897, n30898, n30899, n30900, n30901, n30902,
         n30903, n30904, n30905, n30906, n30907, n30908, n30909, n30910,
         n30911, n30912, n30913, n30914, n30915, n30916, n30917, n30918,
         n30919, n30920, n30921, n30922, n30923, n30924, n30925, n30926,
         n30927, n30928, n30929, n30930, n30931, n30932, n30933, n30934,
         n30935, n30936, n30937, n30938, n30939, n30940, n30941, n30942,
         n30943, n30944, n30945, n30946, n30947, n30948, n30949, n30950,
         n30951, n30952, n30953, n30954, n30955, n30956, n30957, n30958,
         n30959, n30960, n30961, n30962, n30963, n30964, n30965, n30966,
         n30967, n30968, n30969, n30970, n30971, n30972, n30973, n30974,
         n30975, n30976, n30977, n30978, n30979, n30980, n30981, n30982,
         n30983, n30984, n30985, n30986, n30987, n30988, n30989, n30990,
         n30991, n30992, n30993, n30994, n30995, n30996, n30997, n30998,
         n30999, n31000, n31001, n31002, n31003, n31004, n31005, n31006,
         n31007, n31008, n31009, n31010, n31011, n31012, n31013, n31014,
         n31015, n31016, n31017, n31018, n31019, n31020, n31021, n31022,
         n31023, n31024, n31025, n31026, n31027, n31028, n31029, n31030,
         n31031, n31032, n31033, n31034, n31035, n31036, n31037, n31038,
         n31039, n31040, n31041, n31042, n31043, n31044, n31045, n31046,
         n31047, n31048, n31049, n31050, n31051, n31052, n31053, n31054,
         n31055, n31056, n31057, n31058, n31059, n31060, n31061, n31062,
         n31063, n31064, n31065, n31066, n31067, n31068, n31069, n31070,
         n31071, n31072, n31073, n31074, n31075, n31076, n31077, n31078,
         n31079, n31080, n31081, n31082, n31083, n31084, n31085, n31086,
         n31087, n31088, n31089, n31090, n31091, n31092, n31093, n31094,
         n31095, n31096, n31097, n31098, n31099, n31100, n31101, n31102,
         n31103, n31104, n31105, n31106, n31107, n31108, n31109, n31110,
         n31111, n31112, n31113, n31114, n31115, n31116, n31117, n31118,
         n31119, n31120, n31121, n31122, n31123, n31124, n31125, n31126,
         n31127, n31128, n31129, n31130, n31131, n31132, n31133, n31134,
         n31135, n31136, n31137, n31138, n31139, n31140, n31141, n31142,
         n31143, n31144, n31145, n31146, n31147, n31148, n31149, n31150,
         n31151, n31152, n31153, n31154, n31155, n31156, n31157, n31158,
         n31159, n31160, n31161, n31162, n31163, n31164, n31165, n31166,
         n31167, n31168, n31169, n31170, n31171, n31172, n31173, n31174,
         n31175, n31176, n31177, n31178, n31179, n31180, n31181, n31182,
         n31183, n31184, n31185, n31186, n31187, n31188, n31189, n31190,
         n31191, n31192, n31193, n31194, n31195, n31196, n31197, n31198,
         n31199, n31200, n31201, n31202, n31203, n31204, n31205, n31206,
         n31207, n31208, n31209, n31210, n31211, n31212, n31213, n31214,
         n31215, n31216, n31217, n31218, n31219, n31220, n31221, n31222,
         n31223, n31224, n31225, n31226, n31227, n31228, n31229, n31230,
         n31231, n31232, n31233, n31234, n31235, n31236, n31237, n31238,
         n31239, n31240, n31241, n31242, n31243, n31244, n31245, n31246,
         n31247, n31248, n31249, n31250, n31251, n31252, n31253, n31254,
         n31255, n31256, n31257, n31258, n31259, n31260, n31261, n31262,
         n31263, n31264, n31265, n31266, n31267, n31268, n31269, n31270,
         n31271, n31272, n31273, n31274, n31275, n31276, n31277, n31278,
         n31279, n31280, n31281, n31282, n31283, n31284, n31285, n31286,
         n31287, n31288, n31289, n31290, n31291, n31292, n31293, n31294,
         n31295, n31296, n31297, n31298, n31299, n31300, n31301, n31302,
         n31303, n31304, n31305, n31306, n31307, n31308, n31309, n31310,
         n31311, n31312, n31313, n31314, n31315, n31316, n31317, n31318,
         n31319, n31320, n31321, n31322, n31323, n31324, n31325, n31326,
         n31327, n31328, n31329, n31330, n31331, n31332, n31333, n31334,
         n31335, n31336, n31337, n31338, n31339, n31340, n31341, n31342,
         n31343, n31344, n31345, n31346, n31347, n31348, n31349, n31350,
         n31351, n31352, n31353, n31354, n31355, n31356, n31357, n31358,
         n31359, n31360, n31361, n31362, n31363, n31364, n31365, n31366,
         n31367, n31368, n31369, n31370, n31371, n31372, n31373, n31374,
         n31375, n31376, n31377, n31378, n31379, n31380, n31381, n31382,
         n31383, n31384, n31385, n31386, n31387, n31388, n31389, n31390,
         n31391, n31392, n31393, n31394, n31395, n31396, n31397, n31398,
         n31399, n31400, n31401, n31402, n31403, n31404, n31405, n31406,
         n31407, n31408, n31409, n31410, n31411, n31412, n31413, n31414,
         n31415, n31416, n31417, n31418, n31419, n31420, n31421, n31422,
         n31423, n31424, n31425, n31426, n31427, n31428, n31429, n31430,
         n31431, n31432, n31433, n31434, n31435, n31436, n31437, n31438,
         n31439, n31440, n31441, n31442, n31443, n31444, n31445, n31446,
         n31447, n31448, n31449, n31450, n31451, n31452, n31453, n31454,
         n31455, n31456, n31457, n31458, n31459, n31460, n31461, n31462,
         n31463, n31464, n31465, n31466, n31467, n31468, n31469, n31470,
         n31471, n31472, n31473, n31474, n31475, n31476, n31477, n31478,
         n31479, n31480, n31481, n31482, n31483, n31484, n31485, n31486,
         n31487, n31488, n31489, n31490, n31491, n31492, n31493, n31494,
         n31495, n31496, n31497, n31498, n31499, n31500, n31501, n31502,
         n31503, n31504, n31505, n31506, n31507, n31508, n31509, n31510,
         n31511, n31512, n31513, n31514, n31515, n31516, n31517, n31518,
         n31519, n31520, n31521, n31522, n31523, n31524, n31525, n31526,
         n31527, n31528, n31529, n31530, n31531, n31532, n31533, n31534,
         n31535, n31536, n31537, n31538, n31539, n31540, n31541, n31542,
         n31543, n31544, n31545, n31546, n31547, n31548, n31549, n31550,
         n31551, n31552, n31553, n31554, n31555, n31556, n31557, n31558,
         n31559, n31560, n31561, n31562, n31563, n31564, n31565, n31566,
         n31567, n31568, n31569, n31570, n31571, n31572, n31573, n31574,
         n31575, n31576, n31577, n31578, n31579, n31580, n31581, n31582,
         n31583, n31584, n31585, n31586, n31587, n31588, n31589, n31590,
         n31591, n31592, n31593, n31594, n31595, n31596, n31597, n31598,
         n31599, n31600, n31601, n31602, n31603, n31604, n31605, n31606,
         n31607, n31608, n31609, n31610, n31611, n31612, n31613, n31614,
         n31615, n31616, n31617, n31618, n31619, n31620, n31621, n31622,
         n31623, n31624, n31625, n31626, n31627, n31628, n31629, n31630,
         n31631, n31632, n31633, n31634, n31635, n31636, n31637, n31638,
         n31639, n31640, n31641, n31642, n31643, n31644, n31645, n31646,
         n31647, n31648, n31649, n31650, n31651, n31652, n31653, n31654,
         n31655, n31656, n31657, n31658, n31659, n31660, n31661, n31662,
         n31663, n31664, n31665, n31666, n31667, n31668, n31669, n31670,
         n31671, n31672, n31673, n31674, n31675, n31676, n31677, n31678,
         n31679, n31680, n31681, n31682, n31683, n31684, n31685, n31686,
         n31687, n31688, n31689, n31690, n31691, n31692, n31693, n31694,
         n31695, n31696, n31697, n31698, n31699, n31700, n31701, n31702,
         n31703, n31704, n31705, n31706, n31707, n31708, n31709, n31710,
         n31711, n31712, n31713, n31714, n31715, n31716, n31717, n31718,
         n31719, n31720, n31721, n31722, n31723, n31724, n31725, n31726,
         n31727, n31728, n31729, n31730, n31731, n31732, n31733, n31734,
         n31735, n31736, n31737, n31738, n31739, n31740, n31741, n31742,
         n31743, n31744, n31745, n31746, n31747, n31748, n31749, n31750,
         n31751, n31752, n31753, n31754, n31755, n31756, n31757, n31758,
         n31759, n31760, n31761, n31762, n31763, n31764, n31765, n31766,
         n31767, n31768, n31769, n31770, n31771, n31772, n31773, n31774,
         n31775, n31776, n31777, n31778, n31779, n31780, n31781, n31782,
         n31783, n31784, n31785, n31786, n31787, n31788, n31789, n31790,
         n31791, n31792, n31793, n31794, n31795, n31796, n31797, n31798,
         n31799, n31800, n31801, n31802, n31803, n31804, n31805, n31806,
         n31807, n31808, n31809, n31810, n31811, n31812, n31813, n31814,
         n31815, n31816, n31817, n31818, n31819, n31820, n31821, n31822,
         n31823, n31824, n31825, n31826, n31827, n31828, n31829, n31830,
         n31831, n31832, n31833, n31834, n31835, n31836, n31837, n31838,
         n31839, n31840, n31841, n31842, n31843, n31844, n31845, n31846,
         n31847, n31848, n31849, n31850, n31851, n31852, n31853, n31854,
         n31855, n31856, n31857, n31858, n31859, n31860, n31861, n31862,
         n31863, n31864, n31865, n31866, n31867, n31868, n31869, n31870,
         n31871, n31872, n31873, n31874, n31875, n31876, n31877, n31878,
         n31879, n31880, n31881, n31882, n31883, n31884, n31885, n31886,
         n31887, n31888, n31889, n31890, n31891, n31892, n31893, n31894,
         n31895, n31896, n31897, n31898, n31899, n31900, n31901, n31902,
         n31903, n31904, n31905, n31906, n31907, n31908, n31909, n31910,
         n31911, n31912, n31913, n31914, n31915, n31916, n31917, n31918,
         n31919, n31920, n31921, n31922, n31923, n31924, n31925, n31926,
         n31927, n31928, n31929, n31930, n31931, n31932, n31933, n31934,
         n31935, n31936, n31937, n31938, n31939, n31940, n31941, n31942,
         n31943, n31944, n31945, n31946, n31947, n31948, n31949, n31950,
         n31951, n31952, n31953, n31954, n31955, n31956, n31957, n31958,
         n31959, n31960, n31961, n31962, n31963, n31964, n31965, n31966,
         n31967, n31968, n31969, n31970, n31971, n31972, n31973, n31974,
         n31975, n31976, n31977, n31978, n31979, n31980, n31981, n31982,
         n31983, n31984, n31985, n31986, n31987, n31988, n31989, n31990,
         n31991, n31992, n31993, n31994, n31995, n31996, n31997, n31998,
         n31999, n32000, n32001, n32002, n32003, n32004, n32005, n32006,
         n32007, n32008, n32009, n32010, n32011, n32012, n32013, n32014,
         n32015, n32016, n32017, n32018, n32019, n32020, n32021, n32022,
         n32023, n32024, n32025, n32026, n32027, n32028, n32029, n32030,
         n32031, n32032, n32033, n32034, n32035, n32036, n32037, n32038,
         n32039, n32040, n32041, n32042, n32043, n32044, n32045, n32046,
         n32047, n32048, n32049, n32050, n32051, n32052, n32053, n32054,
         n32055, n32056, n32057, n32058, n32059, n32060, n32061, n32062,
         n32063, n32064, n32065, n32066, n32067, n32068, n32069, n32070,
         n32071, n32072, n32073, n32074, n32075, n32076, n32077, n32078,
         n32079, n32080, n32081, n32082, n32083, n32084, n32085, n32086,
         n32087, n32088, n32089, n32090, n32091, n32092, n32093, n32094,
         n32095, n32096, n32097, n32098, n32099, n32100, n32101, n32102,
         n32103, n32104, n32105, n32106, n32107, n32108, n32109, n32110,
         n32111, n32112, n32113, n32114, n32115, n32116, n32117, n32118,
         n32119, n32120, n32121, n32122, n32123, n32124, n32125, n32126,
         n32127, n32128, n32129, n32130, n32131, n32132, n32133, n32134,
         n32135, n32136, n32137, n32138, n32139, n32140, n32141, n32142,
         n32143, n32144, n32145, n32146, n32147, n32148, n32149, n32150,
         n32151, n32152, n32153, n32154, n32155, n32156, n32157, n32158,
         n32159, n32160, n32161, n32162, n32163, n32164, n32165, n32166,
         n32167, n32168, n32169, n32170, n32171, n32172, n32173, n32174,
         n32175, n32176, n32177, n32178, n32179, n32180, n32181, n32182,
         n32183, n32184, n32185, n32186, n32187, n32188, n32189, n32190,
         n32191, n32192, n32193, n32194, n32195, n32196, n32197, n32198,
         n32199, n32200, n32201, n32202, n32203, n32204, n32205, n32206,
         n32207, n32208, n32209, n32210, n32211, n32212, n32213, n32214,
         n32215, n32216, n32217, n32218, n32219, n32220, n32221, n32222,
         n32223, n32224, n32225, n32226, n32227, n32228, n32229, n32230,
         n32231, n32232, n32233, n32234, n32235, n32236, n32237, n32238,
         n32239, n32240, n32241, n32242, n32243, n32244, n32245, n32246,
         n32247, n32248, n32249, n32250, n32251, n32252, n32253, n32254,
         n32255, n32256, n32257, n32258, n32259, n32260, n32261, n32262,
         n32263, n32264, n32265, n32266, n32267, n32268, n32269, n32270,
         n32271, n32272, n32273, n32274, n32275, n32276, n32277, n32278,
         n32279, n32280, n32281, n32282, n32283, n32284, n32285, n32286,
         n32287, n32288, n32289, n32290, n32291, n32292, n32293, n32294,
         n32295, n32296, n32297, n32298, n32299, n32300, n32301, n32302,
         n32303, n32304, n32305, n32306, n32307, n32308, n32309, n32310,
         n32311, n32312, n32313, n32314, n32315, n32316, n32317, n32318,
         n32319, n32320, n32321, n32322, n32323, n32324, n32325, n32326,
         n32327, n32328, n32329, n32330, n32331, n32332, n32333, n32334,
         n32335, n32336, n32337, n32338, n32339, n32340, n32341, n32342,
         n32343, n32344, n32345, n32346, n32347, n32348, n32349, n32350,
         n32351, n32352, n32353, n32354, n32355, n32356, n32357, n32358,
         n32359, n32360, n32361, n32362, n32363, n32364, n32365, n32366,
         n32367, n32368, n32369, n32370, n32371, n32372, n32373, n32374,
         n32375, n32376, n32377, n32378, n32379, n32380, n32381, n32382,
         n32383, n32384, n32385, n32386, n32387, n32388, n32389, n32390,
         n32391, n32392, n32393, n32394, n32395, n32396, n32397, n32398,
         n32399, n32400, n32401, n32402, n32403, n32404, n32405, n32406,
         n32407, n32408, n32409, n32410, n32411, n32412, n32413, n32414,
         n32415, n32416, n32417, n32418, n32419, n32420, n32421, n32422,
         n32423, n32424, n32425, n32426, n32427, n32428, n32429, n32430,
         n32431, n32432, n32433, n32434, n32435, n32436, n32437, n32438,
         n32439, n32440, n32441, n32442, n32443, n32444, n32445, n32446,
         n32447, n32448, n32449, n32450, n32451, n32452, n32453, n32454,
         n32455, n32456, n32457, n32458, n32459, n32460, n32461, n32462,
         n32463, n32464, n32465, n32466, n32467, n32468, n32469, n32470,
         n32471, n32472, n32473, n32474, n32475, n32476, n32477, n32478,
         n32479, n32480, n32481, n32482, n32483, n32484, n32485, n32486,
         n32487, n32488, n32489, n32490, n32491, n32492, n32493, n32494,
         n32495, n32496, n32497, n32498, n32499, n32500, n32501, n32502,
         n32503, n32504, n32505, n32506, n32507, n32508, n32509, n32510,
         n32511, n32512, n32513, n32514, n32515, n32516, n32517, n32518,
         n32519, n32520, n32521, n32522, n32523, n32524, n32525, n32526,
         n32527, n32528, n32529, n32530, n32531, n32532, n32533, n32534,
         n32535, n32536, n32537, n32538, n32539, n32540, n32541, n32542,
         n32543, n32544, n32545, n32546, n32547, n32548, n32549, n32550,
         n32551, n32552, n32553, n32554, n32555, n32556, n32557, n32558,
         n32559, n32560, n32561, n32562, n32563, n32564, n32565, n32566,
         n32567, n32568, n32569, n32570, n32571, n32572, n32573, n32574,
         n32575, n32576, n32577, n32578, n32579, n32580, n32581, n32582,
         n32583, n32584, n32585, n32586, n32587, n32588, n32589, n32590,
         n32591, n32592, n32593, n32594, n32595, n32596, n32597, n32598,
         n32599, n32600, n32601, n32602, n32603, n32604, n32605, n32606,
         n32607, n32608, n32609, n32610, n32611, n32612, n32613, n32614,
         n32615, n32616, n32617, n32618, n32619, n32620, n32621, n32622,
         n32623, n32624, n32625, n32626, n32627, n32628, n32629, n32630,
         n32631, n32632, n32633, n32634, n32635, n32636, n32637, n32638,
         n32639, n32640, n32641, n32642, n32643, n32644, n32645, n32646,
         n32647, n32648, n32649, n32650, n32651, n32652, n32653, n32654,
         n32655, n32656, n32657, n32658, n32659, n32660, n32661, n32662,
         n32663, n32664, n32665, n32666, n32667, n32668, n32669, n32670,
         n32671, n32672, n32673, n32674, n32675, n32676, n32677, n32678,
         n32679, n32680, n32681, n32682, n32683, n32684, n32685, n32686,
         n32687, n32688, n32689, n32690, n32691, n32692, n32693, n32694,
         n32695, n32696, n32697, n32698, n32699, n32700, n32701, n32702,
         n32703, n32704, n32705, n32706, n32707, n32708, n32709, n32710,
         n32711, n32712, n32713, n32714, n32715, n32716, n32717, n32718,
         n32719, n32720, n32721, n32722, n32723, n32724, n32725, n32726,
         n32727, n32728, n32729, n32730, n32731, n32732, n32733, n32734,
         n32735, n32736, n32737, n32738, n32739, n32740, n32741, n32742,
         n32743, n32744, n32745, n32746, n32747, n32748, n32749, n32750,
         n32751, n32752, n32753, n32754, n32755, n32756, n32757, n32758,
         n32759, n32760, n32761, n32762, n32763, n32764, n32765, n32766,
         n32767, n32768, n32769, n32770, n32771, n32772, n32773, n32774,
         n32775, n32776, n32777, n32778, n32779, n32780, n32781, n32782,
         n32783, n32784, n32785, n32786, n32787, n32788, n32789, n32790,
         n32791, n32792, n32793, n32794, n32795, n32796, n32797, n32798,
         n32799, n32800, n32801, n32802, n32803, n32804, n32805, n32806,
         n32807, n32808, n32809, n32810, n32811, n32812, n32813, n32814,
         n32815, n32816, n32817, n32818, n32819, n32820, n32821, n32822,
         n32823, n32824, n32825, n32826, n32827, n32828, n32829, n32830,
         n32831, n32832, n32833, n32834, n32835, n32836, n32837, n32838,
         n32839, n32840, n32841, n32842, n32843, n32844, n32845, n32846,
         n32847, n32848, n32849, n32850, n32851, n32852, n32853, n32854,
         n32855, n32856, n32857, n32858, n32859, n32860, n32861, n32862,
         n32863, n32864, n32865, n32866, n32867, n32868, n32869, n32870,
         n32871, n32872, n32873, n32874, n32875, n32876, n32877, n32878,
         n32879, n32880, n32881, n32882, n32883, n32884, n32885, n32886,
         n32887, n32888, n32889, n32890, n32891, n32892, n32893, n32894,
         n32895, n32896, n32897, n32898, n32899, n32900, n32901, n32902,
         n32903, n32904, n32905, n32906, n32907, n32908, n32909, n32910,
         n32911, n32912, n32913, n32914, n32915, n32916, n32917, n32918,
         n32919, n32920, n32921, n32922, n32923, n32924, n32925, n32926,
         n32927, n32928, n32929, n32930, n32931, n32932, n32933, n32934,
         n32935, n32936, n32937, n32938, n32939, n32940, n32941, n32942,
         n32943, n32944, n32945, n32946, n32947, n32948, n32949, n32950,
         n32951, n32952, n32953, n32954, n32955, n32956, n32957, n32958,
         n32959, n32960, n32961, n32962, n32963, n32964, n32965, n32966,
         n32967, n32968, n32969, n32970, n32971, n32972, n32973, n32974,
         n32975, n32976, n32977, n32978, n32979, n32980, n32981, n32982,
         n32983, n32984, n32985, n32986, n32987, n32988, n32989, n32990,
         n32991, n32992, n32993, n32994, n32995, n32996, n32997, n32998,
         n32999, n33000, n33001, n33002, n33003, n33004, n33005, n33006,
         n33007, n33008, n33009, n33010, n33011, n33012, n33013, n33014,
         n33015, n33016, n33017, n33018, n33019, n33020, n33021, n33022,
         n33023, n33024, n33025, n33026, n33027, n33028, n33029, n33030,
         n33031, n33032, n33033, n33034, n33035, n33036, n33037, n33038,
         n33039, n33040, n33041, n33042, n33043, n33044, n33045, n33046,
         n33047, n33048, n33049, n33050, n33051, n33052, n33053, n33054,
         n33055, n33056, n33057, n33058, n33059, n33060, n33061, n33062,
         n33063, n33064, n33065, n33066, n33067, n33068, n33069, n33070,
         n33071, n33072, n33073, n33074, n33075, n33076, n33077, n33078,
         n33079, n33080, n33081, n33082, n33083, n33084, n33085, n33086,
         n33087, n33088, n33089, n33090, n33091, n33092, n33093, n33094,
         n33095, n33096, n33097, n33098, n33099, n33100, n33101, n33102,
         n33103, n33104, n33105, n33106, n33107, n33108, n33109, n33110,
         n33111, n33112, n33113, n33114, n33115, n33116, n33117, n33118,
         n33119, n33120, n33121, n33122, n33123, n33124, n33125, n33126,
         n33127, n33128, n33129, n33130, n33131, n33132, n33133, n33134,
         n33135, n33136, n33137, n33138, n33139, n33140, n33141, n33142,
         n33143, n33144, n33145, n33146, n33147, n33148, n33149, n33150,
         n33151, n33152, n33153, n33154, n33155, n33156, n33157, n33158,
         n33159, n33160, n33161, n33162, n33163, n33164, n33165, n33166,
         n33167, n33168, n33169, n33170, n33171, n33172, n33173, n33174,
         n33175, n33176, n33177, n33178, n33179, n33180, n33181, n33182,
         n33183, n33184, n33185, n33186, n33187, n33188, n33189, n33190,
         n33191, n33192, n33193, n33194, n33195, n33196, n33197, n33198,
         n33199, n33200, n33201, n33202, n33203, n33204, n33205, n33206,
         n33207, n33208, n33209, n33210, n33211, n33212, n33213, n33214,
         n33215, n33216, n33217, n33218, n33219, n33220, n33221, n33222,
         n33223, n33224, n33225, n33226, n33227, n33228, n33229, n33230,
         n33231, n33232, n33233, n33234, n33235, n33236, n33237, n33238,
         n33239, n33240, n33241, n33242, n33243, n33244, n33245, n33246,
         n33247, n33248, n33249, n33250, n33251, n33252, n33253, n33254,
         n33255, n33256, n33257, n33258, n33259, n33260, n33261, n33262,
         n33263, n33264, n33265, n33266, n33267, n33268, n33269, n33270,
         n33271, n33272, n33273, n33274, n33275, n33276, n33277, n33278,
         n33279, n33280, n33281, n33282, n33283, n33284, n33285, n33286,
         n33287, n33288, n33289, n33290, n33291, n33292, n33293, n33294,
         n33295, n33296, n33297, n33298, n33299, n33300, n33301, n33302,
         n33303, n33304, n33305, n33306, n33307, n33308, n33309, n33310,
         n33311, n33312, n33313, n33314, n33315, n33316, n33317, n33318,
         n33319, n33320, n33321, n33322, n33323, n33324, n33325, n33326,
         n33327, n33328, n33329, n33330, n33331, n33332, n33333, n33334,
         n33335, n33336, n33337, n33338, n33339, n33340, n33341, n33342,
         n33343, n33344, n33345, n33346, n33347, n33348, n33349, n33350,
         n33351, n33352, n33353, n33354, n33355, n33356, n33357, n33358,
         n33359, n33360, n33361, n33362, n33363, n33364, n33365, n33366,
         n33367, n33368, n33369, n33370, n33371, n33372, n33373, n33374,
         n33375, n33376, n33377, n33378, n33379, n33380, n33381, n33382,
         n33383, n33384, n33385, n33386, n33387, n33388, n33389, n33390,
         n33391, n33392, n33393, n33394, n33395, n33396, n33397, n33398,
         n33399, n33400, n33401, n33402, n33403, n33404, n33405, n33406,
         n33407, n33408, n33409, n33410, n33411, n33412, n33413, n33414,
         n33415, n33416, n33417, n33418, n33419, n33420, n33421, n33422,
         n33423, n33424, n33425, n33426, n33427, n33428, n33429, n33430,
         n33431, n33432, n33433, n33434, n33435, n33436, n33437, n33438,
         n33439, n33440, n33441, n33442, n33443, n33444, n33445, n33446,
         n33447, n33448, n33449, n33450, n33451, n33452, n33453, n33454,
         n33455, n33456, n33457, n33458, n33459, n33460, n33461, n33462,
         n33463, n33464, n33465, n33466, n33467, n33468, n33469, n33470,
         n33471, n33472, n33473, n33474, n33475, n33476, n33477, n33478,
         n33479, n33480, n33481, n33482, n33483, n33484, n33485, n33486,
         n33487, n33488, n33489, n33490, n33491, n33492, n33493, n33494,
         n33495, n33496, n33497, n33498, n33499, n33500, n33501, n33502,
         n33503, n33504, n33505, n33506, n33507, n33508, n33509, n33510,
         n33511, n33512, n33513, n33514, n33515, n33516, n33517, n33518,
         n33519, n33520, n33521, n33522, n33523, n33524, n33525, n33526,
         n33527, n33528, n33529, n33530, n33531, n33532, n33533, n33534,
         n33535, n33536, n33537, n33538, n33539, n33540, n33541, n33542,
         n33543, n33544, n33545, n33546, n33547, n33548, n33549, n33550,
         n33551, n33552, n33553, n33554, n33555, n33556, n33557, n33558,
         n33559, n33560, n33561, n33562, n33563, n33564, n33565, n33566,
         n33567, n33568, n33569, n33570, n33571, n33572, n33573, n33574,
         n33575, n33576, n33577, n33578, n33579, n33580, n33581, n33582,
         n33583, n33584, n33585, n33586, n33587, n33588, n33589, n33590,
         n33591, n33592, n33593, n33594, n33595, n33596, n33597, n33598,
         n33599, n33600, n33601, n33602, n33603, n33604, n33605, n33606,
         n33607, n33608, n33609, n33610, n33611, n33612, n33613, n33614,
         n33615, n33616, n33617, n33618, n33619, n33620, n33621, n33622,
         n33623, n33624, n33625, n33626, n33627, n33628, n33629, n33630,
         n33631, n33632, n33633, n33634, n33635, n33636, n33637, n33638,
         n33639, n33640, n33641, n33642, n33643, n33644, n33645, n33646,
         n33647, n33648, n33649, n33650, n33651, n33652, n33653, n33654,
         n33655, n33656, n33657, n33658, n33659, n33660, n33661, n33662,
         n33663, n33664, n33665, n33666, n33667, n33668, n33669, n33670,
         n33671, n33672, n33673, n33674, n33675, n33676, n33677, n33678,
         n33679, n33680, n33681, n33682, n33683, n33684, n33685, n33686,
         n33687, n33688, n33689, n33690, n33691, n33692, n33693, n33694,
         n33695, n33696, n33697, n33698, n33699, n33700, n33701, n33702,
         n33703, n33704, n33705, n33706, n33707, n33708, n33709, n33710,
         n33711, n33712, n33713, n33714, n33715, n33716, n33717, n33718,
         n33719, n33720, n33721, n33722, n33723, n33724, n33725, n33726,
         n33727, n33728, n33729, n33730, n33731, n33732, n33733, n33734,
         n33735, n33736, n33737, n33738, n33739, n33740, n33741, n33742,
         n33743, n33744, n33745, n33746, n33747, n33748, n33749, n33750,
         n33751, n33752, n33753, n33754, n33755, n33756, n33757, n33758,
         n33759, n33760, n33761, n33762, n33763, n33764, n33765, n33766,
         n33767, n33768, n33769, n33770, n33771, n33772, n33773, n33774,
         n33775, n33776, n33777, n33778, n33779, n33780, n33781, n33782,
         n33783, n33784, n33785, n33786, n33787, n33788, n33789, n33790,
         n33791, n33792, n33793, n33794, n33795, n33796, n33797, n33798,
         n33799, n33800, n33801, n33802, n33803, n33804, n33805, n33806,
         n33807, n33808, n33809, n33810, n33811, n33812, n33813, n33814,
         n33815, n33816, n33817, n33818, n33819, n33820, n33821, n33822,
         n33823, n33824, n33825, n33826, n33827, n33828, n33829, n33830,
         n33831, n33832, n33833, n33834, n33835, n33836, n33837, n33838,
         n33839, n33840, n33841, n33842, n33843, n33844, n33845, n33846,
         n33847, n33848, n33849, n33850, n33851, n33852, n33853, n33854,
         n33855, n33856, n33857, n33858, n33859, n33860, n33861, n33862,
         n33863, n33864, n33865, n33866, n33867, n33868, n33869, n33870,
         n33871, n33872, n33873, n33874, n33875, n33876, n33877, n33878,
         n33879, n33880, n33881, n33882, n33883, n33884, n33885, n33886,
         n33887, n33888, n33889, n33890, n33891, n33892, n33893, n33894,
         n33895, n33896, n33897, n33898, n33899, n33900, n33901, n33902,
         n33903, n33904, n33905, n33906, n33907, n33908, n33909, n33910,
         n33911, n33912, n33913, n33914, n33915, n33916, n33917, n33918,
         n33919, n33920, n33921, n33922, n33923, n33924, n33925, n33926,
         n33927, n33928, n33929, n33930, n33931, n33932, n33933, n33934,
         n33935, n33936, n33937, n33938, n33939, n33940, n33941, n33942,
         n33943, n33944, n33945, n33946, n33947, n33948, n33949, n33950,
         n33951, n33952, n33953, n33954, n33955, n33956, n33957, n33958,
         n33959, n33960, n33961, n33962, n33963, n33964, n33965, n33966,
         n33967, n33968, n33969, n33970, n33971, n33972, n33973, n33974,
         n33975, n33976, n33977, n33978, n33979, n33980, n33981, n33982,
         n33983, n33984, n33985, n33986, n33987, n33988, n33989, n33990,
         n33991, n33992, n33993, n33994, n33995, n33996, n33997, n33998,
         n33999, n34000, n34001, n34002, n34003, n34004, n34005, n34006,
         n34007, n34008, n34009, n34010, n34011, n34012, n34013, n34014,
         n34015, n34016, n34017, n34018, n34019, n34020, n34021, n34022,
         n34023, n34024, n34025, n34026, n34027, n34028, n34029, n34030,
         n34031, n34032, n34033, n34034, n34035, n34036, n34037, n34038,
         n34039, n34040, n34041, n34042, n34043, n34044, n34045, n34046,
         n34047, n34048, n34049, n34050, n34051, n34052, n34053, n34054,
         n34055, n34056, n34057, n34058, n34059, n34060, n34061, n34062,
         n34063, n34064, n34065, n34066, n34067, n34068, n34069, n34070,
         n34071, n34072, n34073, n34074, n34075, n34076, n34077, n34078,
         n34079, n34080, n34081, n34082, n34083, n34084, n34085, n34086,
         n34087, n34088, n34089, n34090, n34091, n34092, n34093, n34094,
         n34095, n34096, n34097, n34098, n34099, n34100, n34101, n34102,
         n34103, n34104, n34105, n34106, n34107, n34108, n34109, n34110,
         n34111, n34112, n34113, n34114, n34115, n34116, n34117, n34118,
         n34119, n34120, n34121, n34122, n34123, n34124, n34125, n34126,
         n34127, n34128, n34129, n34130, n34131, n34132, n34133, n34134,
         n34135, n34136, n34137, n34138, n34139, n34140, n34141, n34142,
         n34143, n34144, n34145, n34146, n34147, n34148, n34149, n34150,
         n34151, n34152, n34153, n34154, n34155, n34156, n34157, n34158,
         n34159, n34160, n34161, n34162, n34163, n34164, n34165, n34166,
         n34167, n34168, n34169, n34170, n34171, n34172, n34173, n34174,
         n34175, n34176, n34177, n34178, n34179, n34180, n34181, n34182,
         n34183, n34184, n34185, n34186, n34187, n34188, n34189, n34190,
         n34191, n34192, n34193, n34194, n34195, n34196, n34197, n34198,
         n34199, n34200, n34201, n34202, n34203, n34204, n34205, n34206,
         n34207, n34208, n34209, n34210, n34211, n34212, n34213, n34214,
         n34215, n34216, n34217, n34218, n34219, n34220, n34221, n34222,
         n34223, n34224, n34225, n34226, n34227, n34228, n34229, n34230,
         n34231, n34232, n34233, n34234, n34235, n34236, n34237, n34238,
         n34239, n34240, n34241, n34242, n34243, n34244, n34245, n34246,
         n34247, n34248, n34249, n34250, n34251, n34252, n34253, n34254,
         n34255, n34256, n34257, n34258, n34259, n34260, n34261, n34262,
         n34263, n34264, n34265, n34266, n34267, n34268, n34269, n34270,
         n34271, n34272, n34273, n34274, n34275, n34276, n34277, n34278,
         n34279, n34280, n34281, n34282, n34283, n34284, n34285, n34286,
         n34287, n34288, n34289, n34290, n34291, n34292, n34293, n34294,
         n34295, n34296, n34297, n34298, n34299, n34300, n34301, n34302,
         n34303, n34304, n34305, n34306, n34307, n34308, n34309, n34310,
         n34311, n34312, n34313, n34314, n34315, n34316, n34317, n34318,
         n34319, n34320, n34321, n34322, n34323, n34324, n34325, n34326,
         n34327, n34328, n34329, n34330, n34331, n34332, n34333, n34334,
         n34335, n34336, n34337, n34338, n34339, n34340, n34341, n34342,
         n34343, n34344, n34345, n34346, n34347, n34348, n34349, n34350,
         n34351, n34352, n34353, n34354, n34355, n34356, n34357, n34358,
         n34359, n34360, n34361, n34362, n34363, n34364, n34365, n34366,
         n34367, n34368, n34369, n34370, n34371, n34372, n34373, n34374,
         n34375, n34376, n34377, n34378, n34379, n34380, n34381, n34382,
         n34383, n34384, n34385, n34386, n34387, n34388, n34389, n34390,
         n34391, n34392, n34393, n34394, n34395, n34396, n34397, n34398,
         n34399, n34400, n34401, n34402, n34403, n34404, n34405, n34406,
         n34407, n34408, n34409, n34410, n34411, n34412, n34413, n34414,
         n34415, n34416, n34417, n34418, n34419, n34420, n34421, n34422,
         n34423, n34424, n34425, n34426, n34427, n34428, n34429, n34430,
         n34431, n34432, n34433, n34434, n34435, n34436, n34437, n34438,
         n34439, n34440, n34441, n34442, n34443, n34444, n34445, n34446,
         n34447, n34448, n34449, n34450, n34451, n34452, n34453, n34454,
         n34455, n34456, n34457, n34458, n34459, n34460, n34461, n34462,
         n34463, n34464, n34465, n34466, n34467, n34468, n34469, n34470,
         n34471, n34472, n34473, n34474, n34475, n34476, n34477, n34478,
         n34479, n34480, n34481, n34482, n34483, n34484, n34485, n34486,
         n34487, n34488, n34489, n34490, n34491, n34492, n34493, n34494,
         n34495, n34496, n34497, n34498, n34499, n34500, n34501, n34502,
         n34503, n34504, n34505, n34506, n34507, n34508, n34509, n34510,
         n34511, n34512, n34513, n34514, n34515, n34516, n34517, n34518,
         n34519, n34520, n34521, n34522, n34523, n34524, n34525, n34526,
         n34527, n34528, n34529, n34530, n34531, n34532, n34533, n34534,
         n34535, n34536, n34537, n34538, n34539, n34540, n34541, n34542,
         n34543, n34544, n34545, n34546, n34547, n34548, n34549, n34550,
         n34551, n34552, n34553, n34554, n34555, n34556, n34557, n34558,
         n34559, n34560, n34561, n34562, n34563, n34564, n34565, n34566,
         n34567, n34568, n34569, n34570, n34571, n34572, n34573, n34574,
         n34575, n34576, n34577, n34578, n34579, n34580, n34581, n34582,
         n34583, n34584, n34585, n34586, n34587, n34588, n34589, n34590,
         n34591, n34592, n34593, n34594, n34595, n34596, n34597, n34598,
         n34599, n34600, n34601, n34602, n34603, n34604, n34605, n34606,
         n34607, n34608, n34609, n34610, n34611, n34612, n34613, n34614,
         n34615, n34616, n34617, n34618, n34619, n34620, n34621, n34622,
         n34623, n34624, n34625, n34626, n34627, n34628, n34629, n34630,
         n34631, n34632, n34633, n34634, n34635, n34636, n34637, n34638,
         n34639, n34640, n34641, n34642, n34643, n34644, n34645, n34646,
         n34647, n34648, n34649, n34650, n34651, n34652, n34653, n34654,
         n34655, n34656, n34657, n34658, n34659, n34660, n34661, n34662,
         n34663, n34664, n34665, n34666, n34667, n34668, n34669, n34670,
         n34671, n34672, n34673, n34674, n34675, n34676, n34677, n34678,
         n34679, n34680, n34681, n34682, n34683, n34684, n34685, n34686,
         n34687, n34688, n34689, n34690, n34691, n34692, n34693, n34694,
         n34695, n34696, n34697, n34698, n34699, n34700, n34701, n34702,
         n34703, n34704, n34705, n34706, n34707, n34708, n34709, n34710,
         n34711, n34712, n34713, n34714, n34715, n34716, n34717, n34718,
         n34719, n34720, n34721, n34722, n34723, n34724, n34725, n34726,
         n34727, n34728, n34729, n34730, n34731, n34732, n34733, n34734,
         n34735, n34736, n34737, n34738, n34739, n34740, n34741, n34742,
         n34743, n34744, n34745, n34746, n34747, n34748, n34749, n34750,
         n34751, n34752, n34753, n34754, n34755, n34756, n34757, n34758,
         n34759, n34760, n34761, n34762, n34763, n34764, n34765, n34766,
         n34767, n34768, n34769, n34770, n34771, n34772, n34773, n34774,
         n34775, n34776, n34777, n34778, n34779, n34780, n34781, n34782,
         n34783, n34784, n34785, n34786, n34787, n34788, n34789, n34790,
         n34791, n34792, n34793, n34794, n34795, n34796, n34797, n34798,
         n34799, n34800, n34801, n34802, n34803, n34804, n34805, n34806,
         n34807, n34808, n34809, n34810, n34811, n34812, n34813, n34814,
         n34815, n34816, n34817, n34818, n34819, n34820, n34821, n34822,
         n34823, n34824, n34825, n34826, n34827, n34828, n34829, n34830,
         n34831, n34832, n34833, n34834, n34835, n34836, n34837, n34838,
         n34839, n34840, n34841, n34842, n34843, n34844, n34845, n34846,
         n34847, n34848, n34849, n34850, n34851, n34852, n34853, n34854,
         n34855, n34856, n34857, n34858, n34859, n34860, n34861, n34862,
         n34863, n34864, n34865, n34866, n34867, n34868, n34869, n34870,
         n34871, n34872, n34873, n34874, n34875, n34876, n34877, n34878,
         n34879, n34880, n34881, n34882, n34883, n34884, n34885, n34886,
         n34887, n34888, n34889, n34890, n34891, n34892, n34893, n34894,
         n34895, n34896, n34897, n34898, n34899, n34900, n34901, n34902,
         n34903, n34904, n34905, n34906, n34907, n34908, n34909, n34910,
         n34911, n34912, n34913, n34914, n34915, n34916, n34917, n34918,
         n34919, n34920, n34921, n34922, n34923, n34924, n34925, n34926,
         n34927, n34928, n34929, n34930, n34931, n34932, n34933, n34934,
         n34935, n34936, n34937, n34938, n34939, n34940, n34941, n34942,
         n34943, n34944, n34945, n34946, n34947, n34948, n34949, n34950,
         n34951, n34952, n34953, n34954, n34955, n34956, n34957, n34958,
         n34959, n34960, n34961, n34962, n34963, n34964, n34965, n34966,
         n34967, n34968, n34969, n34970, n34971, n34972, n34973, n34974,
         n34975, n34976, n34977, n34978, n34979, n34980, n34981, n34982,
         n34983, n34984, n34985, n34986, n34987, n34988, n34989, n34990,
         n34991, n34992, n34993, n34994, n34995, n34996, n34997, n34998,
         n34999, n35000, n35001, n35002, n35003, n35004, n35005, n35006,
         n35007, n35008, n35009, n35010, n35011, n35012, n35013, n35014,
         n35015, n35016, n35017, n35018, n35019, n35020, n35021, n35022,
         n35023, n35024, n35025, n35026, n35027, n35028, n35029, n35030,
         n35031, n35032, n35033, n35034, n35035, n35036, n35037, n35038,
         n35039, n35040, n35041, n35042, n35043, n35044, n35045, n35046,
         n35047, n35048, n35049, n35050, n35051, n35052, n35053, n35054,
         n35055, n35056, n35057, n35058, n35059, n35060, n35061, n35062,
         n35063, n35064, n35065, n35066, n35067, n35068, n35069, n35070,
         n35071, n35072, n35073, n35074, n35075, n35076, n35077, n35078,
         n35079, n35080, n35081, n35082, n35083, n35084, n35085, n35086,
         n35087, n35088, n35089, n35090, n35091, n35092, n35093, n35094,
         n35095, n35096, n35097, n35098, n35099, n35100, n35101, n35102,
         n35103, n35104, n35105, n35106, n35107, n35108, n35109, n35110,
         n35111, n35112, n35113, n35114, n35115, n35116, n35117, n35118,
         n35119, n35120, n35121, n35122, n35123, n35124, n35125, n35126,
         n35127, n35128, n35129, n35130, n35131, n35132, n35133, n35134,
         n35135, n35136, n35137, n35138, n35139, n35140, n35141, n35142,
         n35143, n35144, n35145, n35146, n35147, n35148, n35149, n35150,
         n35151, n35152, n35153, n35154, n35155, n35156, n35157, n35158,
         n35159, n35160, n35161, n35162, n35163, n35164, n35165, n35166,
         n35167, n35168, n35169, n35170, n35171, n35172, n35173, n35174,
         n35175, n35176, n35177, n35178, n35179, n35180, n35181, n35182,
         n35183, n35184, n35185, n35186, n35187, n35188, n35189, n35190,
         n35191, n35192, n35193, n35194, n35195, n35196, n35197, n35198,
         n35199, n35200, n35201, n35202, n35203, n35204, n35205, n35206,
         n35207, n35208, n35209, n35210, n35211, n35212, n35213, n35214,
         n35215, n35216, n35217, n35218, n35219, n35220, n35221, n35222,
         n35223, n35224, n35225, n35226, n35227, n35228, n35229, n35230,
         n35231, n35232, n35233, n35234, n35235, n35236, n35237, n35238,
         n35239, n35240, n35241, n35242, n35243, n35244, n35245, n35246,
         n35247, n35248, n35249, n35250, n35251, n35252, n35253, n35254,
         n35255, n35256, n35257, n35258, n35259, n35260, n35261, n35262,
         n35263, n35264, n35265, n35266, n35267, n35268, n35269, n35270,
         n35271, n35272, n35273, n35274, n35275, n35276, n35277, n35278,
         n35279, n35280, n35281, n35282, n35283, n35284, n35285, n35286,
         n35287, n35288, n35289, n35290, n35291, n35292, n35293, n35294,
         n35295, n35296, n35297, n35298, n35299, n35300, n35301, n35302,
         n35303, n35304, n35305, n35306, n35307, n35308, n35309, n35310,
         n35311, n35312, n35313, n35314, n35315, n35316, n35317, n35318,
         n35319, n35320, n35321, n35322, n35323, n35324, n35325, n35326,
         n35327, n35328, n35329, n35330, n35331, n35332, n35333, n35334,
         n35335, n35336, n35337, n35338, n35339, n35340, n35341, n35342,
         n35343, n35344, n35345, n35346, n35347, n35348, n35349, n35350,
         n35351, n35352, n35353, n35354, n35355, n35356, n35357, n35358,
         n35359, n35360, n35361, n35362, n35363, n35364, n35365, n35366,
         n35367, n35368, n35369, n35370, n35371, n35372, n35373, n35374,
         n35375, n35376, n35377, n35378, n35379, n35380, n35381, n35382,
         n35383, n35384, n35385, n35386, n35387, n35388, n35389, n35390,
         n35391, n35392, n35393, n35394, n35395, n35396, n35397, n35398,
         n35399, n35400, n35401, n35402, n35403, n35404, n35405, n35406,
         n35407, n35408, n35409, n35410, n35411, n35412, n35413, n35414,
         n35415, n35416, n35417, n35418, n35419, n35420, n35421, n35422,
         n35423, n35424, n35425, n35426, n35427, n35428, n35429, n35430,
         n35431, n35432, n35433, n35434, n35435, n35436, n35437, n35438,
         n35439, n35440, n35441, n35442, n35443, n35444, n35445, n35446,
         n35447, n35448, n35449, n35450, n35451, n35452, n35453, n35454,
         n35455, n35456, n35457, n35458, n35459, n35460, n35461, n35462,
         n35463, n35464, n35465, n35466, n35467, n35468, n35469, n35470,
         n35471, n35472, n35473, n35474, n35475, n35476, n35477, n35478,
         n35479, n35480, n35481, n35482, n35483, n35484, n35485, n35486,
         n35487, n35488, n35489, n35490, n35491, n35492, n35493, n35494,
         n35495, n35496, n35497, n35498, n35499, n35500, n35501, n35502,
         n35503, n35504, n35505, n35506, n35507, n35508, n35509, n35510,
         n35511, n35512, n35513, n35514, n35515, n35516, n35517, n35518,
         n35519, n35520, n35521, n35522, n35523, n35524, n35525, n35526,
         n35527, n35528, n35529, n35530, n35531, n35532, n35533, n35534,
         n35535, n35536, n35537, n35538, n35539, n35540, n35541, n35542,
         n35543, n35544, n35545, n35546, n35547, n35548, n35549, n35550,
         n35551, n35552, n35553, n35554, n35555, n35556, n35557, n35558,
         n35559, n35560, n35561, n35562, n35563, n35564, n35565, n35566,
         n35567, n35568, n35569, n35570, n35571, n35572, n35573, n35574,
         n35575, n35576, n35577, n35578, n35579, n35580, n35581, n35582,
         n35583, n35584, n35585, n35586, n35587, n35588, n35589, n35590,
         n35591, n35592, n35593, n35594, n35595, n35596, n35597, n35598,
         n35599, n35600, n35601, n35602, n35603, n35604, n35605, n35606,
         n35607, n35608, n35609, n35610, n35611, n35612, n35613, n35614,
         n35615, n35616, n35617, n35618, n35619, n35620, n35621, n35622,
         n35623, n35624, n35625, n35626, n35627, n35628, n35629, n35630,
         n35631, n35632, n35633, n35634, n35635, n35636, n35637, n35638,
         n35639, n35640, n35641, n35642, n35643, n35644, n35645, n35646,
         n35647, n35648, n35649, n35650, n35651, n35652, n35653, n35654,
         n35655, n35656, n35657, n35658, n35659, n35660, n35661, n35662,
         n35663, n35664, n35665, n35666, n35667, n35668, n35669, n35670,
         n35671, n35672, n35673, n35674, n35675, n35676, n35677, n35678,
         n35679, n35680, n35681, n35682, n35683, n35684, n35685, n35686,
         n35687, n35688, n35689, n35690, n35691, n35692, n35693, n35694,
         n35695, n35696, n35697, n35698, n35699, n35700, n35701, n35702,
         n35703, n35704, n35705, n35706, n35707, n35708, n35709, n35710,
         n35711, n35712, n35713, n35714, n35715, n35716, n35717, n35718,
         n35719, n35720, n35721, n35722, n35723, n35724, n35725, n35726,
         n35727, n35728, n35729, n35730, n35731, n35732, n35733, n35734,
         n35735, n35736, n35737, n35738, n35739, n35740, n35741, n35742,
         n35743, n35744, n35745, n35746, n35747, n35748, n35749, n35750,
         n35751, n35752, n35753, n35754, n35755, n35756, n35757, n35758,
         n35759, n35760, n35761, n35762, n35763, n35764, n35765, n35766,
         n35767, n35768, n35769, n35770, n35771, n35772, n35773, n35774,
         n35775, n35776, n35777, n35778, n35779, n35780, n35781, n35782,
         n35783, n35784, n35785, n35786, n35787, n35788, n35789, n35790,
         n35791, n35792, n35793, n35794, n35795, n35796, n35797, n35798,
         n35799, n35800, n35801, n35802, n35803, n35804, n35805, n35806,
         n35807, n35808, n35809, n35810, n35811, n35812, n35813, n35814,
         n35815, n35816, n35817, n35818, n35819, n35820, n35821, n35822,
         n35823, n35824, n35825, n35826, n35827, n35828, n35829, n35830,
         n35831, n35832, n35833, n35834, n35835, n35836, n35837, n35838,
         n35839, n35840, n35841, n35842, n35843, n35844, n35845, n35846,
         n35847, n35848, n35849, n35850, n35851, n35852, n35853, n35854,
         n35855, n35856, n35857, n35858, n35859, n35860, n35861, n35862,
         n35863, n35864, n35865, n35866, n35867, n35868, n35869, n35870,
         n35871, n35872, n35873, n35874, n35875, n35876, n35877, n35878,
         n35879, n35880, n35881, n35882, n35883, n35884, n35885, n35886,
         n35887, n35888, n35889, n35890, n35891, n35892, n35893, n35894,
         n35895, n35896, n35897, n35898, n35899, n35900, n35901, n35902,
         n35903, n35904, n35905, n35906, n35907, n35908, n35909, n35910,
         n35911, n35912, n35913, n35914, n35915, n35916, n35917, n35918,
         n35919, n35920, n35921, n35922, n35923, n35924, n35925, n35926,
         n35927, n35928, n35929, n35930, n35931, n35932, n35933, n35934,
         n35935, n35936, n35937, n35938, n35939, n35940, n35941, n35942,
         n35943, n35944, n35945, n35946, n35947, n35948, n35949, n35950,
         n35951, n35952, n35953, n35954, n35955, n35956, n35957, n35958,
         n35959, n35960, n35961, n35962, n35963, n35964, n35965, n35966,
         n35967, n35968, n35969, n35970, n35971, n35972, n35973, n35974,
         n35975, n35976, n35977, n35978, n35979, n35980, n35981, n35982,
         n35983, n35984, n35985, n35986, n35987, n35988, n35989, n35990,
         n35991, n35992, n35993, n35994, n35995, n35996, n35997, n35998,
         n35999, n36000, n36001, n36002, n36003, n36004, n36005, n36006,
         n36007, n36008, n36009, n36010, n36011, n36012, n36013, n36014,
         n36015, n36016, n36017, n36018, n36019, n36020, n36021, n36022,
         n36023, n36024, n36025, n36026, n36027, n36028, n36029, n36030,
         n36031, n36032, n36033, n36034, n36035, n36036, n36037, n36038,
         n36039, n36040, n36041, n36042, n36043, n36044, n36045, n36046,
         n36047, n36048, n36049, n36050, n36051, n36052, n36053, n36054,
         n36055, n36056, n36057, n36058, n36059, n36060, n36061, n36062,
         n36063, n36064, n36065, n36066, n36067, n36068, n36069, n36070,
         n36071, n36072, n36073, n36074, n36075, n36076, n36077, n36078,
         n36079, n36080, n36081, n36082, n36083, n36084, n36085, n36086,
         n36087, n36088, n36089, n36090, n36091, n36092, n36093, n36094,
         n36095, n36096, n36097, n36098, n36099, n36100, n36101, n36102,
         n36103, n36104, n36105, n36106, n36107, n36108, n36109, n36110,
         n36111, n36112, n36113, n36114, n36115, n36116, n36117, n36118,
         n36119, n36120, n36121, n36122, n36123, n36124, n36125, n36126,
         n36127, n36128, n36129, n36130, n36131, n36132, n36133, n36134,
         n36135, n36136, n36137, n36138, n36139, n36140, n36141, n36142,
         n36143, n36144, n36145, n36146, n36147, n36148, n36149, n36150,
         n36151, n36152, n36153, n36154, n36155, n36156, n36157, n36158,
         n36159, n36160, n36161, n36162, n36163, n36164, n36165, n36166,
         n36167, n36168, n36169, n36170, n36171, n36172, n36173, n36174,
         n36175, n36176, n36177, n36178, n36179, n36180, n36181, n36182,
         n36183, n36184, n36185, n36186, n36187, n36188, n36189, n36190,
         n36191, n36192, n36193, n36194, n36195, n36196, n36197, n36198,
         n36199, n36200, n36201, n36202, n36203, n36204, n36205, n36206,
         n36207, n36208, n36209, n36210, n36211, n36212, n36213, n36214,
         n36215, n36216, n36217, n36218, n36219, n36220, n36221, n36222,
         n36223, n36224, n36225, n36226, n36227, n36228, n36229, n36230,
         n36231, n36232, n36233, n36234, n36235, n36236, n36237, n36238,
         n36239, n36240, n36241, n36242, n36243, n36244, n36245, n36246,
         n36247, n36248, n36249, n36250, n36251, n36252, n36253, n36254,
         n36255, n36256, n36257, n36258, n36259, n36260, n36261, n36262,
         n36263, n36264, n36265, n36266, n36267, n36268, n36269, n36270,
         n36271, n36272, n36273, n36274, n36275, n36276, n36277, n36278,
         n36279, n36280, n36281, n36282, n36283, n36284, n36285, n36286,
         n36287, n36288, n36289, n36290, n36291, n36292, n36293, n36294,
         n36295, n36296, n36297, n36298, n36299, n36300, n36301, n36302,
         n36303, n36304, n36305, n36306, n36307, n36308, n36309, n36310,
         n36311, n36312, n36313, n36314, n36315, n36316, n36317, n36318,
         n36319, n36320, n36321, n36322, n36323, n36324, n36325, n36326,
         n36327, n36328, n36329, n36330, n36331, n36332, n36333, n36334,
         n36335, n36336, n36337, n36338, n36339, n36340, n36341, n36342,
         n36343, n36344, n36345, n36346, n36347, n36348, n36349, n36350,
         n36351, n36352, n36353, n36354, n36355, n36356, n36357, n36358,
         n36359, n36360, n36361, n36362, n36363, n36364, n36365, n36366,
         n36367, n36368, n36369, n36370, n36371, n36372, n36373, n36374,
         n36375, n36376, n36377, n36378, n36379, n36380, n36381, n36382,
         n36383, n36384, n36385, n36386, n36387, n36388, n36389, n36390,
         n36391, n36392, n36393, n36394, n36395, n36396, n36397, n36398,
         n36399, n36400, n36401, n36402, n36403, n36404, n36405, n36406,
         n36407, n36408, n36409, n36410, n36411, n36412, n36413, n36414,
         n36415, n36416, n36417, n36418, n36419, n36420, n36421, n36422,
         n36423, n36424, n36425, n36426, n36427, n36428, n36429, n36430,
         n36431, n36432, n36433, n36434, n36435, n36436, n36437, n36438,
         n36439, n36440, n36441, n36442, n36443, n36444, n36445, n36446,
         n36447, n36448, n36449, n36450, n36451, n36452, n36453, n36454,
         n36455, n36456, n36457, n36458, n36459, n36460, n36461, n36462,
         n36463, n36464, n36465, n36466, n36467, n36468, n36469, n36470,
         n36471, n36472, n36473, n36474, n36475, n36476, n36477, n36478,
         n36479, n36480, n36481, n36482, n36483, n36484, n36485, n36486,
         n36487, n36488, n36489, n36490, n36491, n36492, n36493, n36494,
         n36495, n36496, n36497, n36498, n36499, n36500, n36501, n36502,
         n36503, n36504, n36505, n36506, n36507, n36508, n36509, n36510,
         n36511, n36512, n36513, n36514, n36515, n36516, n36517, n36518,
         n36519, n36520, n36521, n36522, n36523, n36524, n36525, n36526,
         n36527, n36528, n36529, n36530, n36531, n36532, n36533, n36534,
         n36535, n36536, n36537, n36538, n36539, n36540, n36541, n36542,
         n36543, n36544, n36545, n36546, n36547, n36548, n36549, n36550,
         n36551, n36552, n36553, n36554, n36555, n36556, n36557, n36558,
         n36559, n36560, n36561, n36562, n36563, n36564, n36565, n36566,
         n36567, n36568, n36569, n36570, n36571, n36572, n36573, n36574,
         n36575, n36576, n36577, n36578, n36579, n36580, n36581, n36582,
         n36583, n36584, n36585, n36586, n36587, n36588, n36589, n36590,
         n36591, n36592, n36593, n36594, n36595, n36596, n36597, n36598,
         n36599, n36600, n36601, n36602, n36603, n36604, n36605, n36606,
         n36607, n36608, n36609, n36610, n36611, n36612, n36613, n36614,
         n36615, n36616, n36617, n36618, n36619, n36620, n36621, n36622,
         n36623, n36624, n36625, n36626, n36627, n36628, n36629, n36630,
         n36631, n36632, n36633, n36634, n36635, n36636, n36637, n36638,
         n36639, n36640, n36641, n36642, n36643, n36644, n36645, n36646,
         n36647, n36648, n36649, n36650, n36651, n36652, n36653, n36654,
         n36655, n36656, n36657, n36658, n36659, n36660, n36661, n36662,
         n36663, n36664, n36665, n36666, n36667, n36668, n36669, n36670,
         n36671, n36672, n36673, n36674, n36675, n36676, n36677, n36678,
         n36679, n36680, n36681, n36682, n36683, n36684, n36685, n36686,
         n36687, n36688, n36689, n36690, n36691, n36692, n36693, n36694,
         n36695, n36696, n36697, n36698, n36699, n36700, n36701, n36702,
         n36703, n36704, n36705, n36706, n36707, n36708, n36709, n36710,
         n36711, n36712, n36713, n36714, n36715, n36716, n36717, n36718,
         n36719, n36720, n36721, n36722, n36723, n36724, n36725, n36726,
         n36727, n36728, n36729, n36730, n36731, n36732, n36733, n36734,
         n36735, n36736, n36737, n36738, n36739, n36740, n36741, n36742,
         n36743, n36744, n36745, n36746, n36747, n36748, n36749, n36750,
         n36751, n36752, n36753, n36754, n36755, n36756, n36757, n36758,
         n36759, n36760, n36761, n36762, n36763, n36764, n36765, n36766,
         n36767, n36768, n36769, n36770, n36771, n36772, n36773, n36774,
         n36775, n36776, n36777, n36778, n36779, n36780, n36781, n36782,
         n36783, n36784, n36785, n36786, n36787, n36788, n36789, n36790,
         n36791, n36792, n36793, n36794, n36795, n36796, n36797, n36798,
         n36799, n36800, n36801, n36802, n36803, n36804, n36805, n36806,
         n36807, n36808, n36809, n36810, n36811, n36812, n36813, n36814,
         n36815, n36816, n36817, n36818, n36819, n36820, n36821, n36822,
         n36823, n36824, n36825, n36826, n36827, n36828, n36829, n36830,
         n36831, n36832, n36833, n36834, n36835, n36836, n36837, n36838,
         n36839, n36840, n36841, n36842, n36843, n36844, n36845, n36846,
         n36847, n36848, n36849, n36850, n36851, n36852, n36853, n36854,
         n36855, n36856, n36857, n36858, n36859, n36860, n36861, n36862,
         n36863, n36864, n36865, n36866, n36867, n36868, n36869, n36870,
         n36871, n36872, n36873, n36874, n36875, n36876, n36877, n36878,
         n36879, n36880, n36881, n36882, n36883, n36884, n36885, n36886,
         n36887, n36888, n36889, n36890, n36891, n36892, n36893, n36894,
         n36895, n36896, n36897, n36898, n36899, n36900, n36901, n36902,
         n36903, n36904, n36905, n36906, n36907, n36908, n36909, n36910,
         n36911, n36912, n36913, n36914, n36915, n36916, n36917, n36918,
         n36919, n36920, n36921, n36922, n36923, n36924, n36925, n36926,
         n36927, n36928, n36929, n36930, n36931, n36932, n36933, n36934,
         n36935, n36936, n36937, n36938, n36939, n36940, n36941, n36942,
         n36943, n36944, n36945, n36946, n36947, n36948, n36949, n36950,
         n36951, n36952, n36953, n36954, n36955, n36956, n36957, n36958,
         n36959, n36960, n36961, n36962, n36963, n36964, n36965, n36966,
         n36967, n36968, n36969, n36970, n36971, n36972, n36973, n36974,
         n36975, n36976, n36977, n36978, n36979, n36980, n36981, n36982,
         n36983, n36984, n36985, n36986, n36987, n36988, n36989, n36990,
         n36991, n36992, n36993, n36994, n36995, n36996, n36997, n36998,
         n36999, n37000, n37001, n37002, n37003, n37004, n37005, n37006,
         n37007, n37008, n37009, n37010, n37011, n37012, n37013, n37014,
         n37015, n37016, n37017, n37018, n37019, n37020, n37021, n37022,
         n37023, n37024, n37025, n37026, n37027, n37028, n37029, n37030,
         n37031, n37032, n37033, n37034, n37035, n37036, n37037, n37038,
         n37039, n37040, n37041, n37042, n37043, n37044, n37045, n37046,
         n37047, n37048, n37049, n37050, n37051, n37052, n37053, n37054,
         n37055, n37056, n37057, n37058, n37059, n37060, n37061, n37062,
         n37063, n37064, n37065, n37066, n37067, n37068, n37069, n37070,
         n37071, n37072, n37073, n37074, n37075, n37076, n37077, n37078,
         n37079, n37080, n37081, n37082, n37083, n37084, n37085, n37086,
         n37087, n37088, n37089, n37090, n37091, n37092, n37093, n37094,
         n37095, n37096, n37097, n37098, n37099, n37100, n37101, n37102,
         n37103, n37104, n37105, n37106, n37107, n37108, n37109, n37110,
         n37111, n37112, n37113, n37114, n37115, n37116, n37117, n37118,
         n37119, n37120, n37121, n37122, n37123, n37124, n37125, n37126,
         n37127, n37128, n37129, n37130, n37131, n37132, n37133, n37134,
         n37135, n37136, n37137, n37138, n37139, n37140, n37141, n37142,
         n37143, n37144, n37145, n37146, n37147, n37148, n37149, n37150,
         n37151, n37152, n37153, n37154, n37155, n37156, n37157, n37158,
         n37159, n37160, n37161, n37162, n37163, n37164, n37165, n37166,
         n37167, n37168, n37169, n37170, n37171, n37172, n37173, n37174,
         n37175, n37176, n37177, n37178, n37179, n37180, n37181, n37182,
         n37183, n37184, n37185, n37186, n37187, n37188, n37189, n37190,
         n37191, n37192, n37193, n37194, n37195, n37196, n37197, n37198,
         n37199, n37200, n37201, n37202, n37203, n37204, n37205, n37206,
         n37207, n37208, n37209, n37210, n37211, n37212, n37213, n37214,
         n37215, n37216, n37217, n37218, n37219, n37220, n37221, n37222,
         n37223, n37224, n37225, n37226, n37227, n37228, n37229, n37230,
         n37231, n37232, n37233, n37234, n37235, n37236, n37237, n37238,
         n37239, n37240, n37241, n37242, n37243, n37244, n37245, n37246,
         n37247, n37248, n37249, n37250, n37251, n37252, n37253, n37254,
         n37255, n37256, n37257, n37258, n37259, n37260, n37261, n37262,
         n37263, n37264, n37265, n37266, n37267, n37268, n37269, n37270,
         n37271, n37272, n37273, n37274, n37275, n37276, n37277, n37278,
         n37279, n37280, n37281, n37282, n37283, n37284, n37285, n37286,
         n37287, n37288, n37289, n37290, n37291, n37292, n37293, n37294,
         n37295, n37296, n37297, n37298, n37299, n37300, n37301, n37302,
         n37303, n37304, n37305, n37306, n37307, n37308, n37309, n37310,
         n37311, n37312, n37313, n37314, n37315, n37316, n37317, n37318,
         n37319, n37320, n37321, n37322, n37323, n37324, n37325, n37326,
         n37327, n37328, n37329, n37330, n37331, n37332, n37333, n37334,
         n37335, n37336, n37337, n37338, n37339, n37340, n37341, n37342,
         n37343, n37344, n37345, n37346, n37347, n37348, n37349, n37350,
         n37351, n37352, n37353, n37354, n37355, n37356, n37357, n37358,
         n37359, n37360, n37361, n37362, n37363, n37364, n37365, n37366,
         n37367, n37368, n37369, n37370, n37371, n37372, n37373, n37374,
         n37375, n37376, n37377, n37378, n37379, n37380, n37381, n37382,
         n37383, n37384, n37385, n37386, n37387, n37388, n37389, n37390,
         n37391, n37392, n37393, n37394, n37395, n37396, n37397, n37398,
         n37399, n37400, n37401, n37402, n37403, n37404, n37405, n37406,
         n37407, n37408, n37409, n37410, n37411, n37412, n37413, n37414,
         n37415, n37416, n37417, n37418, n37419, n37420, n37421, n37422,
         n37423, n37424, n37425, n37426, n37427, n37428, n37429, n37430,
         n37431, n37432, n37433, n37434, n37435, n37436, n37437, n37438,
         n37439, n37440, n37441, n37442, n37443, n37444, n37445, n37446,
         n37447, n37448, n37449, n37450, n37451, n37452, n37453, n37454,
         n37455, n37456, n37457, n37458, n37459, n37460, n37461, n37462,
         n37463, n37464, n37465, n37466, n37467, n37468, n37469, n37470,
         n37471, n37472, n37473, n37474, n37475, n37476, n37477, n37478,
         n37479, n37480, n37481, n37482, n37483, n37484, n37485, n37486,
         n37487, n37488, n37489, n37490, n37491, n37492, n37493, n37494,
         n37495, n37496, n37497, n37498, n37499, n37500, n37501, n37502,
         n37503, n37504, n37505, n37506, n37507, n37508, n37509, n37510,
         n37511, n37512, n37513, n37514, n37515, n37516, n37517, n37518,
         n37519, n37520, n37521, n37522, n37523, n37524, n37525, n37526,
         n37527, n37528, n37529, n37530, n37531, n37532, n37533, n37534,
         n37535, n37536, n37537, n37538, n37539, n37540, n37541, n37542,
         n37543, n37544, n37545, n37546, n37547, n37548, n37549, n37550,
         n37551, n37552, n37553, n37554, n37555, n37556, n37557, n37558,
         n37559, n37560, n37561, n37562, n37563, n37564, n37565, n37566,
         n37567, n37568, n37569, n37570, n37571, n37572, n37573, n37574,
         n37575, n37576, n37577, n37578, n37579, n37580, n37581, n37582,
         n37583, n37584, n37585, n37586, n37587, n37588, n37589, n37590,
         n37591, n37592, n37593, n37594, n37595, n37596, n37597, n37598,
         n37599, n37600, n37601, n37602, n37603, n37604, n37605, n37606,
         n37607, n37608, n37609, n37610, n37611, n37612, n37613, n37614,
         n37615, n37616, n37617, n37618, n37619, n37620, n37621, n37622,
         n37623, n37624, n37625, n37626, n37627, n37628, n37629, n37630,
         n37631, n37632, n37633, n37634, n37635, n37636, n37637, n37638,
         n37639, n37640, n37641, n37642, n37643, n37644, n37645, n37646,
         n37647, n37648, n37649, n37650, n37651, n37652, n37653, n37654,
         n37655, n37656, n37657, n37658, n37659, n37660, n37661, n37662,
         n37663, n37664, n37665, n37666, n37667, n37668, n37669, n37670,
         n37671, n37672, n37673, n37674, n37675, n37676, n37677, n37678,
         n37679, n37680, n37681, n37682, n37683, n37684, n37685, n37686,
         n37687, n37688, n37689, n37690, n37691, n37692, n37693, n37694,
         n37695, n37696, n37697, n37698, n37699, n37700, n37701, n37702,
         n37703, n37704, n37705, n37706, n37707, n37708, n37709, n37710,
         n37711, n37712, n37713, n37714, n37715, n37716, n37717, n37718,
         n37719, n37720, n37721, n37722, n37723, n37724, n37725, n37726,
         n37727, n37728, n37729, n37730, n37731, n37732, n37733, n37734,
         n37735, n37736, n37737, n37738, n37739, n37740, n37741, n37742,
         n37743, n37744, n37745, n37746, n37747, n37748, n37749, n37750,
         n37751, n37752, n37753, n37754, n37755, n37756, n37757, n37758,
         n37759, n37760, n37761, n37762, n37763, n37764, n37765, n37766,
         n37767, n37768, n37769, n37770, n37771, n37772, n37773, n37774,
         n37775, n37776, n37777, n37778, n37779, n37780, n37781, n37782,
         n37783, n37784, n37785, n37786, n37787, n37788, n37789, n37790,
         n37791, n37792, n37793, n37794, n37795, n37796, n37797, n37798,
         n37799, n37800, n37801, n37802, n37803, n37804, n37805, n37806,
         n37807, n37808, n37809, n37810, n37811, n37812, n37813, n37814,
         n37815, n37816, n37817, n37818, n37819, n37820, n37821, n37822,
         n37823, n37824, n37825, n37826, n37827, n37828, n37829, n37830,
         n37831, n37832, n37833, n37834, n37835, n37836, n37837, n37838,
         n37839, n37840, n37841, n37842, n37843, n37844, n37845, n37846,
         n37847, n37848, n37849, n37850, n37851, n37852, n37853, n37854,
         n37855, n37856, n37857, n37858, n37859, n37860, n37861, n37862,
         n37863, n37864, n37865, n37866, n37867, n37868, n37869, n37870,
         n37871, n37872, n37873, n37874, n37875, n37876, n37877, n37878,
         n37879, n37880, n37881, n37882, n37883, n37884, n37885, n37886,
         n37887, n37888, n37889, n37890, n37891, n37892, n37893, n37894,
         n37895, n37896, n37897, n37898, n37899, n37900, n37901, n37902,
         n37903, n37904, n37905, n37906, n37907, n37908, n37909, n37910,
         n37911, n37912, n37913, n37914, n37915, n37916, n37917, n37918,
         n37919, n37920, n37921, n37922, n37923, n37924, n37925, n37926,
         n37927, n37928, n37929, n37930, n37931, n37932, n37933, n37934,
         n37935, n37936, n37937, n37938, n37939, n37940, n37941, n37942,
         n37943, n37944, n37945, n37946, n37947, n37948, n37949, n37950,
         n37951, n37952, n37953, n37954, n37955, n37956, n37957, n37958,
         n37959, n37960, n37961, n37962, n37963, n37964, n37965, n37966,
         n37967, n37968, n37969, n37970, n37971, n37972, n37973, n37974,
         n37975, n37976, n37977, n37978, n37979, n37980, n37981, n37982,
         n37983, n37984, n37985, n37986, n37987, n37988, n37989, n37990,
         n37991, n37992, n37993, n37994, n37995, n37996, n37997, n37998,
         n37999, n38000, n38001, n38002, n38003, n38004, n38005, n38006,
         n38007, n38008, n38009, n38010, n38011, n38012, n38013, n38014,
         n38015, n38016, n38017, n38018, n38019, n38020, n38021, n38022,
         n38023, n38024, n38025, n38026, n38027, n38028, n38029, n38030,
         n38031, n38032, n38033, n38034, n38035, n38036, n38037, n38038,
         n38039, n38040, n38041, n38042, n38043, n38044, n38045, n38046,
         n38047, n38048, n38049, n38050, n38051, n38052, n38053, n38054,
         n38055, n38056, n38057, n38058, n38059, n38060, n38061, n38062,
         n38063, n38064, n38065, n38066, n38067, n38068, n38069, n38070,
         n38071, n38072, n38073, n38074, n38075, n38076, n38077, n38078,
         n38079, n38080, n38081, n38082, n38083, n38084, n38085, n38086,
         n38087, n38088, n38089, n38090, n38091, n38092, n38093, n38094,
         n38095, n38096, n38097, n38098, n38099, n38100, n38101, n38102,
         n38103, n38104, n38105, n38106, n38107, n38108, n38109, n38110,
         n38111, n38112, n38113, n38114, n38115, n38116, n38117, n38118,
         n38119, n38120, n38121, n38122, n38123, n38124, n38125, n38126,
         n38127, n38128, n38129, n38130, n38131, n38132, n38133, n38134,
         n38135, n38136, n38137, n38138, n38139, n38140, n38141, n38142,
         n38143, n38144, n38145, n38146, n38147, n38148, n38149, n38150,
         n38151, n38152, n38153, n38154, n38155, n38156, n38157, n38158,
         n38159, n38160, n38161, n38162, n38163, n38164, n38165, n38166,
         n38167, n38168, n38169, n38170, n38171, n38172, n38173, n38174,
         n38175, n38176, n38177, n38178, n38179, n38180, n38181, n38182,
         n38183, n38184, n38185, n38186, n38187, n38188, n38189, n38190,
         n38191, n38192, n38193, n38194, n38195, n38196, n38197, n38198,
         n38199, n38200, n38201, n38202, n38203, n38204, n38205, n38206,
         n38207, n38208, n38209, n38210, n38211, n38212, n38213, n38214,
         n38215, n38216, n38217, n38218, n38219, n38220, n38221, n38222,
         n38223, n38224, n38225, n38226, n38227, n38228, n38229, n38230,
         n38231, n38232, n38233, n38234, n38235, n38236, n38237, n38238,
         n38239, n38240, n38241, n38242, n38243, n38244, n38245, n38246,
         n38247, n38248, n38249, n38250, n38251, n38252, n38253, n38254,
         n38255, n38256, n38257, n38258, n38259, n38260, n38261, n38262,
         n38263, n38264, n38265, n38266, n38267, n38268, n38269, n38270,
         n38271, n38272, n38273, n38274, n38275, n38276, n38277, n38278,
         n38279, n38280, n38281, n38282, n38283, n38284, n38285, n38286,
         n38287, n38288, n38289, n38290, n38291, n38292, n38293, n38294,
         n38295, n38296, n38297, n38298, n38299, n38300, n38301, n38302,
         n38303, n38304, n38305, n38306, n38307, n38308, n38309, n38310,
         n38311, n38312, n38313, n38314, n38315, n38316, n38317, n38318,
         n38319, n38320, n38321, n38322, n38323, n38324, n38325, n38326,
         n38327, n38328, n38329, n38330, n38331, n38332, n38333, n38334,
         n38335, n38336, n38337, n38338, n38339, n38340, n38341, n38342,
         n38343, n38344, n38345, n38346, n38347, n38348, n38349, n38350,
         n38351, n38352, n38353, n38354, n38355, n38356, n38357, n38358,
         n38359, n38360, n38361, n38362, n38363, n38364, n38365, n38366,
         n38367, n38368, n38369, n38370, n38371, n38372, n38373, n38374,
         n38375, n38376, n38377, n38378, n38379, n38380, n38381, n38382,
         n38383, n38384, n38385, n38386, n38387, n38388, n38389, n38390,
         n38391, n38392, n38393, n38394, n38395, n38396, n38397, n38398,
         n38399, n38400, n38401, n38402, n38403, n38404, n38405, n38406,
         n38407, n38408, n38409, n38410, n38411, n38412, n38413, n38414,
         n38415, n38416, n38417, n38418, n38419, n38420, n38421, n38422,
         n38423, n38424, n38425, n38426, n38427, n38428, n38429, n38430,
         n38431, n38432, n38433, n38434, n38435, n38436, n38437, n38438,
         n38439, n38440, n38441, n38442, n38443, n38444, n38445, n38446,
         n38447, n38448, n38449, n38450, n38451, n38452, n38453, n38454,
         n38455, n38456, n38457, n38458, n38459, n38460, n38461, n38462,
         n38463, n38464, n38465, n38466, n38467, n38468, n38469, n38470,
         n38471, n38472, n38473, n38474, n38475, n38476, n38477, n38478,
         n38479, n38480, n38481, n38482, n38483, n38484, n38485, n38486,
         n38487, n38488, n38489, n38490, n38491, n38492, n38493, n38494,
         n38495, n38496, n38497, n38498, n38499, n38500, n38501, n38502,
         n38503, n38504, n38505, n38506, n38507, n38508, n38509, n38510,
         n38511, n38512, n38513, n38514, n38515, n38516, n38517, n38518,
         n38519, n38520, n38521, n38522, n38523, n38524, n38525, n38526,
         n38527, n38528, n38529, n38530, n38531, n38532, n38533, n38534,
         n38535, n38536, n38537, n38538, n38539, n38540, n38541, n38542,
         n38543, n38544, n38545, n38546, n38547, n38548, n38549, n38550,
         n38551, n38552, n38553, n38554, n38555, n38556, n38557, n38558,
         n38559, n38560, n38561, n38562, n38563, n38564, n38565, n38566,
         n38567, n38568, n38569, n38570, n38571, n38572, n38573, n38574,
         n38575, n38576, n38577, n38578, n38579, n38580, n38581, n38582,
         n38583, n38584, n38585, n38586, n38587, n38588, n38589, n38590,
         n38591, n38592, n38593, n38594, n38595, n38596, n38597, n38598,
         n38599, n38600, n38601, n38602, n38603, n38604, n38605, n38606,
         n38607, n38608, n38609, n38610, n38611, n38612, n38613, n38614,
         n38615, n38616, n38617, n38618, n38619, n38620, n38621, n38622,
         n38623, n38624, n38625, n38626, n38627, n38628, n38629, n38630,
         n38631, n38632, n38633, n38634, n38635, n38636, n38637, n38638,
         n38639, n38640, n38641, n38642, n38643, n38644, n38645, n38646,
         n38647, n38648, n38649, n38650, n38651, n38652, n38653, n38654,
         n38655, n38656, n38657, n38658, n38659, n38660, n38661, n38662,
         n38663, n38664, n38665, n38666, n38667, n38668, n38669, n38670,
         n38671, n38672, n38673, n38674, n38675, n38676, n38677, n38678,
         n38679, n38680, n38681, n38682, n38683, n38684, n38685, n38686,
         n38687, n38688, n38689, n38690, n38691, n38692, n38693, n38694,
         n38695, n38696, n38697, n38698, n38699, n38700, n38701, n38702,
         n38703, n38704, n38705, n38706, n38707, n38708, n38709, n38710,
         n38711, n38712, n38713, n38714, n38715, n38716, n38717, n38718,
         n38719, n38720, n38721, n38722, n38723, n38724, n38725, n38726,
         n38727, n38728, n38729, n38730, n38731, n38732, n38733, n38734,
         n38735, n38736, n38737, n38738, n38739, n38740, n38741, n38742,
         n38743, n38744, n38745, n38746, n38747, n38748, n38749, n38750,
         n38751, n38752, n38753, n38754, n38755, n38756, n38757, n38758,
         n38759, n38760, n38761, n38762, n38763, n38764, n38765, n38766,
         n38767, n38768, n38769, n38770, n38771, n38772, n38773, n38774,
         n38775, n38776, n38777, n38778, n38779, n38780, n38781, n38782,
         n38783, n38784, n38785, n38786, n38787, n38788, n38789, n38790,
         n38791, n38792, n38793, n38794, n38795, n38796, n38797, n38798,
         n38799, n38800, n38801, n38802, n38803, n38804, n38805, n38806,
         n38807, n38808, n38809, n38810, n38811, n38812, n38813, n38814,
         n38815, n38816, n38817, n38818, n38819, n38820, n38821, n38822,
         n38823, n38824, n38825, n38826, n38827, n38828, n38829, n38830,
         n38831, n38832, n38833, n38834, n38835, n38836, n38837, n38838,
         n38839, n38840, n38841, n38842, n38843, n38844, n38845, n38846,
         n38847, n38848, n38849, n38850, n38851, n38852, n38853, n38854,
         n38855, n38856, n38857, n38858, n38859, n38860, n38861, n38862,
         n38863, n38864, n38865, n38866, n38867, n38868, n38869, n38870,
         n38871, n38872, n38873, n38874, n38875, n38876, n38877, n38878,
         n38879, n38880, n38881, n38882, n38883, n38884, n38885, n38886,
         n38887, n38888, n38889, n38890, n38891, n38892, n38893, n38894,
         n38895, n38896, n38897, n38898, n38899, n38900, n38901, n38902,
         n38903, n38904, n38905, n38906, n38907, n38908, n38909, n38910,
         n38911, n38912, n38913, n38914, n38915, n38916, n38917, n38918,
         n38919, n38920, n38921, n38922, n38923, n38924, n38925, n38926,
         n38927, n38928, n38929, n38930, n38931, n38932, n38933, n38934,
         n38935, n38936, n38937, n38938, n38939, n38940, n38941, n38942,
         n38943, n38944, n38945, n38946, n38947, n38948, n38949, n38950,
         n38951, n38952, n38953, n38954, n38955, n38956, n38957, n38958,
         n38959, n38960, n38961, n38962, n38963, n38964, n38965, n38966,
         n38967, n38968, n38969, n38970, n38971, n38972, n38973, n38974,
         n38975, n38976, n38977, n38978, n38979, n38980, n38981, n38982,
         n38983, n38984, n38985, n38986, n38987, n38988, n38989, n38990,
         n38991, n38992, n38993, n38994, n38995, n38996, n38997, n38998,
         n38999, n39000, n39001, n39002, n39003, n39004, n39005, n39006,
         n39007, n39008, n39009, n39010, n39011, n39012, n39013, n39014,
         n39015, n39016, n39017, n39018, n39019, n39020, n39021, n39022,
         n39023, n39024, n39025, n39026, n39027, n39028, n39029, n39030,
         n39031, n39032, n39033, n39034, n39035, n39036, n39037, n39038,
         n39039, n39040, n39041, n39042, n39043, n39044, n39045, n39046,
         n39047, n39048, n39049, n39050, n39051, n39052, n39053, n39054,
         n39055, n39056, n39057, n39058, n39059, n39060, n39061, n39062,
         n39063, n39064, n39065, n39066, n39067, n39068, n39069, n39070,
         n39071, n39072, n39073, n39074, n39075, n39076, n39077, n39078,
         n39079, n39080, n39081, n39082, n39083, n39084, n39085, n39086,
         n39087, n39088, n39089, n39090, n39091, n39092, n39093, n39094,
         n39095, n39096, n39097, n39098, n39099, n39100, n39101, n39102,
         n39103, n39104, n39105, n39106, n39107, n39108, n39109, n39110,
         n39111, n39112, n39113, n39114, n39115, n39116, n39117, n39118,
         n39119, n39120, n39121, n39122, n39123, n39124, n39125, n39126,
         n39127, n39128, n39129, n39130, n39131, n39132, n39133, n39134,
         n39135, n39136, n39137, n39138, n39139, n39140, n39141, n39142,
         n39143, n39144, n39145, n39146, n39147, n39148, n39149, n39150,
         n39151, n39152, n39153, n39154, n39155, n39156, n39157, n39158,
         n39159, n39160, n39161, n39162, n39163, n39164, n39165, n39166,
         n39167, n39168, n39169, n39170, n39171, n39172, n39173, n39174,
         n39175, n39176, n39177, n39178, n39179, n39180, n39181, n39182,
         n39183, n39184, n39185, n39186, n39187, n39188, n39189, n39190,
         n39191, n39192, n39193, n39194, n39195, n39196, n39197, n39198,
         n39199, n39200, n39201, n39202, n39203, n39204, n39205, n39206,
         n39207, n39208, n39209, n39210, n39211, n39212, n39213, n39214,
         n39215, n39216, n39217, n39218, n39219, n39220, n39221, n39222,
         n39223, n39224, n39225, n39226, n39227, n39228, n39229, n39230,
         n39231, n39232, n39233, n39234, n39235, n39236, n39237, n39238,
         n39239, n39240, n39241, n39242, n39243, n39244, n39245, n39246,
         n39247, n39248, n39249, n39250, n39251, n39252, n39253, n39254,
         n39255, n39256, n39257, n39258, n39259, n39260, n39261, n39262,
         n39263, n39264, n39265, n39266, n39267, n39268, n39269, n39270,
         n39271, n39272, n39273, n39274, n39275, n39276, n39277, n39278,
         n39279, n39280, n39281, n39282, n39283, n39284, n39285, n39286,
         n39287, n39288, n39289, n39290, n39291, n39292, n39293, n39294,
         n39295, n39296, n39297, n39298, n39299, n39300, n39301, n39302,
         n39303, n39304, n39305, n39306, n39307, n39308, n39309, n39310,
         n39311, n39312, n39313, n39314, n39315, n39316, n39317, n39318,
         n39319, n39320, n39321, n39322, n39323, n39324, n39325, n39326,
         n39327, n39328, n39329, n39330, n39331, n39332, n39333, n39334,
         n39335, n39336, n39337, n39338, n39339, n39340, n39341, n39342,
         n39343, n39344, n39345, n39346, n39347, n39348, n39349, n39350,
         n39351, n39352, n39353, n39354, n39355, n39356, n39357, n39358,
         n39359, n39360, n39361, n39362, n39363, n39364, n39365, n39366,
         n39367, n39368, n39369, n39370, n39371, n39372, n39373, n39374,
         n39375, n39376, n39377, n39378, n39379, n39380, n39381, n39382,
         n39383, n39384, n39385, n39386, n39387, n39388, n39389, n39390,
         n39391, n39392, n39393, n39394, n39395, n39396, n39397, n39398,
         n39399, n39400, n39401, n39402, n39403, n39404, n39405, n39406,
         n39407, n39408, n39409, n39410, n39411, n39412, n39413, n39414,
         n39415, n39416, n39417, n39418, n39419, n39420, n39421, n39422,
         n39423, n39424, n39425, n39426, n39427, n39428, n39429, n39430,
         n39431, n39432, n39433, n39434, n39435, n39436, n39437, n39438,
         n39439, n39440, n39441, n39442, n39443, n39444, n39445, n39446,
         n39447, n39448, n39449, n39450, n39451, n39452, n39453, n39454,
         n39455, n39456, n39457, n39458, n39459, n39460, n39461, n39462,
         n39463, n39464, n39465, n39466, n39467, n39468, n39469, n39470,
         n39471, n39472, n39473, n39474, n39475, n39476, n39477, n39478,
         n39479, n39480, n39481, n39482, n39483, n39484, n39485, n39486,
         n39487, n39488, n39489, n39490, n39491, n39492, n39493, n39494,
         n39495, n39496, n39497, n39498, n39499, n39500, n39501, n39502,
         n39503, n39504, n39505, n39506, n39507, n39508, n39509, n39510,
         n39511, n39512, n39513, n39514, n39515, n39516, n39517, n39518,
         n39519, n39520, n39521, n39522, n39523, n39524, n39525, n39526,
         n39527, n39528, n39529, n39530, n39531, n39532, n39533, n39534,
         n39535, n39536, n39537, n39538, n39539, n39540, n39541, n39542,
         n39543, n39544, n39545, n39546, n39547, n39548, n39549, n39550,
         n39551, n39552, n39553, n39554, n39555, n39556, n39557, n39558,
         n39559, n39560, n39561, n39562, n39563, n39564, n39565, n39566,
         n39567, n39568, n39569, n39570, n39571, n39572, n39573, n39574,
         n39575, n39576, n39577, n39578, n39579, n39580, n39581, n39582,
         n39583, n39584, n39585, n39586, n39587, n39588, n39589, n39590,
         n39591, n39592, n39593, n39594, n39595, n39596, n39597, n39598,
         n39599, n39600, n39601, n39602, n39603, n39604, n39605, n39606,
         n39607, n39608, n39609, n39610, n39611, n39612, n39613, n39614,
         n39615, n39616, n39617, n39618, n39619, n39620, n39621, n39622,
         n39623, n39624, n39625, n39626, n39627, n39628, n39629, n39630,
         n39631, n39632, n39633, n39634, n39635, n39636, n39637, n39638,
         n39639, n39640, n39641, n39642, n39643, n39644, n39645, n39646,
         n39647, n39648, n39649, n39650, n39651, n39652, n39653, n39654,
         n39655, n39656, n39657, n39658, n39659, n39660, n39661, n39662,
         n39663, n39664, n39665, n39666, n39667, n39668, n39669, n39670,
         n39671, n39672, n39673, n39674, n39675, n39676, n39677, n39678,
         n39679, n39680, n39681, n39682, n39683, n39684, n39685, n39686,
         n39687, n39688, n39689, n39690, n39691, n39692, n39693, n39694,
         n39695, n39696, n39697, n39698, n39699, n39700, n39701, n39702,
         n39703, n39704, n39705, n39706, n39707, n39708, n39709, n39710,
         n39711, n39712, n39713, n39714, n39715, n39716, n39717, n39718,
         n39719, n39720, n39721, n39722, n39723, n39724, n39725, n39726,
         n39727, n39728, n39729, n39730, n39731, n39732, n39733, n39734,
         n39735, n39736, n39737, n39738, n39739, n39740, n39741, n39742,
         n39743, n39744, n39745, n39746, n39747, n39748, n39749, n39750,
         n39751, n39752, n39753, n39754, n39755, n39756, n39757, n39758,
         n39759, n39760, n39761, n39762, n39763, n39764, n39765, n39766,
         n39767, n39768, n39769, n39770, n39771, n39772, n39773, n39774,
         n39775, n39776, n39777, n39778, n39779, n39780, n39781, n39782,
         n39783, n39784, n39785, n39786, n39787, n39788, n39789, n39790,
         n39791, n39792, n39793, n39794, n39795, n39796, n39797, n39798,
         n39799, n39800, n39801, n39802, n39803, n39804, n39805, n39806,
         n39807, n39808, n39809, n39810, n39811, n39812, n39813, n39814,
         n39815, n39816, n39817, n39818, n39819, n39820, n39821, n39822,
         n39823, n39824, n39825, n39826, n39827, n39828, n39829, n39830,
         n39831, n39832, n39833, n39834, n39835, n39836, n39837, n39838,
         n39839, n39840, n39841, n39842, n39843, n39844, n39845, n39846,
         n39847, n39848, n39849, n39850, n39851, n39852, n39853, n39854,
         n39855, n39856, n39857, n39858, n39859, n39860, n39861, n39862,
         n39863, n39864, n39865, n39866, n39867, n39868, n39869, n39870,
         n39871, n39872, n39873, n39874, n39875, n39876, n39877, n39878,
         n39879, n39880, n39881, n39882, n39883, n39884, n39885, n39886,
         n39887, n39888, n39889, n39890, n39891, n39892, n39893, n39894,
         n39895, n39896, n39897, n39898, n39899, n39900, n39901, n39902,
         n39903, n39904, n39905, n39906, n39907, n39908, n39909, n39910,
         n39911, n39912, n39913, n39914, n39915, n39916, n39917, n39918,
         n39919, n39920, n39921, n39922, n39923, n39924, n39925, n39926,
         n39927, n39928, n39929, n39930, n39931, n39932, n39933, n39934,
         n39935, n39936, n39937, n39938, n39939, n39940, n39941, n39942,
         n39943, n39944, n39945, n39946, n39947, n39948, n39949, n39950,
         n39951, n39952, n39953, n39954, n39955, n39956, n39957, n39958,
         n39959, n39960, n39961, n39962, n39963, n39964, n39965, n39966,
         n39967, n39968, n39969, n39970, n39971, n39972, n39973, n39974,
         n39975, n39976, n39977, n39978, n39979, n39980, n39981, n39982,
         n39983, n39984, n39985, n39986, n39987, n39988, n39989, n39990,
         n39991, n39992, n39993, n39994, n39995, n39996, n39997, n39998,
         n39999, n40000, n40001, n40002, n40003, n40004, n40005, n40006,
         n40007, n40008, n40009, n40010, n40011, n40012, n40013, n40014,
         n40015, n40016, n40017, n40018, n40019, n40020, n40021, n40022,
         n40023, n40024, n40025, n40026, n40027, n40028, n40029, n40030,
         n40031, n40032, n40033, n40034, n40035, n40036, n40037, n40038,
         n40039, n40040, n40041, n40042, n40043, n40044, n40045, n40046,
         n40047, n40048, n40049, n40050, n40051, n40052, n40053, n40054,
         n40055, n40056, n40057, n40058, n40059, n40060, n40061, n40062,
         n40063, n40064, n40065, n40066, n40067, n40068, n40069, n40070,
         n40071, n40072, n40073, n40074, n40075, n40076, n40077, n40078,
         n40079, n40080, n40081, n40082, n40083, n40084, n40085, n40086,
         n40087, n40088, n40089, n40090, n40091, n40092, n40093, n40094,
         n40095, n40096, n40097, n40098, n40099, n40100, n40101, n40102,
         n40103, n40104, n40105, n40106, n40107, n40108, n40109, n40110,
         n40111, n40112, n40113, n40114, n40115, n40116, n40117, n40118,
         n40119, n40120, n40121, n40122, n40123, n40124, n40125, n40126,
         n40127, n40128, n40129, n40130, n40131, n40132, n40133, n40134,
         n40135, n40136, n40137, n40138, n40139, n40140, n40141, n40142,
         n40143, n40144, n40145, n40146, n40147, n40148, n40149, n40150,
         n40151, n40152, n40153, n40154, n40155, n40156, n40157, n40158,
         n40159, n40160, n40161, n40162, n40163, n40164, n40165, n40166,
         n40167, n40168, n40169, n40170, n40171, n40172, n40173, n40174,
         n40175, n40176, n40177, n40178, n40179, n40180, n40181, n40182,
         n40183, n40184, n40185, n40186, n40187, n40188, n40189, n40190,
         n40191, n40192, n40193, n40194, n40195, n40196, n40197, n40198,
         n40199, n40200, n40201, n40202, n40203, n40204, n40205, n40206,
         n40207, n40208, n40209, n40210, n40211, n40212, n40213, n40214,
         n40215, n40216, n40217, n40218, n40219, n40220, n40221, n40222,
         n40223, n40224, n40225, n40226, n40227, n40228, n40229, n40230,
         n40231, n40232, n40233, n40234, n40235, n40236, n40237, n40238,
         n40239, n40240, n40241, n40242, n40243, n40244, n40245, n40246,
         n40247, n40248, n40249, n40250, n40251, n40252, n40253, n40254,
         n40255, n40256, n40257, n40258, n40259, n40260, n40261, n40262,
         n40263, n40264, n40265, n40266, n40267, n40268, n40269, n40270,
         n40271, n40272, n40273, n40274, n40275, n40276, n40277, n40278,
         n40279, n40280, n40281, n40282, n40283, n40284, n40285, n40286,
         n40287, n40288, n40289, n40290, n40291, n40292, n40293, n40294,
         n40295, n40296, n40297, n40298, n40299, n40300, n40301, n40302,
         n40303, n40304, n40305, n40306, n40307, n40308, n40309, n40310,
         n40311, n40312, n40313, n40314, n40315, n40316, n40317, n40318,
         n40319, n40320, n40321, n40322, n40323, n40324, n40325, n40326,
         n40327, n40328, n40329, n40330, n40331, n40332, n40333, n40334,
         n40335, n40336, n40337, n40338, n40339, n40340, n40341, n40342,
         n40343, n40344, n40345, n40346, n40347, n40348, n40349, n40350,
         n40351, n40352, n40353, n40354, n40355, n40356, n40357, n40358,
         n40359, n40360, n40361, n40362, n40363, n40364, n40365, n40366,
         n40367, n40368, n40369, n40370, n40371, n40372, n40373, n40374,
         n40375, n40376, n40377, n40378, n40379, n40380, n40381, n40382,
         n40383, n40384, n40385, n40386, n40387, n40388, n40389, n40390,
         n40391, n40392, n40393, n40394, n40395, n40396, n40397, n40398,
         n40399, n40400, n40401, n40402, n40403, n40404, n40405, n40406,
         n40407, n40408, n40409, n40410, n40411, n40412, n40413, n40414,
         n40415, n40416, n40417, n40418, n40419, n40420, n40421, n40422,
         n40423, n40424, n40425, n40426, n40427, n40428, n40429, n40430,
         n40431, n40432, n40433, n40434, n40435, n40436, n40437, n40438,
         n40439, n40440, n40441, n40442, n40443, n40444, n40445, n40446,
         n40447, n40448, n40449, n40450, n40451, n40452, n40453, n40454,
         n40455, n40456, n40457, n40458, n40459, n40460, n40461, n40462,
         n40463, n40464, n40465, n40466, n40467, n40468, n40469, n40470,
         n40471, n40472, n40473, n40474, n40475, n40476, n40477, n40478,
         n40479, n40480, n40481, n40482, n40483, n40484, n40485, n40486,
         n40487, n40488, n40489, n40490, n40491, n40492, n40493, n40494,
         n40495, n40496, n40497, n40498, n40499, n40500, n40501, n40502,
         n40503, n40504, n40505, n40506, n40507, n40508, n40509, n40510,
         n40511, n40512, n40513, n40514, n40515, n40516, n40517, n40518,
         n40519, n40520, n40521, n40522, n40523, n40524, n40525, n40526,
         n40527, n40528, n40529, n40530, n40531, n40532, n40533, n40534,
         n40535, n40536, n40537, n40538, n40539, n40540, n40541, n40542,
         n40543, n40544, n40545, n40546, n40547, n40548, n40549, n40550,
         n40551, n40552, n40553, n40554, n40555, n40556, n40557, n40558,
         n40559, n40560, n40561, n40562, n40563, n40564, n40565, n40566,
         n40567, n40568, n40569, n40570, n40571, n40572, n40573, n40574,
         n40575, n40576, n40577, n40578, n40579, n40580, n40581, n40582,
         n40583, n40584, n40585, n40586, n40587, n40588, n40589, n40590,
         n40591, n40592, n40593, n40594, n40595, n40596, n40597, n40598,
         n40599, n40600, n40601, n40602, n40603, n40604, n40605, n40606,
         n40607, n40608, n40609, n40610, n40611, n40612, n40613, n40614,
         n40615, n40616, n40617, n40618, n40619, n40620, n40621, n40622,
         n40623, n40624, n40625, n40626, n40627, n40628, n40629, n40630,
         n40631, n40632, n40633, n40634, n40635, n40636, n40637, n40638,
         n40639, n40640, n40641, n40642, n40643, n40644, n40645, n40646,
         n40647, n40648, n40649, n40650, n40651, n40652, n40653, n40654,
         n40655, n40656, n40657, n40658, n40659, n40660, n40661, n40662,
         n40663, n40664, n40665, n40666, n40667, n40668, n40669, n40670,
         n40671, n40672, n40673, n40674, n40675, n40676, n40677, n40678,
         n40679, n40680, n40681, n40682, n40683, n40684, n40685, n40686,
         n40687, n40688, n40689, n40690, n40691, n40692, n40693, n40694,
         n40695, n40696, n40697, n40698, n40699, n40700, n40701, n40702,
         n40703, n40704, n40705, n40706, n40707, n40708, n40709, n40710,
         n40711, n40712, n40713, n40714, n40715, n40716, n40717, n40718,
         n40719, n40720, n40721, n40722, n40723, n40724, n40725, n40726,
         n40727, n40728, n40729, n40730, n40731, n40732, n40733, n40734,
         n40735, n40736, n40737, n40738, n40739, n40740, n40741, n40742,
         n40743, n40744, n40745, n40746, n40747, n40748, n40749, n40750,
         n40751, n40752, n40753, n40754, n40755, n40756, n40757, n40758,
         n40759, n40760, n40761, n40762, n40763, n40764, n40765, n40766,
         n40767, n40768, n40769, n40770, n40771, n40772, n40773, n40774,
         n40775, n40776, n40777, n40778, n40779, n40780, n40781, n40782,
         n40783, n40784, n40785, n40786, n40787, n40788, n40789, n40790,
         n40791, n40792, n40793, n40794, n40795, n40796, n40797, n40798,
         n40799, n40800, n40801, n40802, n40803, n40804, n40805, n40806,
         n40807, n40808, n40809, n40810, n40811, n40812, n40813, n40814,
         n40815, n40816, n40817, n40818, n40819, n40820, n40821, n40822,
         n40823, n40824, n40825, n40826, n40827, n40828, n40829, n40830,
         n40831, n40832, n40833, n40834, n40835, n40836, n40837, n40838,
         n40839, n40840, n40841, n40842, n40843, n40844, n40845, n40846,
         n40847, n40848, n40849, n40850, n40851, n40852, n40853, n40854,
         n40855, n40856, n40857, n40858, n40859, n40860, n40861, n40862,
         n40863, n40864, n40865, n40866, n40867, n40868, n40869, n40870,
         n40871, n40872, n40873, n40874, n40875, n40876, n40877, n40878,
         n40879, n40880, n40881, n40882, n40883, n40884, n40885, n40886,
         n40887, n40888, n40889, n40890, n40891, n40892, n40893, n40894,
         n40895, n40896, n40897, n40898, n40899, n40900, n40901, n40902,
         n40903, n40904, n40905, n40906, n40907, n40908, n40909, n40910,
         n40911, n40912, n40913, n40914, n40915, n40916, n40917, n40918,
         n40919, n40920, n40921, n40922, n40923, n40924, n40925, n40926,
         n40927, n40928, n40929, n40930, n40931, n40932, n40933, n40934,
         n40935, n40936, n40937, n40938, n40939, n40940, n40941, n40942,
         n40943, n40944, n40945, n40946, n40947, n40948, n40949, n40950,
         n40951, n40952, n40953, n40954, n40955, n40956, n40957, n40958,
         n40959, n40960, n40961, n40962, n40963, n40964, n40965, n40966,
         n40967, n40968, n40969, n40970, n40971, n40972, n40973, n40974,
         n40975, n40976, n40977, n40978, n40979, n40980, n40981, n40982,
         n40983, n40984, n40985, n40986, n40987, n40988, n40989, n40990,
         n40991, n40992, n40993, n40994, n40995, n40996, n40997, n40998,
         n40999, n41000;
  wire   [31:0] Data_in;
  wire   [5:0] opcode_i;
  wire   [4:0] \u_DataPath/regfile_addr_out_towb_i ;
  wire   [31:0] \u_DataPath/from_alu_data_out_i ;
  wire   [31:0] \u_DataPath/from_mem_data_out_i ;
  wire   [2:0] \u_DataPath/cw_towb_i ;
  wire   [4:0] \u_DataPath/RFaddr_out_memwb_i ;
  wire   [31:0] \u_DataPath/dataOut_exe_i ;
  wire   [2:0] \u_DataPath/cw_memwb_i ;
  wire   [31:0] \u_DataPath/mem_writedata_out_i ;
  wire   [10:0] \u_DataPath/cw_tomem_i ;
  wire   [10:0] \u_DataPath/cw_exmem_i ;
  wire   [4:0] \u_DataPath/rs_ex_i ;
  wire   [31:0] \u_DataPath/data_read_ex_2_i ;
  wire   [31:0] \u_DataPath/data_read_ex_1_i ;
  wire   [31:0] \u_DataPath/pc_4_to_ex_i ;
  wire   [21:0] \u_DataPath/cw_to_ex_i ;
  wire   [31:0] \u_DataPath/immediate_ext_dec_i ;
  wire   [31:0] \u_DataPath/pc4_to_idexreg_i ;
  wire   [31:0] \u_DataPath/jaddr_i ;
  wire   [4:0] \u_DataPath/idex_rt_i ;
  wire   [31:0] \u_DataPath/pc_4_i ;
  wire   [31:0] \u_DataPath/branch_target_i ;
  wire   [31:0] \u_DataPath/jump_address_i ;
  wire   [1:0] \u_DataPath/u_decode_unit/hdu_0/current_state ;
  wire   [31:0] \u_DataPath/u_execute/psw_status_i ;
  wire   [31:0] \u_DataPath/u_execute/A_inALU_i ;
  wire   [31:0] \u_DataPath/u_execute/link_value_i ;
  wire   [31:0] addr_to_iram;
  assign Address_toRAM[30] = 1'b0;
  assign Address_toRAM[31] = 1'b0;
  assign addr_to_iram[30] = 1'b0;
  assign addr_to_iram[31] = 1'b0;
  assign addr_to_iram[0] = n17639;
  assign addr_to_iram[3] = n18093;
  assign addr_to_iram[2] = n18094;
  assign addr_to_iram[4] = n18095;
  assign addr_to_iram[5] = n18096;
  assign addr_to_iram[7] = n18097;
  assign addr_to_iram[6] = n18098;
  assign addr_to_iram[9] = n18099;
  assign addr_to_iram[8] = n18100;
  assign addr_to_iram[11] = n18101;
  assign addr_to_iram[10] = n18102;
  assign addr_to_iram[13] = n18103;
  assign addr_to_iram[12] = n18104;
  assign addr_to_iram[15] = n18105;
  assign addr_to_iram[14] = n18106;
  assign addr_to_iram[17] = n18107;
  assign addr_to_iram[16] = n18108;
  assign addr_to_iram[19] = n18109;
  assign addr_to_iram[18] = n18110;
  assign addr_to_iram[21] = n18111;
  assign addr_to_iram[20] = n18112;
  assign addr_to_iram[23] = n18113;
  assign addr_to_iram[22] = n18114;
  assign addr_to_iram[25] = n18115;
  assign addr_to_iram[24] = n18116;
  assign addr_to_iram[27] = n18117;
  assign addr_to_iram[26] = n18118;
  assign addr_to_iram[28] = n18119;
  assign addr_to_iram[29] = n18120;
  assign addr_to_iram[1] = n18156;
  assign Address_toRAM[16] = n29562;
  assign Address_toRAM[14] = n29563;
  assign Address_toRAM[15] = n29564;
  assign Address_toRAM[13] = n29565;
  assign Address_toRAM[11] = n29566;
  assign Address_toRAM[10] = n29567;
  assign Address_toRAM[9] = n29568;
  assign Address_toRAM[8] = n29569;
  assign Address_toRAM[7] = n29570;
  assign Address_toRAM[4] = n29571;
  assign Address_toRAM[3] = n29572;
  assign Address_toRAM[5] = n29573;
  assign Address_toRAM[6] = n29574;
  assign Address_toRAM[2] = n29575;
  assign Address_toRAM[1] = n29576;
  assign Data_in[28] = n29577;
  assign Data_in[31] = n29578;
  assign Data_in[27] = n29579;
  assign Data_in[23] = n29580;
  assign Data_in[24] = n29581;
  assign Data_in[25] = n29582;
  assign Data_in[26] = n29583;
  assign Address_toRAM[17] = n29584;
  assign Data_in[30] = n29585;
  assign Data_in[29] = n29586;
  assign nibble[0] = n29587;
  assign nibble[1] = n29588;
  assign write_op = n29589;
  assign Data_in[0] = n29590;
  assign Data_in[3] = n29591;
  assign Data_in[4] = n29592;
  assign Data_in[1] = n29593;
  assign Data_in[2] = n29594;
  assign Data_in[5] = n29595;
  assign Data_in[6] = n29596;
  assign read_op = n29597;
  assign Address_toRAM[12] = n29598;
  assign Data_in[7] = n29599;
  assign Address_toRAM[18] = n29600;
  assign Address_toRAM[19] = n29654;
  assign Data_in[16] = n29656;
  assign Data_in[17] = n29658;
  assign Data_in[18] = n29660;
  assign Data_in[19] = n29662;
  assign Data_in[20] = n29664;
  assign Data_in[21] = n29666;
  assign Data_in[22] = n29668;
  assign Data_in[11] = n29670;
  assign Data_in[15] = n29672;
  assign Address_toRAM[0] = n29674;
  assign Data_in[9] = n29676;
  assign Data_in[12] = n29678;
  assign Data_in[13] = n29680;
  assign Data_in[14] = n29682;
  assign Data_in[8] = n29684;
  assign Data_in[10] = n29686;
  assign Address_toRAM[20] = n29688;
  assign write_byte = n29690;

  HS65_LH_MUX21X4 U1 ( .D0(n38707), .D1(\u_DataPath/u_ifidreg/N52 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/jaddr_i [16]) );
  HS65_LH_MUX21X4 U2 ( .D0(n17692), .D1(\u_DataPath/u_ifidreg/N67 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(opcode_i[5]) );
  HS65_LH_MUX21X4 U3 ( .D0(n40159), .D1(\u_DataPath/u_ifidreg/N66 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(opcode_i[4]) );
  HS65_LH_MUX21X4 U4 ( .D0(n36976), .D1(\u_DataPath/u_ifidreg/N65 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(opcode_i[3]) );
  HS65_LH_MUX21X4 U5 ( .D0(n17642), .D1(\u_DataPath/u_ifidreg/N64 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(opcode_i[2]) );
  HS65_LH_MUX21X4 U6 ( .D0(n17630), .D1(\u_DataPath/u_ifidreg/N63 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(opcode_i[1]) );
  HS65_LH_MUX21X4 U7 ( .D0(n29702), .D1(\u_DataPath/u_ifidreg/N62 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(opcode_i[0]) );
  HS65_LH_MUX21X4 U8 ( .D0(n38702), .D1(\u_DataPath/u_ifidreg/N61 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/jaddr_i [25]) );
  HS65_LH_MUX21X4 U9 ( .D0(n38717), .D1(\u_DataPath/u_ifidreg/N60 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/jaddr_i [24]) );
  HS65_LH_MUX21X4 U10 ( .D0(n38714), .D1(\u_DataPath/u_ifidreg/N59 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/jaddr_i [23]) );
  HS65_LH_MUX21X4 U11 ( .D0(n38711), .D1(\u_DataPath/u_ifidreg/N58 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/jaddr_i [22]) );
  HS65_LH_MUX21X4 U12 ( .D0(n17701), .D1(\u_DataPath/u_ifidreg/N57 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/jaddr_i [21]) );
  HS65_LH_MUX21X4 U13 ( .D0(n38699), .D1(\u_DataPath/u_ifidreg/N56 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/jaddr_i [20]) );
  HS65_LH_MUX21X4 U14 ( .D0(n38720), .D1(\u_DataPath/u_ifidreg/N55 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/jaddr_i [19]) );
  HS65_LH_MUX21X4 U15 ( .D0(n38703), .D1(\u_DataPath/u_ifidreg/N54 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/jaddr_i [18]) );
  HS65_LH_MUX21X4 U16 ( .D0(n38706), .D1(\u_DataPath/u_ifidreg/N53 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/jaddr_i [17]) );
  HS65_LH_MUX21X4 U17 ( .D0(n17649), .D1(\u_DataPath/u_ifidreg/N35 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/pc4_to_idexreg_i [31]) );
  HS65_LH_MUX21X4 U18 ( .D0(n17652), .D1(\u_DataPath/u_ifidreg/N34 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/pc4_to_idexreg_i [30]) );
  HS65_LH_MUX21X4 U19 ( .D0(n17653), .D1(\u_DataPath/u_ifidreg/N33 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/pc4_to_idexreg_i [29]) );
  HS65_LH_MUX21X4 U20 ( .D0(n17654), .D1(\u_DataPath/u_ifidreg/N32 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/pc4_to_idexreg_i [28]) );
  HS65_LH_MUX21X4 U21 ( .D0(n17655), .D1(\u_DataPath/u_ifidreg/N31 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/pc4_to_idexreg_i [27]) );
  HS65_LH_MUX21X4 U22 ( .D0(n17711), .D1(\u_DataPath/u_ifidreg/N30 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/pc4_to_idexreg_i [26]) );
  HS65_LH_MUX21X4 U23 ( .D0(n17712), .D1(\u_DataPath/u_ifidreg/N29 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/pc4_to_idexreg_i [25]) );
  HS65_LH_MUX21X4 U24 ( .D0(n17713), .D1(\u_DataPath/u_ifidreg/N28 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/pc4_to_idexreg_i [24]) );
  HS65_LH_MUX21X4 U25 ( .D0(n17715), .D1(\u_DataPath/u_ifidreg/N27 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/pc4_to_idexreg_i [23]) );
  HS65_LH_MUX21X4 U26 ( .D0(n17717), .D1(\u_DataPath/u_ifidreg/N26 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/pc4_to_idexreg_i [22]) );
  HS65_LH_MUX21X4 U27 ( .D0(n17719), .D1(\u_DataPath/u_ifidreg/N25 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/pc4_to_idexreg_i [21]) );
  HS65_LH_MUX21X4 U28 ( .D0(n17721), .D1(\u_DataPath/u_ifidreg/N24 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/pc4_to_idexreg_i [20]) );
  HS65_LH_MUX21X4 U29 ( .D0(n17723), .D1(\u_DataPath/u_ifidreg/N23 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/pc4_to_idexreg_i [19]) );
  HS65_LH_MUX21X4 U30 ( .D0(n17657), .D1(\u_DataPath/u_ifidreg/N22 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/pc4_to_idexreg_i [18]) );
  HS65_LH_MUX21X4 U31 ( .D0(n17659), .D1(\u_DataPath/u_ifidreg/N21 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/pc4_to_idexreg_i [17]) );
  HS65_LH_MUX21X4 U32 ( .D0(n17660), .D1(\u_DataPath/u_ifidreg/N20 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/pc4_to_idexreg_i [16]) );
  HS65_LH_MUX21X4 U33 ( .D0(n17663), .D1(\u_DataPath/u_ifidreg/N19 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/pc4_to_idexreg_i [15]) );
  HS65_LH_MUX21X4 U34 ( .D0(n17664), .D1(\u_DataPath/u_ifidreg/N18 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/pc4_to_idexreg_i [14]) );
  HS65_LH_MUX21X4 U35 ( .D0(n17667), .D1(\u_DataPath/u_ifidreg/N17 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/pc4_to_idexreg_i [13]) );
  HS65_LH_MUX21X4 U36 ( .D0(n17668), .D1(\u_DataPath/u_ifidreg/N16 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/pc4_to_idexreg_i [12]) );
  HS65_LH_MUX21X4 U37 ( .D0(n17671), .D1(\u_DataPath/u_ifidreg/N15 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/pc4_to_idexreg_i [11]) );
  HS65_LH_MUX21X4 U38 ( .D0(n17672), .D1(\u_DataPath/u_ifidreg/N14 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/pc4_to_idexreg_i [10]) );
  HS65_LH_MUX21X4 U39 ( .D0(n17675), .D1(\u_DataPath/u_ifidreg/N13 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/pc4_to_idexreg_i [9]) );
  HS65_LH_MUX21X4 U40 ( .D0(n17676), .D1(\u_DataPath/u_ifidreg/N12 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/pc4_to_idexreg_i [8]) );
  HS65_LH_MUX21X4 U41 ( .D0(n17679), .D1(\u_DataPath/u_ifidreg/N11 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/pc4_to_idexreg_i [7]) );
  HS65_LH_MUX21X4 U42 ( .D0(n17681), .D1(\u_DataPath/u_ifidreg/N10 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/pc4_to_idexreg_i [6]) );
  HS65_LH_MUX21X4 U43 ( .D0(n17683), .D1(\u_DataPath/u_ifidreg/N9 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/pc4_to_idexreg_i [5]) );
  HS65_LH_MUX21X4 U44 ( .D0(n17684), .D1(\u_DataPath/u_ifidreg/N8 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/pc4_to_idexreg_i [4]) );
  HS65_LH_MUX21X4 U45 ( .D0(n17822), .D1(\u_DataPath/u_ifidreg/N7 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/pc4_to_idexreg_i [3]) );
  HS65_LH_MUX21X4 U46 ( .D0(n17686), .D1(\u_DataPath/u_ifidreg/N6 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/pc4_to_idexreg_i [2]) );
  HS65_LH_MUX21X4 U47 ( .D0(n17688), .D1(\u_DataPath/u_ifidreg/N5 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/pc4_to_idexreg_i [1]) );
  HS65_LH_MUX21X4 U48 ( .D0(n17690), .D1(\u_DataPath/u_ifidreg/N4 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/pc4_to_idexreg_i [0]) );
  HS65_LH_MUX21X4 U49 ( .D0(n38700), .D1(\u_DataPath/u_ifidreg/N51 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/immediate_ext_dec_i [15])
         );
  HS65_LH_MUX21X4 U50 ( .D0(n17731), .D1(\u_DataPath/u_ifidreg/N50 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/immediate_ext_dec_i [14])
         );
  HS65_LH_MUX21X4 U51 ( .D0(n17730), .D1(\u_DataPath/u_ifidreg/N49 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/immediate_ext_dec_i [13])
         );
  HS65_LH_MUX21X4 U52 ( .D0(n17732), .D1(\u_DataPath/u_ifidreg/N48 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/immediate_ext_dec_i [12])
         );
  HS65_LH_MUX21X4 U53 ( .D0(n17733), .D1(\u_DataPath/u_ifidreg/N47 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/immediate_ext_dec_i [11])
         );
  HS65_LH_MUX21X4 U54 ( .D0(n17734), .D1(\u_DataPath/u_ifidreg/N46 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/immediate_ext_dec_i [10])
         );
  HS65_LH_MUX21X4 U55 ( .D0(n17735), .D1(\u_DataPath/u_ifidreg/N45 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/immediate_ext_dec_i [9])
         );
  HS65_LH_MUX21X4 U56 ( .D0(n17736), .D1(\u_DataPath/u_ifidreg/N44 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/immediate_ext_dec_i [8])
         );
  HS65_LH_MUX21X4 U57 ( .D0(n17737), .D1(\u_DataPath/u_ifidreg/N43 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/immediate_ext_dec_i [7])
         );
  HS65_LH_MUX21X4 U58 ( .D0(n17738), .D1(\u_DataPath/u_ifidreg/N42 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/immediate_ext_dec_i [6])
         );
  HS65_LH_MUX21X4 U59 ( .D0(n17739), .D1(\u_DataPath/u_ifidreg/N41 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/immediate_ext_dec_i [5])
         );
  HS65_LH_MUX21X4 U60 ( .D0(n17740), .D1(\u_DataPath/u_ifidreg/N40 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/immediate_ext_dec_i [4])
         );
  HS65_LH_MUX21X4 U61 ( .D0(n38697), .D1(\u_DataPath/u_ifidreg/N39 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/immediate_ext_dec_i [3])
         );
  HS65_LH_MUX21X4 U62 ( .D0(n40161), .D1(\u_DataPath/u_ifidreg/N38 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/immediate_ext_dec_i [2])
         );
  HS65_LH_MUX21X4 U63 ( .D0(n17725), .D1(\u_DataPath/u_ifidreg/N37 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/immediate_ext_dec_i [1])
         );
  HS65_LH_MUX21X4 U64 ( .D0(n38698), .D1(\u_DataPath/u_ifidreg/N36 ), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(\u_DataPath/immediate_ext_dec_i [0])
         );
  HS65_LH_AO222X4 U72 ( .A(n17691), .B(n70), .C(n68), .D(n29703), .E(n69), .F(
        n29704), .Z(\u_DataPath/pc_4_i [0]) );
  HS65_LH_AO222X4 U73 ( .A(n70), .B(n17689), .C(n69), .D(n29770), .E(n29771), 
        .F(n68), .Z(\u_DataPath/pc_4_i [1]) );
  HS65_LH_AO222X4 U74 ( .A(n70), .B(n38493), .C(n69), .D(n38497), .E(n38563), 
        .F(n68), .Z(n17244) );
  HS65_LH_AO222X4 U75 ( .A(n70), .B(n29772), .C(n69), .D(n29773), .E(n29863), 
        .F(n68), .Z(n17243) );
  HS65_LH_AO222X4 U76 ( .A(n70), .B(n30647), .C(n69), .D(n30646), .E(n30645), 
        .F(n68), .Z(n17242) );
  HS65_LH_AO222X4 U77 ( .A(n70), .B(n30830), .C(n69), .D(n30831), .E(n30890), 
        .F(n68), .Z(n17241) );
  HS65_LH_AO222X4 U78 ( .A(n70), .B(n30738), .C(n69), .D(n30739), .E(n30829), 
        .F(n68), .Z(n17240) );
  HS65_LH_AO222X4 U79 ( .A(n70), .B(n30521), .C(n69), .D(n30522), .E(n30581), 
        .F(n68), .Z(n17239) );
  HS65_LH_AO222X4 U80 ( .A(n70), .B(n30374), .C(n69), .D(n30373), .E(n30372), 
        .F(n68), .Z(n17238) );
  HS65_LH_AO222X4 U81 ( .A(n70), .B(n30583), .C(n69), .D(n30584), .E(n30643), 
        .F(n68), .Z(n17237) );
  HS65_LH_AO222X4 U82 ( .A(n70), .B(n30240), .C(n69), .D(n30239), .E(n30238), 
        .F(n68), .Z(n17236) );
  HS65_LH_AO222X4 U83 ( .A(n70), .B(n30465), .C(n69), .D(n30466), .E(n38777), 
        .F(n68), .Z(n17235) );
  HS65_LH_AO222X4 U84 ( .A(n70), .B(n30127), .C(n69), .D(n30126), .E(n30125), 
        .F(n68), .Z(n17234) );
  HS65_LH_AO222X4 U85 ( .A(n70), .B(n30324), .C(n69), .D(n30325), .E(n38895), 
        .F(n68), .Z(n17233) );
  HS65_LH_AO222X4 U86 ( .A(n70), .B(n30029), .C(n69), .D(n30028), .E(n30027), 
        .F(n68), .Z(n17232) );
  HS65_LH_AO222X4 U87 ( .A(n70), .B(n30199), .C(n69), .D(n30200), .E(n38995), 
        .F(n68), .Z(n17231) );
  HS65_LH_AO222X4 U88 ( .A(n70), .B(n29956), .C(n69), .D(n29955), .E(n29954), 
        .F(n68), .Z(n17230) );
  HS65_LH_AO222X4 U89 ( .A(n70), .B(n30092), .C(n69), .D(n30093), .E(n39043), 
        .F(n68), .Z(n17229) );
  HS65_LH_AO222X4 U90 ( .A(n70), .B(n29906), .C(n69), .D(n29909), .E(n38967), 
        .F(n68), .Z(n17228) );
  HS65_LH_AO222X4 U91 ( .A(n70), .B(n30003), .C(n69), .D(n30005), .E(n30024), 
        .F(n68), .Z(n17227) );
  HS65_LH_AO222X4 U92 ( .A(n70), .B(n29878), .C(n69), .D(n29879), .E(n38868), 
        .F(n68), .Z(n17226) );
  HS65_LH_AO222X4 U93 ( .A(n70), .B(n29935), .C(n69), .D(n29939), .E(n38897), 
        .F(n68), .Z(n17225) );
  HS65_LH_AO222X4 U94 ( .A(n70), .B(n29865), .C(n69), .D(n29868), .E(n39116), 
        .F(n68), .Z(n17224) );
  HS65_LH_AO222X4 U95 ( .A(n70), .B(n29901), .C(n69), .D(n29902), .E(n29903), 
        .F(n68), .Z(n17223) );
  HS65_LH_AO222X4 U96 ( .A(n70), .B(n30893), .C(n69), .D(n30894), .E(n37034), 
        .F(n68), .Z(n17222) );
  HS65_LH_AO222X4 U97 ( .A(n70), .B(n39499), .C(n69), .D(n39498), .E(n39626), 
        .F(n68), .Z(n17221) );
  HS65_LH_AO222X4 U98 ( .A(n70), .B(n31115), .C(n69), .D(n31116), .E(n31178), 
        .F(n68), .Z(n17220) );
  HS65_LH_AO222X4 U99 ( .A(n70), .B(n39209), .C(n69), .D(n39207), .E(n39266), 
        .F(n68), .Z(n17219) );
  HS65_LH_AO222X4 U100 ( .A(n70), .B(n31050), .C(n69), .D(n31051), .E(n31113), 
        .F(n68), .Z(n17218) );
  HS65_LH_AO222X4 U101 ( .A(n70), .B(n39269), .C(n69), .D(n39267), .E(n39353), 
        .F(n68), .Z(n17217) );
  HS65_LH_AO222X4 U102 ( .A(n70), .B(n30986), .C(n69), .D(n30987), .E(n31049), 
        .F(n68), .Z(n17216) );
  HS65_LH_AO222X4 U103 ( .A(n70), .B(n30899), .C(n69), .D(n30898), .E(n30985), 
        .F(n68), .Z(n17215) );
  HS65_LH_AND2X4 U104 ( .A(n70), .B(iram_data[0]), .Z(
        \u_DataPath/u_ifidreg/N36 ) );
  HS65_LH_AND2X4 U105 ( .A(n70), .B(iram_data[1]), .Z(
        \u_DataPath/u_ifidreg/N37 ) );
  HS65_LH_AND2X4 U106 ( .A(n70), .B(iram_data[2]), .Z(
        \u_DataPath/u_ifidreg/N38 ) );
  HS65_LH_AND2X4 U107 ( .A(n70), .B(iram_data[3]), .Z(
        \u_DataPath/u_ifidreg/N39 ) );
  HS65_LH_AND2X4 U108 ( .A(n70), .B(iram_data[4]), .Z(
        \u_DataPath/u_ifidreg/N40 ) );
  HS65_LH_AND2X4 U109 ( .A(n70), .B(iram_data[5]), .Z(
        \u_DataPath/u_ifidreg/N41 ) );
  HS65_LH_AND2X4 U110 ( .A(n70), .B(iram_data[6]), .Z(
        \u_DataPath/u_ifidreg/N42 ) );
  HS65_LH_AND2X4 U111 ( .A(n70), .B(iram_data[7]), .Z(
        \u_DataPath/u_ifidreg/N43 ) );
  HS65_LH_AND2X4 U112 ( .A(n70), .B(iram_data[8]), .Z(
        \u_DataPath/u_ifidreg/N44 ) );
  HS65_LH_AND2X4 U113 ( .A(n70), .B(iram_data[9]), .Z(
        \u_DataPath/u_ifidreg/N45 ) );
  HS65_LH_AND2X4 U114 ( .A(n70), .B(iram_data[10]), .Z(
        \u_DataPath/u_ifidreg/N46 ) );
  HS65_LH_AND2X4 U115 ( .A(n70), .B(iram_data[11]), .Z(
        \u_DataPath/u_ifidreg/N47 ) );
  HS65_LH_AND2X4 U116 ( .A(n70), .B(iram_data[12]), .Z(
        \u_DataPath/u_ifidreg/N48 ) );
  HS65_LH_AND2X4 U117 ( .A(n70), .B(iram_data[13]), .Z(
        \u_DataPath/u_ifidreg/N49 ) );
  HS65_LH_AND2X4 U118 ( .A(n70), .B(iram_data[14]), .Z(
        \u_DataPath/u_ifidreg/N50 ) );
  HS65_LH_AND2X4 U119 ( .A(n70), .B(iram_data[15]), .Z(
        \u_DataPath/u_ifidreg/N51 ) );
  HS65_LH_AND2X4 U120 ( .A(n70), .B(iram_data[16]), .Z(
        \u_DataPath/u_ifidreg/N52 ) );
  HS65_LH_AND2X4 U121 ( .A(n70), .B(iram_data[17]), .Z(
        \u_DataPath/u_ifidreg/N53 ) );
  HS65_LH_AND2X4 U122 ( .A(n70), .B(iram_data[18]), .Z(
        \u_DataPath/u_ifidreg/N54 ) );
  HS65_LH_AND2X4 U123 ( .A(n70), .B(iram_data[19]), .Z(
        \u_DataPath/u_ifidreg/N55 ) );
  HS65_LH_AND2X4 U124 ( .A(n70), .B(iram_data[20]), .Z(
        \u_DataPath/u_ifidreg/N56 ) );
  HS65_LH_AND2X4 U125 ( .A(n70), .B(iram_data[21]), .Z(
        \u_DataPath/u_ifidreg/N57 ) );
  HS65_LH_AND2X4 U126 ( .A(n70), .B(iram_data[22]), .Z(
        \u_DataPath/u_ifidreg/N58 ) );
  HS65_LH_AND2X4 U127 ( .A(n70), .B(iram_data[23]), .Z(
        \u_DataPath/u_ifidreg/N59 ) );
  HS65_LH_AND2X4 U128 ( .A(n70), .B(iram_data[24]), .Z(
        \u_DataPath/u_ifidreg/N60 ) );
  HS65_LH_AND2X4 U129 ( .A(n70), .B(iram_data[25]), .Z(
        \u_DataPath/u_ifidreg/N61 ) );
  HS65_LH_NAND2AX4 U130 ( .A(iram_data[26]), .B(n70), .Z(
        \u_DataPath/u_ifidreg/N62 ) );
  HS65_LH_AND2X4 U131 ( .A(n70), .B(iram_data[27]), .Z(
        \u_DataPath/u_ifidreg/N63 ) );
  HS65_LH_NAND2AX4 U132 ( .A(iram_data[28]), .B(n70), .Z(
        \u_DataPath/u_ifidreg/N64 ) );
  HS65_LH_AND2X4 U133 ( .A(n70), .B(iram_data[29]), .Z(
        \u_DataPath/u_ifidreg/N65 ) );
  HS65_LH_NAND2AX4 U134 ( .A(iram_data[30]), .B(n70), .Z(
        \u_DataPath/u_ifidreg/N66 ) );
  HS65_LH_AND2X4 U135 ( .A(n70), .B(iram_data[31]), .Z(
        \u_DataPath/u_ifidreg/N67 ) );
  HS65_LH_CNIVX3 U151 ( .A(rst), .Z(n2733) );
  HS65_LH_AO22X4 U153 ( .A(n17841), .B(n74), .C(n73), .D(n17840), .Z(
        \u_DataPath/RFaddr_out_memwb_i [0]) );
  HS65_LH_AO22X4 U154 ( .A(n17838), .B(n74), .C(n73), .D(n17837), .Z(
        \u_DataPath/RFaddr_out_memwb_i [1]) );
  HS65_LH_AO22X4 U155 ( .A(n17835), .B(n74), .C(n73), .D(n17834), .Z(
        \u_DataPath/RFaddr_out_memwb_i [2]) );
  HS65_LH_AO22X4 U156 ( .A(n17831), .B(n74), .C(n73), .D(n17832), .Z(
        \u_DataPath/RFaddr_out_memwb_i [3]) );
  HS65_LH_AO22X4 U157 ( .A(n17829), .B(n74), .C(n73), .D(n17828), .Z(
        \u_DataPath/RFaddr_out_memwb_i [4]) );
  HS65_LH_AND2X4 U508 ( .A(\u_DataPath/u_execute/ovf_i ), .B(n2733), .Z(
        \u_DataPath/u_execute/psw_status_i [1]) );
  HS65_LH_OR3X4 U550 ( .A(\u_DataPath/u_idexreg/N13 ), .B(n180), .C(
        \u_DataPath/u_idexreg/N11 ), .Z(\u_DataPath/u_idexreg/N10 ) );
  HS65_LH_MX41X4 U604 ( .D0(n35219), .S0(\u_DataPath/u_idexreg/N19 ), .D1(
        n35267), .S1(n214), .D2(n35231), .S2(n227), .D3(n244), .S3(n35218), 
        .Z(\u_DataPath/cw_to_ex_i [0]) );
  HS65_LH_OAI21X2 U628 ( .A(\u_DataPath/u_idexreg/N8 ), .B(n227), .C(n35419), 
        .Z(n228) );
  HS65_LH_OAI222X2 U643 ( .A(n254), .B(n40524), .C(n253), .D(n34580), .E(n284), 
        .F(n34670), .Z(\u_DataPath/cw_to_ex_i [4]) );
  HS65_LH_NAND3AX3 U645 ( .A(n34002), .B(n33995), .C(n255), .Z(n283) );
  HS65_LH_NOR4ABX2 U659 ( .A(\u_DataPath/u_idexreg/N19 ), .B(n33918), .C(
        n33916), .D(n33929), .Z(\u_DataPath/cw_to_ex_i [15]) );
  HS65_LH_NOR3AX2 U660 ( .A(n34016), .B(n279), .C(n34017), .Z(
        \u_DataPath/u_idexreg/N20 ) );
  HS65_LH_AND2X4 U662 ( .A(\u_DataPath/u_idexreg/N8 ), .B(n17774), .Z(
        \u_DataPath/cw_to_ex_i [19]) );
  HS65_LH_NAND4ABX3 U664 ( .A(\u_DataPath/u_idexreg/N21 ), .B(
        \u_DataPath/u_idexreg/N20 ), .C(n285), .D(n284), .Z(
        \u_DataPath/cw_exmem_i [10]) );
  HS65_LH_AND2X4 U699 ( .A(n40481), .B(n2733), .Z(\u_DataPath/reg_write_i ) );
  HS65_LH_AND2X4 U700 ( .A(n40474), .B(n2733), .Z(\u_DataPath/cw_towb_i [1])
         );
  HS65_LH_AND2X4 U701 ( .A(n34053), .B(n2733), .Z(\u_DataPath/cw_towb_i [0])
         );
  HS65_LH_OAI21X2 U713 ( .A(n292), .B(n307), .C(n320), .Z(
        \u_DataPath/from_mem_data_out_i [31]) );
  HS65_LH_OAI21X2 U715 ( .A(n293), .B(n307), .C(n320), .Z(
        \u_DataPath/from_mem_data_out_i [30]) );
  HS65_LH_OAI21X2 U717 ( .A(n294), .B(n307), .C(n320), .Z(
        \u_DataPath/from_mem_data_out_i [29]) );
  HS65_LH_OAI21X2 U719 ( .A(n295), .B(n307), .C(n320), .Z(
        \u_DataPath/from_mem_data_out_i [28]) );
  HS65_LH_OAI21X2 U721 ( .A(n296), .B(n307), .C(n320), .Z(
        \u_DataPath/from_mem_data_out_i [27]) );
  HS65_LH_OAI21X2 U723 ( .A(n297), .B(n307), .C(n320), .Z(
        \u_DataPath/from_mem_data_out_i [26]) );
  HS65_LH_OAI21X2 U725 ( .A(n298), .B(n307), .C(n320), .Z(
        \u_DataPath/from_mem_data_out_i [25]) );
  HS65_LH_OAI21X2 U727 ( .A(n299), .B(n307), .C(n320), .Z(
        \u_DataPath/from_mem_data_out_i [24]) );
  HS65_LH_OAI21X2 U729 ( .A(n300), .B(n307), .C(n320), .Z(
        \u_DataPath/from_mem_data_out_i [23]) );
  HS65_LH_OAI21X2 U731 ( .A(n301), .B(n307), .C(n320), .Z(
        \u_DataPath/from_mem_data_out_i [22]) );
  HS65_LH_OAI21X2 U733 ( .A(n302), .B(n307), .C(n320), .Z(
        \u_DataPath/from_mem_data_out_i [21]) );
  HS65_LH_OAI21X2 U735 ( .A(n303), .B(n307), .C(n320), .Z(
        \u_DataPath/from_mem_data_out_i [20]) );
  HS65_LH_OAI21X2 U737 ( .A(n304), .B(n307), .C(n320), .Z(
        \u_DataPath/from_mem_data_out_i [19]) );
  HS65_LH_OAI21X2 U739 ( .A(n305), .B(n307), .C(n320), .Z(
        \u_DataPath/from_mem_data_out_i [18]) );
  HS65_LH_OAI21X2 U741 ( .A(n306), .B(n307), .C(n320), .Z(
        \u_DataPath/from_mem_data_out_i [17]) );
  HS65_LH_OAI21X2 U743 ( .A(n308), .B(n307), .C(n320), .Z(
        \u_DataPath/from_mem_data_out_i [16]) );
  HS65_LH_CB4I1X4 U745 ( .A(n33944), .B(n33955), .C(n33951), .D(n309), .Z(n335) );
  HS65_LH_AO222X4 U765 ( .A(n34227), .B(n337), .C(Data_out_fromRAM[23]), .D(
        n336), .E(Data_out_fromRAM[7]), .F(n335), .Z(
        \u_DataPath/from_mem_data_out_i [7]) );
  HS65_LH_AO222X4 U767 ( .A(n325), .B(n337), .C(n336), .D(Data_out_fromRAM[22]), .E(n335), .F(Data_out_fromRAM[6]), .Z(\u_DataPath/from_mem_data_out_i [6])
         );
  HS65_LH_AO222X4 U769 ( .A(n33893), .B(n337), .C(n336), .D(
        Data_out_fromRAM[21]), .E(n335), .F(Data_out_fromRAM[5]), .Z(
        \u_DataPath/from_mem_data_out_i [5]) );
  HS65_LH_AO222X4 U771 ( .A(n33901), .B(n337), .C(n336), .D(
        Data_out_fromRAM[20]), .E(n335), .F(Data_out_fromRAM[4]), .Z(
        \u_DataPath/from_mem_data_out_i [4]) );
  HS65_LH_AO222X4 U773 ( .A(n33934), .B(n337), .C(n336), .D(
        Data_out_fromRAM[19]), .E(n335), .F(Data_out_fromRAM[3]), .Z(
        \u_DataPath/from_mem_data_out_i [3]) );
  HS65_LH_AO222X4 U775 ( .A(n33952), .B(n337), .C(n336), .D(
        Data_out_fromRAM[18]), .E(n335), .F(Data_out_fromRAM[2]), .Z(
        \u_DataPath/from_mem_data_out_i [2]) );
  HS65_LH_AO222X4 U777 ( .A(n33909), .B(n337), .C(n336), .D(
        Data_out_fromRAM[17]), .E(n335), .F(Data_out_fromRAM[1]), .Z(
        \u_DataPath/from_mem_data_out_i [1]) );
  HS65_LH_AO222X4 U779 ( .A(n33888), .B(n337), .C(n336), .D(
        Data_out_fromRAM[16]), .E(n335), .F(Data_out_fromRAM[0]), .Z(
        \u_DataPath/from_mem_data_out_i [0]) );
  HS65_LH_AND2X4 U847 ( .A(n33829), .B(n2733), .Z(\u_DataPath/cw_memwb_i [2])
         );
  HS65_LH_AND2X4 U849 ( .A(n33969), .B(n2733), .Z(\u_DataPath/cw_tomem_i [8])
         );
  HS65_LH_AND2X4 U850 ( .A(n34262), .B(n2733), .Z(\u_DataPath/cw_tomem_i [7])
         );
  HS65_LH_AND2X4 U851 ( .A(n31929), .B(n2733), .Z(\u_DataPath/cw_tomem_i [6])
         );
  HS65_LH_AND2X4 U852 ( .A(n33961), .B(n2733), .Z(\u_DataPath/cw_tomem_i [5])
         );
  HS65_LH_AND2X4 U853 ( .A(n31928), .B(n2733), .Z(\u_DataPath/cw_tomem_i [4])
         );
  HS65_LH_AND2X4 U855 ( .A(n17790), .B(n2733), .Z(\u_DataPath/cw_memwb_i [0])
         );
  HS65_LH_AND2X4 U856 ( .A(n34372), .B(n2733), .Z(\u_DataPath/jump_i ) );
  HS65_LH_AND2X4 U857 ( .A(n39422), .B(n2733), .Z(\u_DataPath/cw_tomem_i [0])
         );
  HS65_LH_AO22X4 U860 ( .A(n15473), .B(n348), .C(n347), .D(n29559), .Z(
        \u_DataPath/jump_address_i [31]) );
  HS65_LH_AO22X4 U861 ( .A(n14192), .B(n348), .C(n347), .D(n15396), .Z(
        \u_DataPath/jump_address_i [30]) );
  HS65_LH_AO22X4 U862 ( .A(n14180), .B(n348), .C(n347), .D(n14031), .Z(
        \u_DataPath/jump_address_i [29]) );
  HS65_LH_AO22X4 U863 ( .A(n14162), .B(n348), .C(n347), .D(n14850), .Z(
        \u_DataPath/jump_address_i [28]) );
  HS65_LH_AO22X4 U864 ( .A(n14212), .B(n348), .C(n347), .D(n14627), .Z(
        \u_DataPath/jump_address_i [27]) );
  HS65_LH_AO22X4 U865 ( .A(n14198), .B(n348), .C(n347), .D(n14553), .Z(
        \u_DataPath/jump_address_i [26]) );
  HS65_LH_AO22X4 U866 ( .A(n14171), .B(n348), .C(n347), .D(n14752), .Z(
        \u_DataPath/jump_address_i [25]) );
  HS65_LH_AO22X4 U867 ( .A(n14165), .B(n348), .C(n347), .D(n14822), .Z(
        \u_DataPath/jump_address_i [24]) );
  HS65_LH_AO22X4 U868 ( .A(n14195), .B(n348), .C(n347), .D(n14642), .Z(
        \u_DataPath/jump_address_i [23]) );
  HS65_LH_AO22X4 U869 ( .A(n14159), .B(n348), .C(n347), .D(n14559), .Z(
        \u_DataPath/jump_address_i [22]) );
  HS65_LH_AO22X4 U870 ( .A(n14177), .B(n348), .C(n347), .D(n15268), .Z(
        \u_DataPath/jump_address_i [21]) );
  HS65_LH_AO22X4 U871 ( .A(n14153), .B(n348), .C(n347), .D(
        \u_DataPath/u_execute/A_inALU_i [20]), .Z(
        \u_DataPath/jump_address_i [20]) );
  HS65_LH_AO22X4 U872 ( .A(n14204), .B(n348), .C(n347), .D(n14388), .Z(
        \u_DataPath/jump_address_i [19]) );
  HS65_LH_AO22X4 U873 ( .A(n14144), .B(n348), .C(n347), .D(n15096), .Z(
        \u_DataPath/jump_address_i [18]) );
  HS65_LH_AO22X4 U874 ( .A(n14147), .B(n348), .C(n347), .D(n15018), .Z(
        \u_DataPath/jump_address_i [17]) );
  HS65_LH_AO22X4 U875 ( .A(n14150), .B(n348), .C(n347), .D(n14997), .Z(
        \u_DataPath/jump_address_i [16]) );
  HS65_LH_AO22X4 U876 ( .A(n14303), .B(n348), .C(n347), .D(n14035), .Z(
        \u_DataPath/jump_address_i [15]) );
  HS65_LH_AO22X4 U877 ( .A(n14306), .B(n348), .C(n347), .D(n14036), .Z(
        \u_DataPath/jump_address_i [14]) );
  HS65_LH_AO22X4 U878 ( .A(n14183), .B(n348), .C(n347), .D(n14032), .Z(
        \u_DataPath/jump_address_i [13]) );
  HS65_LH_AO22X4 U879 ( .A(n14189), .B(n348), .C(n347), .D(
        \u_DataPath/u_execute/A_inALU_i [12]), .Z(
        \u_DataPath/jump_address_i [12]) );
  HS65_LH_AO22X4 U880 ( .A(n14208), .B(n348), .C(n347), .D(n14358), .Z(
        \u_DataPath/jump_address_i [11]) );
  HS65_LH_AO22X4 U881 ( .A(n14201), .B(n348), .C(n347), .D(n14033), .Z(
        \u_DataPath/jump_address_i [10]) );
  HS65_LH_AO22X4 U882 ( .A(n18007), .B(n348), .C(n347), .D(n14545), .Z(
        \u_DataPath/jump_address_i [9]) );
  HS65_LH_AO22X4 U883 ( .A(n18011), .B(n348), .C(n347), .D(n14030), .Z(
        \u_DataPath/jump_address_i [8]) );
  HS65_LH_AO22X4 U884 ( .A(n18001), .B(n348), .C(n347), .D(n14583), .Z(
        \u_DataPath/jump_address_i [7]) );
  HS65_LH_AO22X4 U885 ( .A(n18015), .B(n348), .C(n347), .D(n14029), .Z(
        \u_DataPath/jump_address_i [6]) );
  HS65_LH_AO22X4 U886 ( .A(n18005), .B(n348), .C(n347), .D(n14734), .Z(
        \u_DataPath/jump_address_i [5]) );
  HS65_LH_AO22X4 U887 ( .A(n17904), .B(n348), .C(n347), .D(n14918), .Z(
        \u_DataPath/jump_address_i [4]) );
  HS65_LH_AO22X4 U888 ( .A(n17974), .B(n348), .C(n347), .D(n15246), .Z(
        \u_DataPath/jump_address_i [3]) );
  HS65_LH_AO22X4 U889 ( .A(n17881), .B(n348), .C(n347), .D(n15324), .Z(
        \u_DataPath/jump_address_i [2]) );
  HS65_LH_AO22X4 U890 ( .A(n17866), .B(n348), .C(n347), .D(n15502), .Z(
        \u_DataPath/jump_address_i [1]) );
  HS65_LH_AO22X4 U891 ( .A(n17863), .B(n348), .C(n347), .D(n15163), .Z(
        \u_DataPath/jump_address_i [0]) );
  HS65_LH_AND2X4 U892 ( .A(n15580), .B(n2733), .Z(
        \u_DataPath/branch_target_i [31]) );
  HS65_LH_AND2X4 U923 ( .A(n34014), .B(n2733), .Z(
        \u_DataPath/branch_target_i [0]) );
  HS65_LH_OAI21X2 U1593 ( .A(n15572), .B(n18157), .C(n17286), .Z(
        \u_DataPath/dataOut_exe_i [31]) );
  HS65_LH_AO222X4 U1594 ( .A(n15577), .B(n17327), .C(n17326), .D(n17953), .E(
        n17951), .F(n17525), .Z(\u_DataPath/dataOut_exe_i [30]) );
  HS65_LH_AO222X4 U1595 ( .A(n17936), .B(n17327), .C(n17326), .D(n17937), .E(
        n17938), .F(n17525), .Z(\u_DataPath/dataOut_exe_i [29]) );
  HS65_LH_AO222X4 U1596 ( .A(n17910), .B(n17327), .C(n17326), .D(n17911), .E(
        n17912), .F(n17525), .Z(\u_DataPath/dataOut_exe_i [28]) );
  HS65_LH_AO222X4 U1597 ( .A(n17990), .B(n17327), .C(n17326), .D(n17992), .E(
        n17993), .F(n17525), .Z(\u_DataPath/dataOut_exe_i [27]) );
  HS65_LH_AO222X4 U1598 ( .A(n17959), .B(n17327), .C(n17326), .D(n17960), .E(
        n17961), .F(n17525), .Z(\u_DataPath/dataOut_exe_i [26]) );
  HS65_LH_OAI21X2 U1600 ( .A(n17924), .B(n18157), .C(n17285), .Z(
        \u_DataPath/dataOut_exe_i [25]) );
  HS65_LH_OAI21X2 U1602 ( .A(n17918), .B(n18157), .C(n17284), .Z(
        \u_DataPath/dataOut_exe_i [24]) );
  HS65_LH_AO222X4 U1603 ( .A(n32609), .B(n1067), .C(n1065), .D(n31219), .E(
        n31216), .F(n1040), .Z(\u_DataPath/dataOut_exe_i [23]) );
  HS65_LH_AO222X4 U1604 ( .A(n31294), .B(n1067), .C(n1065), .D(n31295), .E(
        n31296), .F(n1040), .Z(\u_DataPath/dataOut_exe_i [22]) );
  HS65_LH_OAI21X2 U1606 ( .A(n31869), .B(n1059), .C(n1033), .Z(
        \u_DataPath/dataOut_exe_i [21]) );
  HS65_LH_AO222X4 U1607 ( .A(n31811), .B(n1067), .C(n1065), .D(n31810), .E(
        n31816), .F(n1040), .Z(\u_DataPath/dataOut_exe_i [20]) );
  HS65_LH_OAI21X2 U1609 ( .A(n32158), .B(n1059), .C(n1036), .Z(
        \u_DataPath/dataOut_exe_i [19]) );
  HS65_LH_AO222X4 U1610 ( .A(n32517), .B(n1067), .C(n1065), .D(n32515), .E(
        n32566), .F(n1040), .Z(\u_DataPath/dataOut_exe_i [18]) );
  HS65_LH_AO222X4 U1611 ( .A(n32710), .B(n1067), .C(n1065), .D(n32711), .E(
        n32771), .F(n1040), .Z(\u_DataPath/dataOut_exe_i [17]) );
  HS65_LH_OAI21X2 U1613 ( .A(n32627), .B(n1059), .C(n1041), .Z(
        \u_DataPath/dataOut_exe_i [16]) );
  HS65_LH_OAI21X2 U1615 ( .A(n32772), .B(n1059), .C(n1043), .Z(
        \u_DataPath/dataOut_exe_i [15]) );
  HS65_LH_AO22X4 U1616 ( .A(n31765), .B(n1065), .C(n1067), .D(n15556), .Z(
        \u_DataPath/dataOut_exe_i [14]) );
  HS65_LH_OAI21X2 U1618 ( .A(n32849), .B(n1059), .C(n1046), .Z(
        \u_DataPath/dataOut_exe_i [13]) );
  HS65_LH_OAI21X2 U1620 ( .A(n32930), .B(n1059), .C(n1048), .Z(
        \u_DataPath/dataOut_exe_i [12]) );
  HS65_LH_AO22X4 U1621 ( .A(n33013), .B(n1065), .C(n1067), .D(n33020), .Z(
        \u_DataPath/dataOut_exe_i [11]) );
  HS65_LH_AO22X4 U1622 ( .A(n33228), .B(n1065), .C(n1067), .D(n29700), .Z(
        \u_DataPath/dataOut_exe_i [10]) );
  HS65_LH_AO22X4 U1623 ( .A(n33472), .B(n1065), .C(n1067), .D(n33471), .Z(
        \u_DataPath/dataOut_exe_i [9]) );
  HS65_LH_AO22X4 U1624 ( .A(n33656), .B(n1065), .C(n1067), .D(n33655), .Z(
        \u_DataPath/dataOut_exe_i [8]) );
  HS65_LH_OAI21X2 U1626 ( .A(n33609), .B(n1059), .C(n1054), .Z(
        \u_DataPath/dataOut_exe_i [7]) );
  HS65_LH_OAI21X2 U1628 ( .A(n33517), .B(n1059), .C(n1056), .Z(
        \u_DataPath/dataOut_exe_i [6]) );
  HS65_LH_OAI21X2 U1630 ( .A(n33553), .B(n1059), .C(n1058), .Z(
        \u_DataPath/dataOut_exe_i [5]) );
  HS65_LH_AO22X4 U1631 ( .A(n33699), .B(n1065), .C(n1067), .D(n33732), .Z(
        \u_DataPath/dataOut_exe_i [4]) );
  HS65_LH_AO22X4 U1632 ( .A(n33787), .B(n1065), .C(n1067), .D(n33796), .Z(
        \u_DataPath/dataOut_exe_i [3]) );
  HS65_LH_AO22X4 U1633 ( .A(n33850), .B(n1065), .C(n1067), .D(n33849), .Z(
        \u_DataPath/dataOut_exe_i [2]) );
  HS65_LH_AND2X4 U1634 ( .A(n32348), .B(n2733), .Z(n1066) );
  HS65_LH_AO222X4 U1635 ( .A(n32349), .B(n1067), .C(n1065), .D(n32343), .E(
        n32341), .F(n1066), .Z(\u_DataPath/dataOut_exe_i [1]) );
  HS65_LH_AO222X4 U1636 ( .A(n32506), .B(n1067), .C(n1066), .D(n32505), .E(
        n1065), .F(n32512), .Z(\u_DataPath/dataOut_exe_i [0]) );
  HS65_LH_AND2X4 U1683 ( .A(n39761), .B(n2733), .Z(\u_DataPath/u_idexreg/N39 )
         );
  HS65_LH_AND2X4 U1684 ( .A(n39739), .B(n2733), .Z(\u_DataPath/u_idexreg/N38 )
         );
  HS65_LH_AND2X4 U1685 ( .A(n38648), .B(n2733), .Z(\u_DataPath/u_idexreg/N37 )
         );
  HS65_LH_AND2X4 U1686 ( .A(n29722), .B(n2733), .Z(\u_DataPath/u_idexreg/N36 )
         );
  HS65_LH_AND2X4 U1687 ( .A(n39828), .B(n2733), .Z(\u_DataPath/u_idexreg/N35 )
         );
  HS65_LH_AND2X4 U1688 ( .A(n39695), .B(n2733), .Z(\u_DataPath/u_idexreg/N34 )
         );
  HS65_LH_AND2X4 U1689 ( .A(n39630), .B(n2733), .Z(\u_DataPath/u_idexreg/N33 )
         );
  HS65_LH_AND2X4 U1690 ( .A(n39651), .B(n2733), .Z(\u_DataPath/u_idexreg/N32 )
         );
  HS65_LH_AND2X4 U1691 ( .A(n39270), .B(n2733), .Z(\u_DataPath/u_idexreg/N31 )
         );
  HS65_LH_NOR2AX3 U1693 ( .A(n40205), .B(rst), .Z(\u_DataPath/u_idexreg/N29 )
         );
  HS65_LH_AND2X4 U1698 ( .A(n39378), .B(n2733), .Z(
        \u_DataPath/pc_4_to_ex_i [31]) );
  HS65_LH_AND2X4 U1699 ( .A(n39356), .B(n2733), .Z(
        \u_DataPath/pc_4_to_ex_i [30]) );
  HS65_LH_AND2X4 U1700 ( .A(n39850), .B(n2733), .Z(
        \u_DataPath/pc_4_to_ex_i [29]) );
  HS65_LH_AND2X4 U1701 ( .A(n39872), .B(n2733), .Z(
        \u_DataPath/pc_4_to_ex_i [28]) );
  HS65_LH_AND2X4 U1702 ( .A(n39894), .B(n2733), .Z(
        \u_DataPath/pc_4_to_ex_i [27]) );
  HS65_LH_AND2X4 U1703 ( .A(n39916), .B(n2733), .Z(
        \u_DataPath/pc_4_to_ex_i [26]) );
  HS65_LH_AND2X4 U1704 ( .A(n39938), .B(n2733), .Z(
        \u_DataPath/pc_4_to_ex_i [25]) );
  HS65_LH_AND2X4 U1705 ( .A(n39400), .B(n2733), .Z(
        \u_DataPath/pc_4_to_ex_i [24]) );
  HS65_LH_AND2X4 U1706 ( .A(n39960), .B(n2733), .Z(
        \u_DataPath/pc_4_to_ex_i [23]) );
  HS65_LH_AND2X4 U1707 ( .A(n39982), .B(n2733), .Z(
        \u_DataPath/pc_4_to_ex_i [22]) );
  HS65_LH_AND2X4 U1708 ( .A(n40004), .B(n2733), .Z(
        \u_DataPath/pc_4_to_ex_i [21]) );
  HS65_LH_AND2X4 U1709 ( .A(n40026), .B(n2733), .Z(
        \u_DataPath/pc_4_to_ex_i [20]) );
  HS65_LH_AND2X4 U1710 ( .A(n40048), .B(n2733), .Z(
        \u_DataPath/pc_4_to_ex_i [19]) );
  HS65_LH_AND2X4 U1711 ( .A(n40070), .B(n2733), .Z(
        \u_DataPath/pc_4_to_ex_i [18]) );
  HS65_LH_AND2X4 U1712 ( .A(n40092), .B(n2733), .Z(
        \u_DataPath/pc_4_to_ex_i [17]) );
  HS65_LH_AND2X4 U1713 ( .A(n39783), .B(n2733), .Z(
        \u_DataPath/pc_4_to_ex_i [16]) );
  HS65_LH_AND2X4 U1714 ( .A(n40114), .B(n2733), .Z(
        \u_DataPath/pc_4_to_ex_i [15]) );
  HS65_LH_AND2X4 U1715 ( .A(n39827), .B(n2733), .Z(
        \u_DataPath/pc_4_to_ex_i [14]) );
  HS65_LH_AND2X4 U1716 ( .A(n40136), .B(n2733), .Z(
        \u_DataPath/pc_4_to_ex_i [13]) );
  HS65_LH_AND2X4 U1717 ( .A(n39805), .B(n2733), .Z(
        \u_DataPath/pc_4_to_ex_i [12]) );
  HS65_LH_AND2X4 U1718 ( .A(n39717), .B(n2733), .Z(
        \u_DataPath/pc_4_to_ex_i [11]) );
  HS65_LH_AND2X4 U1719 ( .A(n39355), .B(n2733), .Z(
        \u_DataPath/pc_4_to_ex_i [10]) );
  HS65_LH_AND2X4 U1720 ( .A(n33090), .B(n2733), .Z(
        \u_DataPath/pc_4_to_ex_i [9]) );
  HS65_LH_AND2X4 U1721 ( .A(n33082), .B(n2733), .Z(
        \u_DataPath/pc_4_to_ex_i [8]) );
  HS65_LH_AND2X4 U1722 ( .A(n33074), .B(n2733), .Z(
        \u_DataPath/pc_4_to_ex_i [7]) );
  HS65_LH_AND2X4 U1723 ( .A(n33080), .B(n2733), .Z(
        \u_DataPath/pc_4_to_ex_i [6]) );
  HS65_LH_AND2X4 U1724 ( .A(n33071), .B(n2733), .Z(
        \u_DataPath/pc_4_to_ex_i [5]) );
  HS65_LH_AND2X4 U1725 ( .A(n33073), .B(n2733), .Z(
        \u_DataPath/pc_4_to_ex_i [4]) );
  HS65_LH_AND2X4 U1726 ( .A(n33079), .B(n2733), .Z(
        \u_DataPath/pc_4_to_ex_i [3]) );
  HS65_LH_AND2X4 U1727 ( .A(n33087), .B(n2733), .Z(
        \u_DataPath/pc_4_to_ex_i [2]) );
  HS65_LH_AND2X4 U1728 ( .A(n33081), .B(n2733), .Z(
        \u_DataPath/u_execute/link_value_i [1]) );
  HS65_LH_AND2X4 U1729 ( .A(n34012), .B(n2733), .Z(
        \u_DataPath/u_execute/link_value_i [0]) );
  HS65_LH_OAI21X2 U1804 ( .A(n40883), .B(n40895), .C(n1895), .Z(n1152) );
  HS65_LH_OAI21X2 U1805 ( .A(n17214), .B(n1952), .C(n1152), .Z(
        \u_DataPath/data_read_ex_1_i [31]) );
  HS65_LH_OAI21X2 U1828 ( .A(n38242), .B(n38239), .C(n1895), .Z(n1175) );
  HS65_LH_OAI21X2 U1829 ( .A(n17214), .B(n1976), .C(n1175), .Z(
        \u_DataPath/data_read_ex_1_i [30]) );
  HS65_LH_OAI21X2 U1852 ( .A(n38327), .B(n38376), .C(n1895), .Z(n1198) );
  HS65_LH_OAI21X2 U1853 ( .A(n17214), .B(n2000), .C(n1198), .Z(
        \u_DataPath/data_read_ex_1_i [29]) );
  HS65_LH_OAI21X2 U1876 ( .A(n37501), .B(n37500), .C(n1895), .Z(n1221) );
  HS65_LH_OAI21X2 U1877 ( .A(n17214), .B(n2024), .C(n1221), .Z(
        \u_DataPath/data_read_ex_1_i [28]) );
  HS65_LH_OAI21X2 U1900 ( .A(n37855), .B(n37853), .C(n1895), .Z(n1244) );
  HS65_LH_OAI21X2 U1901 ( .A(n17214), .B(n2048), .C(n1244), .Z(
        \u_DataPath/data_read_ex_1_i [27]) );
  HS65_LH_OAI21X2 U1924 ( .A(n38181), .B(n38233), .C(n1895), .Z(n1267) );
  HS65_LH_OAI21X2 U1925 ( .A(n17214), .B(n2072), .C(n1267), .Z(
        \u_DataPath/data_read_ex_1_i [26]) );
  HS65_LH_OAI21X2 U1948 ( .A(n37341), .B(n37338), .C(n1895), .Z(n1290) );
  HS65_LH_OAI21X2 U1949 ( .A(n17214), .B(n2096), .C(n1290), .Z(
        \u_DataPath/data_read_ex_1_i [25]) );
  HS65_LH_OAI21X2 U1972 ( .A(n37718), .B(n37715), .C(n1895), .Z(n1313) );
  HS65_LH_OAI21X2 U1973 ( .A(n17214), .B(n2120), .C(n1313), .Z(
        \u_DataPath/data_read_ex_1_i [24]) );
  HS65_LH_OAI21X2 U1996 ( .A(n37422), .B(n37421), .C(n1895), .Z(n1336) );
  HS65_LH_OAI21X2 U1997 ( .A(n17214), .B(n2144), .C(n1336), .Z(
        \u_DataPath/data_read_ex_1_i [23]) );
  HS65_LH_OAI21X2 U2020 ( .A(n37586), .B(n37588), .C(n1895), .Z(n1359) );
  HS65_LH_OAI21X2 U2021 ( .A(n17214), .B(n2168), .C(n1359), .Z(
        \u_DataPath/data_read_ex_1_i [22]) );
  HS65_LH_OAI21X2 U2044 ( .A(n37665), .B(n37664), .C(n1895), .Z(n1382) );
  HS65_LH_OAI21X2 U2045 ( .A(n17214), .B(n2192), .C(n1382), .Z(
        \u_DataPath/data_read_ex_1_i [21]) );
  HS65_LH_OAI21X2 U2068 ( .A(n38099), .B(n38098), .C(n1895), .Z(n1405) );
  HS65_LH_OAI21X2 U2069 ( .A(n17214), .B(n2216), .C(n1405), .Z(
        \u_DataPath/data_read_ex_1_i [20]) );
  HS65_LH_OAI21X2 U2092 ( .A(n37803), .B(n37802), .C(n1895), .Z(n1428) );
  HS65_LH_OAI21X2 U2093 ( .A(n17214), .B(n2240), .C(n1428), .Z(
        \u_DataPath/data_read_ex_1_i [19]) );
  HS65_LH_OAI21X2 U2116 ( .A(n37124), .B(n37126), .C(n1895), .Z(n1451) );
  HS65_LH_OAI21X2 U2117 ( .A(n17213), .B(n2264), .C(n1451), .Z(
        \u_DataPath/data_read_ex_1_i [18]) );
  HS65_LH_OAI21X2 U2140 ( .A(n37071), .B(n37074), .C(n1895), .Z(n1474) );
  HS65_LH_OAI21X2 U2141 ( .A(n17213), .B(n2288), .C(n1474), .Z(
        \u_DataPath/data_read_ex_1_i [17]) );
  HS65_LH_OAI21X2 U2164 ( .A(n37259), .B(n37258), .C(n1895), .Z(n1497) );
  HS65_LH_OAI21X2 U2165 ( .A(n17213), .B(n2312), .C(n1497), .Z(
        \u_DataPath/data_read_ex_1_i [16]) );
  HS65_LH_OAI21X2 U2188 ( .A(n32574), .B(n32577), .C(n1895), .Z(n1520) );
  HS65_LH_OAI21X2 U2189 ( .A(n17213), .B(n2336), .C(n1520), .Z(
        \u_DataPath/data_read_ex_1_i [15]) );
  HS65_LH_OAI21X2 U2212 ( .A(n31770), .B(n31764), .C(n1895), .Z(n1543) );
  HS65_LH_OAI21X2 U2213 ( .A(n17213), .B(n2360), .C(n1543), .Z(
        \u_DataPath/data_read_ex_1_i [14]) );
  HS65_LH_OAI21X2 U2236 ( .A(n32814), .B(n32847), .C(n1895), .Z(n1566) );
  HS65_LH_OAI21X2 U2237 ( .A(n17213), .B(n2384), .C(n1566), .Z(
        \u_DataPath/data_read_ex_1_i [13]) );
  HS65_LH_OAI21X2 U2260 ( .A(n32888), .B(n32887), .C(n1895), .Z(n1589) );
  HS65_LH_OAI21X2 U2261 ( .A(n17213), .B(n2408), .C(n1589), .Z(
        \u_DataPath/data_read_ex_1_i [12]) );
  HS65_LH_OAI21X2 U2284 ( .A(n32962), .B(n32963), .C(n1895), .Z(n1612) );
  HS65_LH_OAI21X2 U2285 ( .A(n17213), .B(n2432), .C(n1612), .Z(
        \u_DataPath/data_read_ex_1_i [11]) );
  HS65_LH_OAI21X2 U2308 ( .A(n33177), .B(n33206), .C(n1895), .Z(n1635) );
  HS65_LH_OAI21X2 U2309 ( .A(n17213), .B(n2456), .C(n1635), .Z(
        \u_DataPath/data_read_ex_1_i [10]) );
  HS65_LH_OAI21X2 U2332 ( .A(n33367), .B(n33395), .C(n1895), .Z(n1658) );
  HS65_LH_OAI21X2 U2333 ( .A(n17213), .B(n2480), .C(n1658), .Z(
        \u_DataPath/data_read_ex_1_i [9]) );
  HS65_LH_OAI21X2 U2356 ( .A(n33400), .B(n33410), .C(n1895), .Z(n1681) );
  HS65_LH_OAI21X2 U2357 ( .A(n17213), .B(n2504), .C(n1681), .Z(
        \u_DataPath/data_read_ex_1_i [8]) );
  HS65_LH_OAI21X2 U2380 ( .A(n33436), .B(n33467), .C(n1895), .Z(n1704) );
  HS65_LH_OAI21X2 U2381 ( .A(n17213), .B(n2528), .C(n1704), .Z(
        \u_DataPath/data_read_ex_1_i [7]) );
  HS65_LH_OAI21X2 U2404 ( .A(n33271), .B(n33272), .C(n1895), .Z(n1727) );
  HS65_LH_OAI21X2 U2405 ( .A(n17213), .B(n2552), .C(n1727), .Z(
        \u_DataPath/data_read_ex_1_i [6]) );
  HS65_LH_OAI21X2 U2428 ( .A(n37207), .B(n37251), .C(n1895), .Z(n1750) );
  HS65_LH_OAI21X2 U2429 ( .A(n17213), .B(n2576), .C(n1750), .Z(
        \u_DataPath/data_read_ex_1_i [5]) );
  HS65_LH_OAI21X2 U2452 ( .A(n38017), .B(n38015), .C(n1895), .Z(n1773) );
  HS65_LH_OAI21X2 U2453 ( .A(n17214), .B(n2600), .C(n1773), .Z(
        \u_DataPath/data_read_ex_1_i [4]) );
  HS65_LH_OAI21X2 U2476 ( .A(n38441), .B(n38443), .C(n1895), .Z(n1796) );
  HS65_LH_OAI21X2 U2477 ( .A(n17214), .B(n2624), .C(n1796), .Z(
        \u_DataPath/data_read_ex_1_i [3]) );
  HS65_LH_OAI21X2 U2500 ( .A(n38383), .B(n38430), .C(n1895), .Z(n1819) );
  HS65_LH_OAI21X2 U2501 ( .A(n17214), .B(n2648), .C(n1819), .Z(
        \u_DataPath/data_read_ex_1_i [2]) );
  HS65_LH_OAI21X2 U2524 ( .A(n37933), .B(n37937), .C(n1895), .Z(n1842) );
  HS65_LH_OAI21X2 U2525 ( .A(n17214), .B(n2672), .C(n1842), .Z(
        \u_DataPath/data_read_ex_1_i [1]) );
  HS65_LH_OAI21X2 U2548 ( .A(n34395), .B(n34392), .C(n1895), .Z(n1898) );
  HS65_LH_OAI21X2 U2549 ( .A(n17213), .B(n2729), .C(n1898), .Z(
        \u_DataPath/data_read_ex_1_i [0]) );
  HS65_LH_OAI21X2 U2623 ( .A(n36896), .B(n36955), .C(n2725), .Z(n1951) );
  HS65_LH_OAI21X2 U2647 ( .A(n36165), .B(n36162), .C(n2725), .Z(n1975) );
  HS65_LH_OAI21X2 U2671 ( .A(n35877), .B(n35876), .C(n2725), .Z(n1999) );
  HS65_LH_OAI21X2 U2695 ( .A(n35974), .B(n36004), .C(n2725), .Z(n2023) );
  HS65_LH_OAI21X2 U2719 ( .A(n35705), .B(n35703), .C(n2725), .Z(n2047) );
  HS65_LH_OAI21X2 U2743 ( .A(n36207), .B(n36206), .C(n2725), .Z(n2071) );
  HS65_LH_OAI21X2 U2767 ( .A(n36828), .B(n36821), .C(n2725), .Z(n2095) );
  HS65_LH_OAI21X2 U2791 ( .A(n35906), .B(n35908), .C(n2725), .Z(n2119) );
  HS65_LH_OAI21X2 U2815 ( .A(n36007), .B(n36039), .C(n2725), .Z(n2143) );
  HS65_LH_OAI21X2 U2839 ( .A(n36396), .B(n36395), .C(n2725), .Z(n2167) );
  HS65_LH_OAI21X2 U2863 ( .A(n35945), .B(n35941), .C(n2725), .Z(n2191) );
  HS65_LH_OAI21X2 U2887 ( .A(n36276), .B(n36272), .C(n2725), .Z(n2215) );
  HS65_LH_OAI21X2 U2911 ( .A(n35843), .B(n35845), .C(n2725), .Z(n2239) );
  HS65_LH_OAI21X2 U2935 ( .A(n36862), .B(n36863), .C(n2725), .Z(n2263) );
  HS65_LH_OAI21X2 U2959 ( .A(n36237), .B(n36271), .C(n2725), .Z(n2287) );
  HS65_LH_OAI21X2 U2983 ( .A(n35813), .B(n35814), .C(n2725), .Z(n2311) );
  HS65_LH_OAI21X2 U3007 ( .A(n36306), .B(n36305), .C(n2725), .Z(n2335) );
  HS65_LH_OAI21X2 U3031 ( .A(n31722), .B(n31716), .C(n2725), .Z(n2359) );
  HS65_LH_OAI21X2 U3055 ( .A(n36575), .B(n36573), .C(n2725), .Z(n2383) );
  HS65_LH_OAI21X2 U3079 ( .A(n36474), .B(n36427), .C(n2725), .Z(n2407) );
  HS65_LH_OAI21X2 U3103 ( .A(n36494), .B(n36484), .C(n2725), .Z(n2431) );
  HS65_LH_OAI21X2 U3127 ( .A(n36769), .B(n36768), .C(n2725), .Z(n2455) );
  HS65_LH_OAI21X2 U3151 ( .A(n36046), .B(n36054), .C(n2725), .Z(n2479) );
  HS65_LH_OAI21X2 U3175 ( .A(n36712), .B(n36757), .C(n2725), .Z(n2503) );
  HS65_LH_OAI21X2 U3199 ( .A(n36704), .B(n36657), .C(n2725), .Z(n2527) );
  HS65_LH_OAI21X2 U3223 ( .A(n35742), .B(n35737), .C(n2725), .Z(n2551) );
  HS65_LH_OAI21X2 U3247 ( .A(n36135), .B(n36127), .C(n2725), .Z(n2575) );
  HS65_LH_OAI21X2 U3271 ( .A(n33302), .B(n33331), .C(n2725), .Z(n2599) );
  HS65_LH_OAI21X2 U3295 ( .A(n33333), .B(n33363), .C(n2725), .Z(n2623) );
  HS65_LH_OAI21X2 U3319 ( .A(n35672), .B(n35702), .C(n2725), .Z(n2647) );
  HS65_LH_OAI21X2 U3343 ( .A(n34033), .B(n34047), .C(n2725), .Z(n2671) );
  HS65_LH_OAI21X2 U3367 ( .A(n32444), .B(n32441), .C(n2725), .Z(n2728) );
  HS65_LH_AND2X4 U3370 ( .A(n14109), .B(n2733), .Z(\u_DataPath/u_ifidreg/N35 )
         );
  HS65_LH_AND2X4 U3371 ( .A(n14105), .B(n2733), .Z(\u_DataPath/u_ifidreg/N34 )
         );
  HS65_LH_AND2X4 U3372 ( .A(n15469), .B(n2733), .Z(\u_DataPath/u_ifidreg/N33 )
         );
  HS65_LH_AND2X4 U3373 ( .A(n14103), .B(n2733), .Z(\u_DataPath/u_ifidreg/N32 )
         );
  HS65_LH_AND2X4 U3374 ( .A(n15466), .B(n2733), .Z(\u_DataPath/u_ifidreg/N31 )
         );
  HS65_LH_AND2X4 U3375 ( .A(n14101), .B(n2733), .Z(\u_DataPath/u_ifidreg/N30 )
         );
  HS65_LH_AND2X4 U3376 ( .A(n15463), .B(n2733), .Z(\u_DataPath/u_ifidreg/N29 )
         );
  HS65_LH_AND2X4 U3377 ( .A(n14099), .B(n2733), .Z(\u_DataPath/u_ifidreg/N28 )
         );
  HS65_LH_AND2X4 U3378 ( .A(n17714), .B(n2733), .Z(\u_DataPath/u_ifidreg/N27 )
         );
  HS65_LH_AND2X4 U3379 ( .A(n17716), .B(n2733), .Z(\u_DataPath/u_ifidreg/N26 )
         );
  HS65_LH_AND2X4 U3380 ( .A(n17718), .B(n2733), .Z(\u_DataPath/u_ifidreg/N25 )
         );
  HS65_LH_AND2X4 U3381 ( .A(n17720), .B(n2733), .Z(\u_DataPath/u_ifidreg/N24 )
         );
  HS65_LH_AND2X4 U3382 ( .A(n17722), .B(n2733), .Z(\u_DataPath/u_ifidreg/N23 )
         );
  HS65_LH_AND2X4 U3383 ( .A(n17656), .B(n2733), .Z(\u_DataPath/u_ifidreg/N22 )
         );
  HS65_LH_AND2X4 U3384 ( .A(n17658), .B(n2733), .Z(\u_DataPath/u_ifidreg/N21 )
         );
  HS65_LH_AND2X4 U3385 ( .A(n17661), .B(n2733), .Z(\u_DataPath/u_ifidreg/N20 )
         );
  HS65_LH_AND2X4 U3386 ( .A(n17662), .B(n2733), .Z(\u_DataPath/u_ifidreg/N19 )
         );
  HS65_LH_AND2X4 U3387 ( .A(n17665), .B(n2733), .Z(\u_DataPath/u_ifidreg/N18 )
         );
  HS65_LH_AND2X4 U3388 ( .A(n17666), .B(n2733), .Z(\u_DataPath/u_ifidreg/N17 )
         );
  HS65_LH_AND2X4 U3389 ( .A(n17669), .B(n2733), .Z(\u_DataPath/u_ifidreg/N16 )
         );
  HS65_LH_AND2X4 U3390 ( .A(n17670), .B(n2733), .Z(\u_DataPath/u_ifidreg/N15 )
         );
  HS65_LH_AND2X4 U3391 ( .A(n17673), .B(n2733), .Z(\u_DataPath/u_ifidreg/N14 )
         );
  HS65_LH_AND2X4 U3392 ( .A(n17674), .B(n2733), .Z(\u_DataPath/u_ifidreg/N13 )
         );
  HS65_LH_AND2X4 U3393 ( .A(n17677), .B(n2733), .Z(\u_DataPath/u_ifidreg/N12 )
         );
  HS65_LH_AND2X4 U3394 ( .A(n17678), .B(n2733), .Z(\u_DataPath/u_ifidreg/N11 )
         );
  HS65_LH_AND2X4 U3395 ( .A(n17680), .B(n2733), .Z(\u_DataPath/u_ifidreg/N10 )
         );
  HS65_LH_AND2X4 U3396 ( .A(n17682), .B(n2733), .Z(\u_DataPath/u_ifidreg/N9 )
         );
  HS65_LH_AND2X4 U3397 ( .A(n17685), .B(n2733), .Z(\u_DataPath/u_ifidreg/N8 )
         );
  HS65_LH_AND2X4 U3398 ( .A(n18021), .B(n2733), .Z(\u_DataPath/u_ifidreg/N7 )
         );
  HS65_LH_AND2X4 U3399 ( .A(n17687), .B(n2733), .Z(\u_DataPath/u_ifidreg/N6 )
         );
  HS65_LH_AND2X4 U3400 ( .A(n17689), .B(n2733), .Z(\u_DataPath/u_ifidreg/N5 )
         );
  HS65_LH_AND2X4 U3401 ( .A(n17691), .B(n2733), .Z(\u_DataPath/u_ifidreg/N4 )
         );
  HS65_LH_LDHQX4 \u_DataPath/u_execute/EXALU/ovf_reg  ( .G(
        \u_DataPath/u_execute/EXALU/N810 ), .D(
        \u_DataPath/u_execute/EXALU/N811 ), .Q(\u_DataPath/u_execute/ovf_i )
         );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][2]  ( 
        .G(rst), .D(\u_DataPath/u_decode_unit/reg_file0/N95 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][2] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][22]  ( 
        .G(rst), .D(\u_DataPath/u_decode_unit/reg_file0/N115 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][22] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][18]  ( 
        .G(rst), .D(\u_DataPath/u_decode_unit/reg_file0/N111 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][18] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][8]  ( 
        .G(rst), .D(\u_DataPath/u_decode_unit/reg_file0/N101 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][8] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][29]  ( 
        .G(rst), .D(\u_DataPath/u_decode_unit/reg_file0/N122 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][29] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][12]  ( 
        .G(rst), .D(\u_DataPath/u_decode_unit/reg_file0/N105 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][12] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][23]  ( 
        .G(rst), .D(\u_DataPath/u_decode_unit/reg_file0/N116 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][23] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][24]  ( 
        .G(rst), .D(\u_DataPath/u_decode_unit/reg_file0/N117 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][24] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][26]  ( 
        .G(rst), .D(\u_DataPath/u_decode_unit/reg_file0/N119 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][26] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][3]  ( 
        .G(rst), .D(\u_DataPath/u_decode_unit/reg_file0/N96 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][3] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][6]  ( 
        .G(rst), .D(\u_DataPath/u_decode_unit/reg_file0/N99 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][6] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][9]  ( 
        .G(rst), .D(\u_DataPath/u_decode_unit/reg_file0/N102 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][9] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][5]  ( 
        .G(rst), .D(\u_DataPath/u_decode_unit/reg_file0/N98 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][5] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][31]  ( 
        .G(rst), .D(\u_DataPath/u_decode_unit/reg_file0/N124 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][31] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][21]  ( 
        .G(rst), .D(\u_DataPath/u_decode_unit/reg_file0/N114 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][21] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][13]  ( 
        .G(rst), .D(\u_DataPath/u_decode_unit/reg_file0/N106 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][13] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][0]  ( 
        .G(rst), .D(\u_DataPath/u_decode_unit/reg_file0/N93 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][0] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][1]  ( 
        .G(rst), .D(\u_DataPath/u_decode_unit/reg_file0/N94 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][1] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][17]  ( 
        .G(rst), .D(\u_DataPath/u_decode_unit/reg_file0/N110 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][17] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][16]  ( 
        .G(rst), .D(\u_DataPath/u_decode_unit/reg_file0/N109 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][16] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][28]  ( 
        .G(rst), .D(\u_DataPath/u_decode_unit/reg_file0/N121 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][28] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][25]  ( 
        .G(rst), .D(\u_DataPath/u_decode_unit/reg_file0/N118 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][25] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][11]  ( 
        .G(rst), .D(\u_DataPath/u_decode_unit/reg_file0/N104 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][11] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][14]  ( 
        .G(rst), .D(\u_DataPath/u_decode_unit/reg_file0/N107 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][14] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][20]  ( 
        .G(rst), .D(\u_DataPath/u_decode_unit/reg_file0/N113 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][20] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][4]  ( 
        .G(rst), .D(\u_DataPath/u_decode_unit/reg_file0/N97 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][4] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][7]  ( 
        .G(rst), .D(\u_DataPath/u_decode_unit/reg_file0/N100 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][7] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][30]  ( 
        .G(rst), .D(\u_DataPath/u_decode_unit/reg_file0/N123 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][30] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][10]  ( 
        .G(rst), .D(\u_DataPath/u_decode_unit/reg_file0/N103 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][10] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][19]  ( 
        .G(rst), .D(\u_DataPath/u_decode_unit/reg_file0/N112 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][19] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][15]  ( 
        .G(rst), .D(\u_DataPath/u_decode_unit/reg_file0/N108 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][15] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][27]  ( 
        .G(rst), .D(\u_DataPath/u_decode_unit/reg_file0/N120 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][27] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N93 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][0] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N93 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][0] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N93 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][0] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N101 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][8] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N124 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][31] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N99 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][6] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N110 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][17] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N109 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][16] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N113 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][20] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N118 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][25] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N97 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][4] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N117 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][24] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N118 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][25] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N114 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][21] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N122 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][29] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N105 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][12] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N100 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][7] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N123 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][30] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N116 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][23] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N103 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][10] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N119 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][26] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N96 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][3] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N112 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][19] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N103 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][10] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N94 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][1] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N110 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][17] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N113 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][20] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N117 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][24] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N118 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][25] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N118 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][25] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N124 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][31] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N101 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][8] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N115 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][22] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N102 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][9] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N122 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][29] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N106 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][13] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N100 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][7] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N116 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][23] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N119 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][26] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N96 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][3] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N104 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][11] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N118 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][25] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N109 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][16] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N124 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][31] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N109 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][16] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N113 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][20] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N101 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][8] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N123 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][30] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N116 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][23] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N116 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][23] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N96 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][3] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N108 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][15] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N114 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][21] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N95 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][2] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N110 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][17] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N97 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][4] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N115 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][22] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N106 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][13] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N107 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][14] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N93 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][0] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N93 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][0] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N93 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][0] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N93 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][0] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N93 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][0] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N93 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][0] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N93 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][0] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N95 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][2] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N101 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][8] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N117 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][24] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N102 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][9] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N98 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][5] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N106 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][13] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N100 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][7] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N119 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][26] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N112 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][19] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N108 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][15] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N124 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][31] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N95 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][2] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N95 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][2] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N110 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][17] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N115 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][22] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N120 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][27] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N93 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][0] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N93 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][0] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N124 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][31] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N94 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][1] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N94 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][1] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N99 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][6] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N111 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][18] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N111 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][18] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N95 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][2] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N110 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][17] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N110 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][17] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N113 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][20] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N113 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][20] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N97 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][4] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N107 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][14] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N107 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][14] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N115 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][22] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N121 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][28] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N121 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][28] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N121 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][28] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N117 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][24] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N117 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][24] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N102 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][9] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N118 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][25] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N98 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][5] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N98 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][5] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N114 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][21] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N114 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][21] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N114 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][21] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N106 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][13] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N100 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][7] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N105 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][12] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N123 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][30] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N119 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][26] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N119 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][26] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N103 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][10] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N103 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][10] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N104 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][11] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N93 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][0] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N106 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][13] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N96 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][3] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N104 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][11] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N108 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][15] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N120 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][27] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N94 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][1] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N122 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][29] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N104 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][11] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N120 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][27] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N94 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][1] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N99 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][6] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N99 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][6] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N111 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][18] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N111 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][18] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N109 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][16] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N101 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][8] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N97 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][4] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N97 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][4] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N115 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][22] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N115 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][22] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N121 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][28] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N102 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][9] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N102 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][9] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N98 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][5] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N122 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][29] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N122 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][29] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N106 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][13] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N100 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][7] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N105 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][12] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N123 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][30] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N116 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][23] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N112 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][19] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N105 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][12] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N103 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][10] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N96 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][3] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N112 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][19] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N104 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][11] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N108 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][15] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N107 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][14] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N107 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][14] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N120 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][27] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N124 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][31] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N99 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][6] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N111 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][18] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N97 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][4] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N98 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][5] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N114 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][21] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N100 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][7] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N123 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][30] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N112 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][19] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N124 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][31] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N124 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][31] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N94 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][1] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N94 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][1] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N94 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][1] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N99 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][6] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N99 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][6] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N99 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][6] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N111 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][18] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N95 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][2] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N110 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][17] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N109 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][16] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N109 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][16] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N113 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][20] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N109 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][16] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N113 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][20] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N113 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][20] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N121 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][28] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N112 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][19] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N101 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][8] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N115 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][22] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N121 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][28] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N117 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][24] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N102 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][9] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N118 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][25] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N118 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][25] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N98 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][5] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N114 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][21] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N122 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][29] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N122 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][29] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N106 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][13] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N106 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][13] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N105 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][12] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N105 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][12] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N105 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][12] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N123 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][30] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N123 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][30] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N116 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][23] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N116 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][23] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N103 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][10] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N96 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][3] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N112 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][19] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N112 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][19] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N104 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][11] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N108 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][15] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N108 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][15] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N107 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][14] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N120 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][27] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N120 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][27] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N119 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][26] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N103 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][10] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N96 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][3] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N120 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][27] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N120 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][27] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N99 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][6] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N110 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][17] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N113 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][20] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N122 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][29] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N120 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][27] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N124 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][31] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N124 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][31] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N99 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][6] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N95 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][2] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N97 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][4] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N97 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][4] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N121 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][28] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N112 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][19] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N104 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][11] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N111 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][18] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N112 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][19] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N104 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][11] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N104 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][11] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N95 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][2] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N109 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][16] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N121 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][28] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N121 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][28] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N117 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][24] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N98 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][5] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N114 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][21] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N106 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][13] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N105 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][12] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N105 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][12] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N123 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][30] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N116 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][23] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N116 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][23] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N119 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][26] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N108 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][15] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N108 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][15] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N107 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][14] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N107 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][14] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N95 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][2] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N111 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][18] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N110 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][17] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N109 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][16] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N101 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][8] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N108 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][15] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N97 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][4] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N97 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][4] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N121 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][28] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N117 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][24] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N121 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][28] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N102 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][9] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N102 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][9] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N98 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][5] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N98 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][5] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N114 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][21] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N100 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][7] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N119 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][26] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N103 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][10] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N100 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][7] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N123 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][30] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N104 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][11] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N104 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][11] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N108 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][15] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N107 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][14] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N107 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][14] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N109 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][16] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N109 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][16] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N113 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][20] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N114 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][21] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N103 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][10] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N108 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][15] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N120 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][27] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N94 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][1] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N94 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][1] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N111 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][18] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N111 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][18] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N111 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][18] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N95 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][2] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N115 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][22] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N94 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][1] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N110 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][17] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N115 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][22] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N115 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][22] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N121 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][28] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N117 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][24] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N102 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][9] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N102 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][9] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N98 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][5] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N98 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][5] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N114 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][21] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N122 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][29] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N106 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][13] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N106 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][13] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N100 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][7] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N100 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][7] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N105 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][12] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N123 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][30] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N123 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][30] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N119 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][26] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N108 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][15] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N107 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][14] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N107 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][14] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N101 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][8] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N101 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][8] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N97 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][4] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N103 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][10] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N96 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][3] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N96 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][3] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N112 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][19] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N120 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][27] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N120 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][27] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N121 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][28] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N103 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][10] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N96 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][3] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N99 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][6] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N99 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][6] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N111 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][18] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N124 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][31] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N111 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][18] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N111 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][18] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N95 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][2] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N110 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][17] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N109 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][16] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N101 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][8] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N101 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][8] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N97 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][4] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N97 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][4] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N97 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][4] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N121 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][28] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N117 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][24] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N117 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][24] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N102 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][9] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N102 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][9] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N118 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][25] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N118 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][25] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N98 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][5] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N98 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][5] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N122 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][29] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N107 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][14] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N94 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][1] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N94 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][1] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N95 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][2] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N109 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][16] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N113 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][20] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N115 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][22] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N115 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][22] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N121 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][28] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N121 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][28] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N114 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][21] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N122 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][29] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N106 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][13] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N100 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][7] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N100 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][7] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N100 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][7] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N105 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][12] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N105 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][12] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N123 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][30] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N119 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][26] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N112 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][19] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N112 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][19] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N104 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][11] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N104 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][11] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N104 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][11] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N108 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][15] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N108 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][15] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N120 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][27] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N120 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][27] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N94 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][1] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N98 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][5] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N122 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][29] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N124 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][31] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N94 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][1] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N99 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][6] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N99 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][6] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N111 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][18] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N95 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][2] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N110 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][17] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N113 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][20] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N101 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][8] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N117 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][24] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N117 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][24] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N102 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][9] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N102 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][9] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N118 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][25] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N98 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][5] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N100 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][7] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N105 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][12] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N116 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][23] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N116 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][23] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N119 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][26] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N119 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][26] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N110 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][17] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N113 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][20] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N114 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][21] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N122 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][29] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N106 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][13] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N105 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][12] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N123 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][30] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N123 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][30] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N119 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][26] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N103 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][10] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N103 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][10] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N103 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][10] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N96 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][3] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N96 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][3] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N112 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][19] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N112 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][19] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N107 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][14] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N104 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][11] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N108 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][15] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N107 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][14] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N120 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][27] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N120 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][27] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N93 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][0] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N93 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][0] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N93 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N93 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N93 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N93 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N93 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N93 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N93 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N93 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N93 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N93 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N93 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N93 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N93 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N93 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N93 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][0] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N124 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][31] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N109 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][16] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N97 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][4] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N97 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][4] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N115 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][22] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N102 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][9] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N118 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][25] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N114 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][21] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N106 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][13] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N100 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][7] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N116 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][23] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N116 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][23] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N119 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][26] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N107 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][14] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N124 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][31] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N94 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N94 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N94 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][1] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N99 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][6] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N99 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N99 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][6] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N111 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N111 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N111 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][18] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N101 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][8] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N101 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][8] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N101 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][8] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N101 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N101 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N97 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N97 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][4] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N115 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][22] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N115 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][22] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N115 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N121 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][28] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N96 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][3] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N112 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N112 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N112 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][19] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N104 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N104 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][11] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N108 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N108 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N108 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N94 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][1] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N95 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][2] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N95 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][2] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N95 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N95 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][2] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N110 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][17] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N110 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][17] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N109 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][16] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N109 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][16] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N113 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][20] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N113 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][20] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N113 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N113 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N113 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N97 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N115 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N121 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N121 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][28] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N117 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][24] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N117 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][24] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N117 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][24] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N102 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N102 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N102 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][9] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N118 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][25] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N118 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][25] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N98 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N98 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N98 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N98 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][5] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N114 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][21] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N114 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N114 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][21] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N122 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][29] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N122 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][29] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N122 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N102 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][9] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N118 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][25] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N118 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N114 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N122 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][29] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N106 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][13] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N106 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][13] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N100 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N100 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N100 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][7] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N105 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][12] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N105 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N105 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][12] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N123 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][30] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N123 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N123 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N123 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N123 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][30] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N116 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][23] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N119 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][26] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N119 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N119 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][26] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N103 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][10] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N103 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N103 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N103 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N103 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][10] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N96 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][3] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N96 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][3] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N96 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][3] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N116 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N96 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N112 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N108 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N107 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N107 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N120 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N120 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N120 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N111 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][18] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N110 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N117 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N102 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N105 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N107 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][14] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N124 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][31] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N124 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N124 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N124 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N124 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N124 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N124 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N94 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N94 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N94 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N94 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N94 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N99 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N99 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N102 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N99 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N99 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N111 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N95 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N95 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N95 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N110 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N100 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N110 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N110 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N110 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N110 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N110 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N109 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N109 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N109 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N109 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N109 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N113 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N113 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N113 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N106 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N106 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N100 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N100 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N105 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][12] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N116 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N116 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N116 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N119 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N119 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N113 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N113 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N101 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N101 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N101 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N101 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N97 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N97 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N115 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N115 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N115 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N115 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N117 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N117 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N117 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N117 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N102 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N102 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N98 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N98 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N111 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N121 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N118 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N118 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N118 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N98 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N98 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N114 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N114 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N114 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N114 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N114 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N122 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N122 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N122 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N106 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N106 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N106 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N105 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N105 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N123 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N123 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N116 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N119 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N119 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N119 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N119 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N103 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N103 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N103 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N103 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N103 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N103 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N96 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N96 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N96 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N96 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N116 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N96 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N112 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N112 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N112 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N112 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N104 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N104 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N104 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N108 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N108 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N108 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N107 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N120 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N120 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N120 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N107 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N94 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N95 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N110 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N115 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N106 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N123 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N119 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N96 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N112 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N104 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N124 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N124 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N124 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N124 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N99 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N99 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N111 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N110 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N110 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N109 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N109 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N109 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N109 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N101 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N101 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N101 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N97 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N115 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N121 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N117 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N102 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N106 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N106 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N105 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N105 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N105 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N123 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N119 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N104 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N104 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N107 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N107 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N124 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N94 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N99 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N99 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N111 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N111 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N113 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N97 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N97 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N97 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N97 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N115 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N115 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N103 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N103 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N112 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N112 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N104 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N104 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N104 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N107 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N120 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N95 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N95 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N110 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N110 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N109 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N101 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N121 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N117 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N117 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N117 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N117 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N102 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N102 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N102 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N118 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N118 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N118 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N98 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N98 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N114 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N114 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N122 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N122 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N122 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N106 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N100 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N100 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N100 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N100 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N105 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N116 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N116 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N116 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N116 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N116 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N119 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N119 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N103 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N96 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N108 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N108 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N107 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N120 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N120 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N124 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N124 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N124 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N121 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N94 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N94 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N94 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N121 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N121 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N117 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N117 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N117 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N124 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N122 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N124 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N99 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N99 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N99 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N99 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N111 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N111 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N111 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N111 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N95 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N113 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N113 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N95 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N95 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N100 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N105 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N110 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N110 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N110 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N113 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N101 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N101 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N101 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N101 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N101 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N97 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N97 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N115 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N115 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N123 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N116 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N96 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N96 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N96 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N97 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N94 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N95 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N95 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N95 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N95 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N109 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N109 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N109 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N109 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N113 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N113 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N113 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N97 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N97 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N115 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N115 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N115 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N121 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N121 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N121 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N121 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N117 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N102 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N102 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N102 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N118 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N118 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N98 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N98 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N98 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N114 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N114 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N114 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N114 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N114 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N114 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N122 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N122 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N122 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N122 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N106 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N111 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N121 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N118 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N118 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N118 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N118 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N98 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N98 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N106 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N106 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N106 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N100 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N100 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N100 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N105 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N105 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N105 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N123 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N123 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N123 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N116 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N116 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N116 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N116 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N119 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N119 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N119 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N119 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N103 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N103 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N103 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N96 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N96 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N112 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N112 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N112 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N112 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N104 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N104 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N104 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N104 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N108 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N108 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N108 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N108 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N107 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N107 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N107 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N120 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N120 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][27] ) );
  HS65_LH_AOI21X2 U1586 ( .A(n17766), .B(n15578), .C(n1017), .Z(
        \u_DataPath/takeBranch_out_i ) );
  HS65_LH_AOI21X2 U637 ( .A(n34435), .B(n34441), .C(n284), .Z(n241) );
  HS65_LH_AOI21X2 U654 ( .A(n34431), .B(n31187), .C(n279), .Z(n272) );
  HS65_LH_NAND2X2 U1614 ( .A(n32806), .B(n1065), .Z(n1043) );
  HS65_LH_NAND2X2 U1617 ( .A(n32848), .B(n1065), .Z(n1046) );
  HS65_LH_NAND2X2 U1619 ( .A(n32925), .B(n1065), .Z(n1048) );
  HS65_LH_NAND2X2 U1627 ( .A(n33519), .B(n1065), .Z(n1056) );
  HS65_LH_NAND2X2 U1629 ( .A(n33558), .B(n1065), .Z(n1058) );
  HS65_LH_NAND2X2 U1625 ( .A(n33610), .B(n1065), .Z(n1054) );
  HS65_LH_NAND2X2 U590 ( .A(n189), .B(n35419), .Z(n253) );
  HS65_LH_AOI22X1 U1592 ( .A(n1065), .B(n35065), .C(n1040), .D(n35106), .Z(
        n1020) );
  HS65_LH_AOI22X1 U1599 ( .A(n1065), .B(n35108), .C(n1040), .D(n35111), .Z(
        n1027) );
  HS65_LH_AOI22X1 U1601 ( .A(n1065), .B(n35152), .C(n1040), .D(n35155), .Z(
        n1029) );
  HS65_LH_AOI22X1 U1605 ( .A(n1065), .B(n31868), .C(n1040), .D(n31874), .Z(
        n1033) );
  HS65_LH_AOI22X1 U1608 ( .A(n1065), .B(n32156), .C(n1040), .D(n32157), .Z(
        n1036) );
  HS65_LH_AOI22X1 U1612 ( .A(n1065), .B(n32628), .C(n1040), .D(n32697), .Z(
        n1041) );
  HS65_LH_NOR3X4 U746 ( .A(n33947), .B(n323), .C(n33942), .Z(n336) );
  HS65_LH_AOI22X1 U749 ( .A(n335), .B(Data_out_fromRAM[14]), .C(n336), .D(
        Data_out_fromRAM[30]), .Z(n314) );
  HS65_LH_NAND2X2 U750 ( .A(n314), .B(n320), .Z(
        \u_DataPath/from_mem_data_out_i [14]) );
  HS65_LH_AOI22X1 U761 ( .A(n335), .B(Data_out_fromRAM[8]), .C(n336), .D(
        Data_out_fromRAM[24]), .Z(n321) );
  HS65_LH_NAND2X2 U762 ( .A(n321), .B(n320), .Z(
        \u_DataPath/from_mem_data_out_i [8]) );
  HS65_LH_AOI22X1 U751 ( .A(n335), .B(Data_out_fromRAM[13]), .C(n336), .D(
        Data_out_fromRAM[29]), .Z(n315) );
  HS65_LH_NAND2X2 U752 ( .A(n315), .B(n320), .Z(
        \u_DataPath/from_mem_data_out_i [13]) );
  HS65_LH_AOI22X1 U757 ( .A(n335), .B(Data_out_fromRAM[10]), .C(n336), .D(
        Data_out_fromRAM[26]), .Z(n318) );
  HS65_LH_NAND2X2 U758 ( .A(n318), .B(n320), .Z(
        \u_DataPath/from_mem_data_out_i [10]) );
  HS65_LH_AOI22X1 U753 ( .A(n335), .B(Data_out_fromRAM[12]), .C(n336), .D(
        Data_out_fromRAM[28]), .Z(n316) );
  HS65_LH_NAND2X2 U754 ( .A(n316), .B(n320), .Z(
        \u_DataPath/from_mem_data_out_i [12]) );
  HS65_LH_AOI22X1 U747 ( .A(Data_out_fromRAM[15]), .B(n335), .C(
        Data_out_fromRAM[31]), .D(n336), .Z(n313) );
  HS65_LH_NAND2X2 U748 ( .A(n313), .B(n320), .Z(
        \u_DataPath/from_mem_data_out_i [15]) );
  HS65_LH_AOI22X1 U759 ( .A(n335), .B(Data_out_fromRAM[9]), .C(n336), .D(
        Data_out_fromRAM[25]), .Z(n319) );
  HS65_LH_NAND2X2 U760 ( .A(n319), .B(n320), .Z(
        \u_DataPath/from_mem_data_out_i [9]) );
  HS65_LH_AOI22X1 U755 ( .A(n335), .B(Data_out_fromRAM[11]), .C(n336), .D(
        Data_out_fromRAM[27]), .Z(n317) );
  HS65_LH_NAND2X2 U756 ( .A(n317), .B(n320), .Z(
        \u_DataPath/from_mem_data_out_i [11]) );
  HS65_LH_NOR2X2 U764 ( .A(n33943), .B(n323), .Z(n337) );
  HS65_LH_CNIVX3 U536 ( .A(n279), .Z(n189) );
  HS65_LH_NOR2X2 U534 ( .A(n279), .B(n35419), .Z(\u_DataPath/u_idexreg/N19 )
         );
  HS65_LH_NAND2X2 U601 ( .A(\u_DataPath/u_idexreg/N19 ), .B(n35216), .Z(n237)
         );
  HS65_LH_CNIVX3 U602 ( .A(n237), .Z(n244) );
  HS65_LH_NAND2X2 U545 ( .A(n189), .B(n31184), .Z(n257) );
  HS65_LH_NAND2X2 U548 ( .A(n189), .B(n31199), .Z(n190) );
  HS65_LH_NOR2X2 U596 ( .A(n31190), .B(n190), .Z(\u_DataPath/u_idexreg/N16 )
         );
  HS65_LH_NAND3X2 U541 ( .A(n189), .B(n35654), .C(n35263), .Z(n281) );
  HS65_LH_NOR3X1 U542 ( .A(n31180), .B(n35425), .C(n281), .Z(
        \u_DataPath/u_idexreg/N13 ) );
  HS65_LH_NOR2X2 U546 ( .A(n35425), .B(n257), .Z(n180) );
  HS65_LH_NOR2X2 U549 ( .A(n31182), .B(n190), .Z(\u_DataPath/u_idexreg/N11 )
         );
  HS65_LH_NOR3X1 U599 ( .A(\u_DataPath/u_idexreg/N16 ), .B(
        \u_DataPath/u_idexreg/N15 ), .C(\u_DataPath/u_idexreg/N10 ), .Z(n193)
         );
  HS65_LH_CBI4I1X3 U600 ( .A(n35220), .B(n35233), .C(n279), .D(n193), .Z(n227)
         );
  HS65_LH_OAI211X1 U629 ( .A(n34273), .B(n253), .C(n229), .D(n228), .Z(
        \u_DataPath/cw_to_ex_i [2]) );
  HS65_LH_CNIVX3 U591 ( .A(n253), .Z(n214) );
  HS65_LH_NOR3X1 U635 ( .A(n237), .B(n34596), .C(n34579), .Z(n246) );
  HS65_LH_CNIVX3 U640 ( .A(n246), .Z(n254) );
  HS65_LH_CNIVX3 U607 ( .A(\u_DataPath/u_idexreg/N19 ), .Z(n284) );
  HS65_LH_AOI312X2 U638 ( .A(n244), .B(n34432), .C(n34436), .D(n40525), .E(
        n246), .F(n241), .Z(n245) );
  HS65_LH_CBI4I6X2 U609 ( .A(n34700), .B(n237), .C(n201), .D(n34690), .Z(n215)
         );
  HS65_LH_AOI22X1 U620 ( .A(n34688), .B(n215), .C(n214), .D(n35029), .Z(n216)
         );
  HS65_LH_CBI4I1X3 U621 ( .A(n34701), .B(n34703), .C(n284), .D(n216), .Z(
        \u_DataPath/cw_to_ex_i [1]) );
  HS65_LH_NOR2X2 U649 ( .A(\u_DataPath/u_idexreg/N16 ), .B(
        \u_DataPath/u_idexreg/N15 ), .Z(n273) );
  HS65_LH_NAND2X2 U656 ( .A(n273), .B(n285), .Z(\u_DataPath/cw_to_ex_i [14])
         );
  HS65_LH_NOR3X1 U647 ( .A(n35425), .B(n33971), .C(n257), .Z(
        \u_DataPath/cw_exmem_i [4]) );
  HS65_LH_NOR3X1 U648 ( .A(n33973), .B(n35420), .C(n257), .Z(
        \u_DataPath/cw_exmem_i [6]) );
  HS65_LH_NOR2X6 U3369 ( .A(n37050), .B(n2731), .Z(\u_DataPath/u_idexreg/N184 ) );
  HS65_LH_NOR2X2 U644 ( .A(n33999), .B(n279), .Z(n255) );
  HS65_LH_NOR2X2 U663 ( .A(n283), .B(n34005), .Z(\u_DataPath/cw_to_ex_i [20])
         );
  HS65_LH_NOR2X6 U1669 ( .A(rst), .B(n39716), .Z(\u_DataPath/u_idexreg/N56 )
         );
  HS65_LH_CNIVX3 U1682 ( .A(n2731), .Z(\u_DataPath/u_idexreg/N40 ) );
  HS65_LH_IVX7 U493 ( .A(n2528), .Z(\u_DataPath/u_decode_unit/reg_file0/N100 )
         );
  HS65_LH_IVX7 U447 ( .A(n1976), .Z(\u_DataPath/u_decode_unit/reg_file0/N123 )
         );
  HS65_LH_IVX7 U457 ( .A(n2096), .Z(\u_DataPath/u_decode_unit/reg_file0/N118 )
         );
  HS65_LH_IVX7 U489 ( .A(n2480), .Z(\u_DataPath/u_decode_unit/reg_file0/N102 )
         );
  HS65_LH_IVX7 U481 ( .A(n2384), .Z(\u_DataPath/u_decode_unit/reg_file0/N106 )
         );
  HS65_LH_IVX7 U449 ( .A(n2000), .Z(\u_DataPath/u_decode_unit/reg_file0/N122 )
         );
  HS65_LH_IVX7 U483 ( .A(n2408), .Z(\u_DataPath/u_decode_unit/reg_file0/N105 )
         );
  HS65_LH_IVX7 U461 ( .A(n2144), .Z(\u_DataPath/u_decode_unit/reg_file0/N116 )
         );
  HS65_LH_IVX7 U491 ( .A(n2504), .Z(\u_DataPath/u_decode_unit/reg_file0/N101 )
         );
  HS65_LH_IVX7 U459 ( .A(n2120), .Z(\u_DataPath/u_decode_unit/reg_file0/N117 )
         );
  HS65_LH_IVX7 U463 ( .A(n2168), .Z(\u_DataPath/u_decode_unit/reg_file0/N115 )
         );
  HS65_LH_IVX7 U451 ( .A(n2024), .Z(\u_DataPath/u_decode_unit/reg_file0/N121 )
         );
  HS65_LH_IVX7 U467 ( .A(n2216), .Z(\u_DataPath/u_decode_unit/reg_file0/N113 )
         );
  HS65_LH_IVX7 U475 ( .A(n2312), .Z(\u_DataPath/u_decode_unit/reg_file0/N109 )
         );
  HS65_LH_IVX7 U473 ( .A(n2288), .Z(\u_DataPath/u_decode_unit/reg_file0/N110 )
         );
  HS65_LH_IVX7 U503 ( .A(n2648), .Z(\u_DataPath/u_decode_unit/reg_file0/N95 )
         );
  HS65_LH_IVX7 U505 ( .A(n2672), .Z(\u_DataPath/u_decode_unit/reg_file0/N94 )
         );
  HS65_LH_IVX7 U477 ( .A(n2336), .Z(\u_DataPath/u_decode_unit/reg_file0/N108 )
         );
  HS65_LH_IVX7 U485 ( .A(n2432), .Z(\u_DataPath/u_decode_unit/reg_file0/N104 )
         );
  HS65_LH_IVX7 U469 ( .A(n2240), .Z(\u_DataPath/u_decode_unit/reg_file0/N112 )
         );
  HS65_LH_IVX7 U471 ( .A(n2264), .Z(\u_DataPath/u_decode_unit/reg_file0/N111 )
         );
  HS65_LH_IVX7 U479 ( .A(n2360), .Z(\u_DataPath/u_decode_unit/reg_file0/N107 )
         );
  HS65_LH_IVX7 U453 ( .A(n2048), .Z(\u_DataPath/u_decode_unit/reg_file0/N120 )
         );
  HS65_LH_IVX7 U495 ( .A(n2552), .Z(\u_DataPath/u_decode_unit/reg_file0/N99 )
         );
  HS65_LH_IVX7 U445 ( .A(n1952), .Z(\u_DataPath/u_decode_unit/reg_file0/N124 )
         );
  HS65_LH_IVX7 U507 ( .A(n2729), .Z(\u_DataPath/u_decode_unit/reg_file0/N93 )
         );
  HS65_LH_NAND2X4 U228 ( .A(n100), .B(n17619), .Z(n99) );
  HS65_LH_NAND2X4 U253 ( .A(n106), .B(n17619), .Z(n104) );
  HS65_LH_NAND2X4 U262 ( .A(n17518), .B(n106), .Z(n113) );
  HS65_LH_NAND2X4 U243 ( .A(n17518), .B(n100), .Z(n101) );
  HS65_LH_OAI12X6 U261 ( .A(n17324), .B(n104), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N147 ) );
  HS65_LH_CNIVX3 U1589 ( .A(n1067), .Z(n1059) );
  HS65_LH_AND2X4 U848 ( .A(n36959), .B(n2733), .Z(\u_DataPath/u_exmemreg/N12 )
         );
  HS65_LH_OR2X4 U704 ( .A(n34069), .B(n323), .Z(n307) );
  HS65_LH_AND2X4 U893 ( .A(n15582), .B(n2733), .Z(
        \u_DataPath/branch_target_i [30]) );
  HS65_LH_AND2X4 U894 ( .A(n15584), .B(n2733), .Z(
        \u_DataPath/branch_target_i [29]) );
  HS65_LH_AND2X4 U895 ( .A(n15586), .B(n2733), .Z(
        \u_DataPath/branch_target_i [28]) );
  HS65_LH_AND2X4 U896 ( .A(n15588), .B(n2733), .Z(
        \u_DataPath/branch_target_i [27]) );
  HS65_LH_NOR3X4 U71 ( .A(rst), .B(n39558), .C(n38496), .Z(n69) );
  HS65_LH_NOR2X6 U70 ( .A(rst), .B(n31114), .Z(n68) );
  HS65_LH_AND2X4 U897 ( .A(n15590), .B(n2733), .Z(
        \u_DataPath/branch_target_i [26]) );
  HS65_LH_AND2X4 U898 ( .A(n15592), .B(n2733), .Z(
        \u_DataPath/branch_target_i [25]) );
  HS65_LH_AND2X4 U899 ( .A(n15594), .B(n2733), .Z(
        \u_DataPath/branch_target_i [24]) );
  HS65_LH_AOI22X1 U627 ( .A(\u_DataPath/u_idexreg/N19 ), .B(n34274), .C(n244), 
        .D(n34032), .Z(n229) );
  HS65_LH_NOR4ABX2 U598 ( .A(n31189), .B(n31188), .C(n279), .D(n31190), .Z(
        \u_DataPath/u_idexreg/N15 ) );
  HS65_LH_NOR2X6 U1803 ( .A(rst), .B(n40889), .Z(n1895) );
  HS65_LH_AND2X4 U900 ( .A(n15596), .B(n2733), .Z(
        \u_DataPath/branch_target_i [23]) );
  HS65_LH_OAI21X2 U3056 ( .A(n36822), .B(n2384), .C(n2383), .Z(
        \u_DataPath/data_read_ex_2_i [13]) );
  HS65_LH_OAI21X2 U3320 ( .A(n36924), .B(n2648), .C(n2647), .Z(
        \u_DataPath/data_read_ex_2_i [2]) );
  HS65_LH_OAI21X2 U3008 ( .A(n36822), .B(n2336), .C(n2335), .Z(
        \u_DataPath/data_read_ex_2_i [15]) );
  HS65_LH_OAI21X2 U3080 ( .A(n36822), .B(n2408), .C(n2407), .Z(
        \u_DataPath/data_read_ex_2_i [12]) );
  HS65_LH_OAI21X2 U3128 ( .A(n36822), .B(n2456), .C(n2455), .Z(
        \u_DataPath/data_read_ex_2_i [10]) );
  HS65_LH_OAI21X2 U3176 ( .A(n36822), .B(n2504), .C(n2503), .Z(
        \u_DataPath/data_read_ex_2_i [8]) );
  HS65_LH_OAI21X2 U3032 ( .A(n36895), .B(n2360), .C(n2359), .Z(
        \u_DataPath/data_read_ex_2_i [14]) );
  HS65_LH_OAI21X2 U3272 ( .A(n33304), .B(n2600), .C(n2599), .Z(
        \u_DataPath/data_read_ex_2_i [4]) );
  HS65_LH_OAI21X2 U3104 ( .A(n36822), .B(n2432), .C(n2431), .Z(
        \u_DataPath/data_read_ex_2_i [11]) );
  HS65_LH_OAI21X2 U3200 ( .A(n36822), .B(n2528), .C(n2527), .Z(
        \u_DataPath/data_read_ex_2_i [7]) );
  HS65_LH_OAI21X2 U3368 ( .A(n36895), .B(n2729), .C(n2728), .Z(
        \u_DataPath/data_read_ex_2_i [0]) );
  HS65_LH_OAI21X2 U3224 ( .A(n36924), .B(n2552), .C(n2551), .Z(
        \u_DataPath/data_read_ex_2_i [6]) );
  HS65_LH_OAI21X2 U3152 ( .A(n36924), .B(n2480), .C(n2479), .Z(
        \u_DataPath/data_read_ex_2_i [9]) );
  HS65_LH_OAI21X2 U3296 ( .A(n36924), .B(n2624), .C(n2623), .Z(
        \u_DataPath/data_read_ex_2_i [3]) );
  HS65_LH_OAI21X2 U3344 ( .A(n36917), .B(n2672), .C(n2671), .Z(
        \u_DataPath/data_read_ex_2_i [1]) );
  HS65_LH_OAI21X2 U3248 ( .A(n36924), .B(n2576), .C(n2575), .Z(
        \u_DataPath/data_read_ex_2_i [5]) );
  HS65_LH_OAI21X2 U2840 ( .A(n36822), .B(n2168), .C(n2167), .Z(
        \u_DataPath/data_read_ex_2_i [22]) );
  HS65_LH_OAI21X2 U2936 ( .A(n36924), .B(n2264), .C(n2263), .Z(
        \u_DataPath/data_read_ex_2_i [18]) );
  HS65_LH_OAI21X2 U2624 ( .A(n36924), .B(n1952), .C(n1951), .Z(
        \u_DataPath/data_read_ex_2_i [31]) );
  HS65_LH_OAI21X2 U2648 ( .A(n36164), .B(n1976), .C(n1975), .Z(
        \u_DataPath/data_read_ex_2_i [30]) );
  HS65_LH_OAI21X2 U2792 ( .A(n36164), .B(n2120), .C(n2119), .Z(
        \u_DataPath/data_read_ex_2_i [24]) );
  HS65_LH_OAI21X2 U2912 ( .A(n36164), .B(n2240), .C(n2239), .Z(
        \u_DataPath/data_read_ex_2_i [19]) );
  HS65_LH_OAI21X2 U2720 ( .A(n36164), .B(n2048), .C(n2047), .Z(
        \u_DataPath/data_read_ex_2_i [27]) );
  HS65_LH_OAI21X2 U2864 ( .A(n36924), .B(n2192), .C(n2191), .Z(
        \u_DataPath/data_read_ex_2_i [21]) );
  HS65_LH_OAI21X2 U2696 ( .A(n36924), .B(n2024), .C(n2023), .Z(
        \u_DataPath/data_read_ex_2_i [28]) );
  HS65_LH_OAI21X2 U2960 ( .A(n36924), .B(n2288), .C(n2287), .Z(
        \u_DataPath/data_read_ex_2_i [17]) );
  HS65_LH_OAI21X2 U2888 ( .A(n36924), .B(n2216), .C(n2215), .Z(
        \u_DataPath/data_read_ex_2_i [20]) );
  HS65_LH_OAI21X2 U2816 ( .A(n36822), .B(n2144), .C(n2143), .Z(
        \u_DataPath/data_read_ex_2_i [23]) );
  HS65_LH_OAI21X2 U2744 ( .A(n36924), .B(n2072), .C(n2071), .Z(
        \u_DataPath/data_read_ex_2_i [26]) );
  HS65_LH_OAI21X2 U2672 ( .A(n36924), .B(n2000), .C(n1999), .Z(
        \u_DataPath/data_read_ex_2_i [29]) );
  HS65_LH_OAI21X2 U2984 ( .A(n36924), .B(n2312), .C(n2311), .Z(
        \u_DataPath/data_read_ex_2_i [16]) );
  HS65_LH_OAI21X2 U2768 ( .A(n36822), .B(n2096), .C(n2095), .Z(
        \u_DataPath/data_read_ex_2_i [25]) );
  HS65_LH_OAI21X2 U639 ( .A(n34431), .B(n253), .C(n245), .Z(
        \u_DataPath/cw_to_ex_i [3]) );
  HS65_LH_NAND3X2 U608 ( .A(n34686), .B(\u_DataPath/u_idexreg/N19 ), .C(n34684), .Z(n201) );
  HS65_LH_AND2X4 U901 ( .A(n15598), .B(n2733), .Z(
        \u_DataPath/branch_target_i [22]) );
  HS65_LH_AND2X4 U902 ( .A(n15600), .B(n2733), .Z(
        \u_DataPath/branch_target_i [21]) );
  HS65_LH_AND2X4 U903 ( .A(n15602), .B(n2733), .Z(
        \u_DataPath/branch_target_i [20]) );
  HS65_LH_AND2X4 U152 ( .A(n17827), .B(n2733), .Z(n73) );
  HS65_LH_AND2X4 U904 ( .A(n15604), .B(n2733), .Z(
        \u_DataPath/branch_target_i [19]) );
  HS65_LH_AND2X4 U914 ( .A(n17752), .B(n2733), .Z(
        \u_DataPath/branch_target_i [9]) );
  HS65_LH_AND2X4 U915 ( .A(n17751), .B(n2733), .Z(
        \u_DataPath/branch_target_i [8]) );
  HS65_LH_AND2X4 U908 ( .A(n15612), .B(n2733), .Z(
        \u_DataPath/branch_target_i [15]) );
  HS65_LH_AND2X4 U920 ( .A(n17746), .B(n2733), .Z(
        \u_DataPath/branch_target_i [3]) );
  HS65_LH_AND2X4 U909 ( .A(n15614), .B(n2733), .Z(
        \u_DataPath/branch_target_i [14]) );
  HS65_LH_AND2X4 U913 ( .A(n15622), .B(n2733), .Z(
        \u_DataPath/branch_target_i [10]) );
  HS65_LH_AND2X4 U905 ( .A(n15606), .B(n2733), .Z(
        \u_DataPath/branch_target_i [18]) );
  HS65_LH_AND2X4 U922 ( .A(n34015), .B(n2733), .Z(
        \u_DataPath/branch_target_i [1]) );
  HS65_LH_AND2X4 U911 ( .A(n15618), .B(n2733), .Z(
        \u_DataPath/branch_target_i [12]) );
  HS65_LH_AND2X4 U910 ( .A(n15616), .B(n2733), .Z(
        \u_DataPath/branch_target_i [13]) );
  HS65_LH_AND2X4 U912 ( .A(n15620), .B(n2733), .Z(
        \u_DataPath/branch_target_i [11]) );
  HS65_LH_AND2X4 U907 ( .A(n15610), .B(n2733), .Z(
        \u_DataPath/branch_target_i [16]) );
  HS65_LH_AND2X4 U919 ( .A(n17747), .B(n2733), .Z(
        \u_DataPath/branch_target_i [4]) );
  HS65_LH_AND2X4 U906 ( .A(n15608), .B(n2733), .Z(
        \u_DataPath/branch_target_i [17]) );
  HS65_LH_AND2X4 U917 ( .A(n17749), .B(n2733), .Z(
        \u_DataPath/branch_target_i [6]) );
  HS65_LH_AND2X4 U916 ( .A(n17750), .B(n2733), .Z(
        \u_DataPath/branch_target_i [7]) );
  HS65_LH_AND2X4 U918 ( .A(n17748), .B(n2733), .Z(
        \u_DataPath/branch_target_i [5]) );
  HS65_LH_AND2X4 U921 ( .A(n17745), .B(n2733), .Z(
        \u_DataPath/branch_target_i [2]) );
  HS65_LH_NOR3X4 U1588 ( .A(n40653), .B(n40712), .C(n1019), .Z(n1067) );
  HS65_LH_NOR3AX4 U1590 ( .A(\u_DataPath/u_exmemreg/N12 ), .B(n40652), .C(
        n40562), .Z(n1065) );
  HS65_LH_NOR2AX3 U1591 ( .A(n40561), .B(n1019), .Z(n1040) );
  HS65_LH_NOR2X6 U69 ( .A(rst), .B(n10452), .Z(n70) );
  HS65_LH_OAI112X11 U439 ( .A(n39446), .B(n39445), .C(n39444), .D(n2733), .Z(
        \u_DataPath/u_fetch/pc1/N3 ) );
  HS65_LH_NOR3X1 U705 ( .A(n34051), .B(n34175), .C(n323), .Z(n309) );
  HS65_LH_NAND4ABX3 U712 ( .A(n34054), .B(n34055), .C(n309), .D(n34052), .Z(
        n320) );
  HS65_LH_NOR2X6 U858 ( .A(rst), .B(n17771), .Z(n348) );
  HS65_LH_AND2X4 U859 ( .A(n17770), .B(n2733), .Z(n347) );
  HS65_LH_NOR2X2 U646 ( .A(n17692), .B(n283), .Z(\u_DataPath/cw_exmem_i [1])
         );
  HS65_LH_NOR2X2 U622 ( .A(n34272), .B(n257), .Z(\u_DataPath/u_idexreg/N8 ) );
  HS65_LH_AND2X4 U2622 ( .A(n36920), .B(n2733), .Z(n2725) );
  HS65_LH_NOR2X2 U661 ( .A(n34351), .B(n281), .Z(\u_DataPath/u_idexreg/N21 )
         );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N93 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][0] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N121 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][28] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N100 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][7] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N107 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][14] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N99 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][6] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N111 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][18] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N105 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][12] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N123 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][30] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N104 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][11] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N107 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][14] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N94 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][1] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N95 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][2] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N110 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][17] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N109 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][16] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N101 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][8] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N115 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][22] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N117 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][24] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N102 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][9] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N118 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][25] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N122 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][29] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N106 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][13] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N106 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][13] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N100 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][7] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N123 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][30] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N116 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][23] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N120 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][27] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N120 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][27] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N107 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][14] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N113 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][20] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N123 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][30] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N99 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][6] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N118 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][25] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N105 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][12] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N112 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][19] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N108 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][15] ) );
  HS65_LH_NOR3X3 U227 ( .A(rst), .B(n17628), .C(n17279), .Z(n100) );
  HS65_LH_NOR3X3 U252 ( .A(rst), .B(n17507), .C(n17279), .Z(n106) );
  HS65_LH_OR2X4 U1587 ( .A(n40652), .B(rst), .Z(n1019) );
  HS65_LH_NAND2X5 U703 ( .A(n34060), .B(n2733), .Z(n323) );
  HS65_LH_CBI4I6X2 U443 ( .A(n39473), .B(n34377), .C(n34378), .D(rst), .Z(
        \u_DataPath/u_decode_unit/hdu_0/current_state [0]) );
  HS65_LH_NAND2X5 U530 ( .A(n2733), .B(n35215), .Z(n279) );
  HS65_LH_AOI211X2 U655 ( .A(n37052), .B(n2733), .C(n272), .D(
        \u_DataPath/u_idexreg/N10 ), .Z(n285) );
  HS65_LH_OAI21X2 U1585 ( .A(n17764), .B(n15578), .C(n18159), .Z(n1017) );
  HS65_LH_NOR2X2 U845 ( .A(rst), .B(n40603), .Z(
        \u_DataPath/regfile_addr_out_towb_i [1]) );
  HS65_LH_NOR2X2 U844 ( .A(rst), .B(n40604), .Z(
        \u_DataPath/regfile_addr_out_towb_i [2]) );
  HS65_LH_NOR2X2 U843 ( .A(rst), .B(n40475), .Z(
        \u_DataPath/regfile_addr_out_towb_i [3]) );
  HS65_LH_NOR2X2 U841 ( .A(rst), .B(n33889), .Z(
        \u_DataPath/from_alu_data_out_i [0]) );
  HS65_LH_NAND2X4 U1681 ( .A(n39672), .B(n2733), .Z(n2731) );
  HS65_LH_NOR2X2 U842 ( .A(rst), .B(n40226), .Z(
        \u_DataPath/regfile_addr_out_towb_i [4]) );
  HS65_LH_NOR2X2 U846 ( .A(rst), .B(n40607), .Z(
        \u_DataPath/regfile_addr_out_towb_i [0]) );
  HS65_LH_NOR2X2 U840 ( .A(rst), .B(n33910), .Z(
        \u_DataPath/from_alu_data_out_i [1]) );
  HS65_LH_NOR2X2 U517 ( .A(rst), .B(n17853), .Z(
        \u_DataPath/u_execute/psw_status_i [0]) );
  HS65_LH_NOR2X2 U1638 ( .A(rst), .B(n32120), .Z(
        \u_DataPath/mem_writedata_out_i [30]) );
  HS65_LH_NOR2X2 U1642 ( .A(rst), .B(n32212), .Z(
        \u_DataPath/mem_writedata_out_i [26]) );
  HS65_LH_NOR2X2 U1662 ( .A(rst), .B(n31930), .Z(
        \u_DataPath/mem_writedata_out_i [6]) );
  HS65_LH_NOR2X2 U1643 ( .A(rst), .B(n32234), .Z(
        \u_DataPath/mem_writedata_out_i [25]) );
  HS65_LH_NOR2X2 U1667 ( .A(rst), .B(n31994), .Z(
        \u_DataPath/mem_writedata_out_i [1]) );
  HS65_LH_NOR2X2 U1668 ( .A(rst), .B(n32057), .Z(
        \u_DataPath/mem_writedata_out_i [0]) );
  HS65_LH_NOR2X2 U1644 ( .A(rst), .B(n32256), .Z(
        \u_DataPath/mem_writedata_out_i [24]) );
  HS65_LH_NOR2X2 U1648 ( .A(rst), .B(n31613), .Z(
        \u_DataPath/mem_writedata_out_i [20]) );
  HS65_LH_NOR2X2 U1649 ( .A(rst), .B(n31634), .Z(
        \u_DataPath/mem_writedata_out_i [19]) );
  HS65_LH_NOR2X2 U1647 ( .A(rst), .B(n31593), .Z(
        \u_DataPath/mem_writedata_out_i [21]) );
  HS65_LH_NOR2X2 U1660 ( .A(rst), .B(n31438), .Z(
        \u_DataPath/mem_writedata_out_i [8]) );
  HS65_LH_NOR2X2 U1664 ( .A(rst), .B(n32014), .Z(
        \u_DataPath/mem_writedata_out_i [4]) );
  HS65_LH_NOR2X2 U1665 ( .A(rst), .B(n32036), .Z(
        \u_DataPath/mem_writedata_out_i [3]) );
  HS65_LH_NOR2X2 U1654 ( .A(rst), .B(n31457), .Z(
        \u_DataPath/mem_writedata_out_i [14]) );
  HS65_LH_NOR2X2 U1656 ( .A(rst), .B(n31496), .Z(
        \u_DataPath/mem_writedata_out_i [12]) );
  HS65_LH_NOR2X2 U1652 ( .A(rst), .B(n31695), .Z(
        \u_DataPath/mem_writedata_out_i [16]) );
  HS65_LH_NOR2X2 U1657 ( .A(rst), .B(n31553), .Z(
        \u_DataPath/mem_writedata_out_i [11]) );
  HS65_LH_NOR2X2 U1663 ( .A(rst), .B(n31951), .Z(
        \u_DataPath/mem_writedata_out_i [5]) );
  HS65_LH_NOR2X2 U1639 ( .A(rst), .B(n32099), .Z(
        \u_DataPath/mem_writedata_out_i [29]) );
  HS65_LH_NOR2X2 U1655 ( .A(rst), .B(n31477), .Z(
        \u_DataPath/mem_writedata_out_i [13]) );
  HS65_LH_NOR2X2 U1651 ( .A(rst), .B(n31675), .Z(
        \u_DataPath/mem_writedata_out_i [17]) );
  HS65_LH_NOR2X2 U1661 ( .A(rst), .B(n31744), .Z(
        \u_DataPath/mem_writedata_out_i [7]) );
  HS65_LH_NOR2X2 U1658 ( .A(rst), .B(n31419), .Z(
        \u_DataPath/mem_writedata_out_i [10]) );
  HS65_LH_NOR2X2 U1650 ( .A(rst), .B(n31654), .Z(
        \u_DataPath/mem_writedata_out_i [18]) );
  HS65_LH_NOR2X2 U442 ( .A(rst), .B(n37036), .Z(
        \u_DataPath/u_decode_unit/hdu_0/current_state [1]) );
  HS65_LH_NOR2X2 U1645 ( .A(rst), .B(n32277), .Z(
        \u_DataPath/mem_writedata_out_i [23]) );
  HS65_LH_NOR2X2 U1646 ( .A(rst), .B(n31572), .Z(
        \u_DataPath/mem_writedata_out_i [22]) );
  HS65_LH_NOR2X2 U1641 ( .A(rst), .B(n32300), .Z(
        \u_DataPath/mem_writedata_out_i [27]) );
  HS65_LH_NOR2X2 U1659 ( .A(rst), .B(n31515), .Z(
        \u_DataPath/mem_writedata_out_i [9]) );
  HS65_LH_NOR2X2 U1653 ( .A(rst), .B(n31534), .Z(
        \u_DataPath/mem_writedata_out_i [15]) );
  HS65_LH_NOR2X2 U1640 ( .A(rst), .B(n32342), .Z(
        \u_DataPath/mem_writedata_out_i [28]) );
  HS65_LH_NOR2X2 U1637 ( .A(rst), .B(n32323), .Z(
        \u_DataPath/mem_writedata_out_i [31]) );
  HS65_LH_IVX7 U465 ( .A(n2192), .Z(\u_DataPath/u_decode_unit/reg_file0/N114 )
         );
  HS65_LH_IVX7 U487 ( .A(n2456), .Z(\u_DataPath/u_decode_unit/reg_file0/N103 )
         );
  HS65_LH_IVX7 U497 ( .A(n2576), .Z(\u_DataPath/u_decode_unit/reg_file0/N98 )
         );
  HS65_LH_IVX7 U499 ( .A(n2600), .Z(\u_DataPath/u_decode_unit/reg_file0/N97 )
         );
  HS65_LH_IVX7 U455 ( .A(n2072), .Z(\u_DataPath/u_decode_unit/reg_file0/N119 )
         );
  HS65_LH_IVX7 U501 ( .A(n2624), .Z(\u_DataPath/u_decode_unit/reg_file0/N96 )
         );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N118 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][25] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N123 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][30] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N108 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][15] ) );
  HS65_LL_IVX18 U3434 ( .A(n14001), .Z(addr_to_iram_1) );
  HS65_LL_IVX18 U3435 ( .A(n14010), .Z(read_op_snps_wire) );
  HS65_LL_IVX18 U3436 ( .A(n13925), .Z(\Address_toRAM[10]_snps_wire ) );
  HS65_LL_IVX18 U3437 ( .A(n13927), .Z(\Address_toRAM[7]_snps_wire ) );
  HS65_LL_IVX18 U3438 ( .A(n13929), .Z(\Address_toRAM[11]_snps_wire ) );
  HS65_LL_IVX18 U3439 ( .A(n13931), .Z(\Address_toRAM[9]_snps_wire ) );
  HS65_LL_IVX18 U3440 ( .A(n13933), .Z(\Address_toRAM[4]_snps_wire ) );
  HS65_LL_IVX18 U3441 ( .A(n13935), .Z(\Address_toRAM[6]_snps_wire ) );
  HS65_LL_IVX18 U3442 ( .A(n13937), .Z(\Address_toRAM[2]_snps_wire ) );
  HS65_LL_IVX18 U3443 ( .A(n13939), .Z(\Address_toRAM[5]_snps_wire ) );
  HS65_LL_IVX18 U3444 ( .A(n14012), .Z(\Data_in[22]_snps_wire ) );
  HS65_LL_IVX18 U3445 ( .A(n14014), .Z(\Data_in[21]_snps_wire ) );
  HS65_LL_IVX18 U3446 ( .A(n14016), .Z(\Data_in[20]_snps_wire ) );
  HS65_LL_IVX18 U3447 ( .A(n14018), .Z(\Data_in[19]_snps_wire ) );
  HS65_LL_IVX18 U3448 ( .A(n14020), .Z(\Data_in[18]_snps_wire ) );
  HS65_LL_IVX18 U3449 ( .A(n14022), .Z(\Data_in[17]_snps_wire ) );
  HS65_LL_IVX18 U3450 ( .A(n14024), .Z(\Data_in[16]_snps_wire ) );
  HS65_LL_IVX18 U3451 ( .A(n13921), .Z(\Data_in[30]_snps_wire ) );
  HS65_LL_IVX18 U3452 ( .A(n13923), .Z(\Data_in[29]_snps_wire ) );
  HS65_LL_IVX18 U3453 ( .A(n13941), .Z(\Address_toRAM[3]_snps_wire ) );
  HS65_LL_IVX18 U3454 ( .A(n14008), .Z(\Data_in[7]_snps_wire ) );
  HS65_LL_IVX18 U3455 ( .A(n13905), .Z(\Data_in[15]_snps_wire ) );
  HS65_LL_IVX18 U3456 ( .A(n13907), .Z(\Data_in[14]_snps_wire ) );
  HS65_LL_IVX18 U3457 ( .A(n13909), .Z(\Data_in[9]_snps_wire ) );
  HS65_LL_IVX18 U3458 ( .A(n13911), .Z(\Data_in[11]_snps_wire ) );
  HS65_LL_IVX18 U3459 ( .A(n13913), .Z(\Data_in[10]_snps_wire ) );
  HS65_LL_IVX18 U3460 ( .A(n13915), .Z(\Data_in[8]_snps_wire ) );
  HS65_LL_IVX18 U3461 ( .A(n13917), .Z(\Data_in[13]_snps_wire ) );
  HS65_LL_IVX18 U3462 ( .A(n13919), .Z(\Data_in[12]_snps_wire ) );
  HS65_LL_NAND3X2 U3463 ( .A(\u_DataPath/regfile_addr_out_towb_i [2]), .B(
        n15714), .C(n15712), .Z(n109) );
  HS65_LH_IVX9 U3464 ( .A(n15665), .Z(n13921) );
  HS65_LH_IVX9 U3465 ( .A(n15664), .Z(n13923) );
  HS65_LH_IVX9 U3466 ( .A(n15671), .Z(n14008) );
  HS65_LH_IVX9 U3467 ( .A(n15661), .Z(n13925) );
  HS65_LH_IVX9 U3468 ( .A(n15657), .Z(n13927) );
  HS65_LH_IVX9 U3469 ( .A(n15645), .Z(n13929) );
  HS65_LH_IVX9 U3470 ( .A(n15655), .Z(n13931) );
  HS65_LH_IVX9 U3471 ( .A(n15653), .Z(n13933) );
  HS65_LH_IVX9 U3472 ( .A(n15647), .Z(n13935) );
  HS65_LH_IVX9 U3473 ( .A(n15659), .Z(n13937) );
  HS65_LH_IVX9 U3474 ( .A(n15649), .Z(n13939) );
  HS65_LH_IVX9 U3475 ( .A(n15676), .Z(n13905) );
  HS65_LH_IVX9 U3476 ( .A(n15684), .Z(n13907) );
  HS65_LH_IVX9 U3477 ( .A(n15678), .Z(n13909) );
  HS65_LH_IVX9 U3478 ( .A(n15673), .Z(n13911) );
  HS65_LH_IVX9 U3479 ( .A(n15689), .Z(n13913) );
  HS65_LH_IVX9 U3480 ( .A(n15686), .Z(n13915) );
  HS65_LH_IVX9 U3481 ( .A(n15682), .Z(n13917) );
  HS65_LH_IVX9 U3482 ( .A(n15680), .Z(n13919) );
  HS65_LH_AND2X4 U3483 ( .A(\u_DataPath/mem_writedata_out_i [7]), .B(
        write_op_snps_wire), .Z(n15671) );
  HS65_LH_NOR2X3 U3484 ( .A(n15700), .B(n15650), .Z(n15651) );
  HS65_LH_NOR2AX3 U3485 ( .A(\u_DataPath/mem_writedata_out_i [30]), .B(n14072), 
        .Z(n15665) );
  HS65_LH_NOR2AX3 U3486 ( .A(\u_DataPath/mem_writedata_out_i [29]), .B(n14072), 
        .Z(n15664) );
  HS65_LH_BFX9 U3487 ( .A(n15675), .Z(n15676) );
  HS65_LH_BFX9 U3488 ( .A(n15683), .Z(n15684) );
  HS65_LH_BFX9 U3489 ( .A(n15677), .Z(n15678) );
  HS65_LH_BFX9 U3490 ( .A(n15672), .Z(n15673) );
  HS65_LH_BFX9 U3491 ( .A(n15688), .Z(n15689) );
  HS65_LH_BFX9 U3492 ( .A(n15685), .Z(n15686) );
  HS65_LH_BFX9 U3493 ( .A(n15681), .Z(n15682) );
  HS65_LH_BFX9 U3494 ( .A(n15679), .Z(n15680) );
  HS65_LH_OAI211X1 U3495 ( .A(n15704), .B(n15703), .C(n15702), .D(n15701), .Z(
        n15705) );
  HS65_LH_NOR2AX3 U3496 ( .A(\u_DataPath/mem_writedata_out_i [16]), .B(n15694), 
        .Z(n15691) );
  HS65_LH_NOR2AX3 U3497 ( .A(\u_DataPath/mem_writedata_out_i [17]), .B(n15694), 
        .Z(n15695) );
  HS65_LH_NOR2AX3 U3498 ( .A(\u_DataPath/mem_writedata_out_i [18]), .B(n15694), 
        .Z(n15693) );
  HS65_LH_NOR2AX3 U3499 ( .A(\u_DataPath/mem_writedata_out_i [19]), .B(n15694), 
        .Z(n15690) );
  HS65_LH_NOR2AX3 U3500 ( .A(\u_DataPath/mem_writedata_out_i [20]), .B(n15694), 
        .Z(n15687) );
  HS65_LH_NOR2AX3 U3501 ( .A(\u_DataPath/mem_writedata_out_i [21]), .B(n15694), 
        .Z(n15692) );
  HS65_LH_NOR2AX3 U3502 ( .A(\u_DataPath/mem_writedata_out_i [22]), .B(n15694), 
        .Z(n15674) );
  HS65_LL_NOR2X6 U3503 ( .A(n15706), .B(n15185), .Z(n14078) );
  HS65_LL_IVX18 U3504 ( .A(n13893), .Z(\nibble[0]_snps_wire ) );
  HS65_LH_IVX9 U3505 ( .A(n13897), .Z(n13898) );
  HS65_LH_IVX9 U3506 ( .A(n13901), .Z(n13902) );
  HS65_LH_IVX9 U3507 ( .A(n13943), .Z(n13944) );
  HS65_LH_IVX9 U3508 ( .A(n13895), .Z(n13896) );
  HS65_LH_IVX9 U3509 ( .A(n13899), .Z(n13900) );
  HS65_LH_IVX9 U3510 ( .A(n13903), .Z(n13904) );
  HS65_LH_IVX9 U3511 ( .A(n16341), .Z(n13901) );
  HS65_LH_IVX9 U3512 ( .A(n17164), .Z(n13903) );
  HS65_LH_IVX9 U3513 ( .A(n17091), .Z(n13943) );
  HS65_LH_IVX9 U3514 ( .A(n16460), .Z(n13897) );
  HS65_LH_IVX9 U3515 ( .A(n14026), .Z(n14027) );
  HS65_LH_IVX9 U3516 ( .A(n16399), .Z(n13899) );
  HS65_LH_IVX9 U3517 ( .A(n16359), .Z(n13895) );
  HS65_LH_IVX9 U3518 ( .A(n14071), .Z(n14026) );
  HS65_LH_AOI21X2 U3519 ( .A(n15696), .B(n9305), .C(n14070), .Z(n14071) );
  HS65_LH_IVX4 U3520 ( .A(n4239), .Z(n14002) );
  HS65_LL_IVX18 U3522 ( .A(n13973), .Z(addr_to_iram_29) );
  HS65_LH_AOI21X2 U3523 ( .A(n15049), .B(n15217), .C(n15048), .Z(n15050) );
  HS65_LH_NOR2X2 U3524 ( .A(n10585), .B(n10589), .Z(n14069) );
  HS65_LL_IVX18 U3525 ( .A(n13997), .Z(addr_to_iram_28) );
  HS65_LL_IVX18 U3526 ( .A(n13999), .Z(addr_to_iram_26) );
  HS65_LL_IVX18 U3527 ( .A(n13969), .Z(addr_to_iram_27) );
  HS65_LL_IVX18 U3528 ( .A(n13993), .Z(addr_to_iram_24) );
  HS65_LL_IVX18 U3529 ( .A(n13967), .Z(addr_to_iram_25) );
  HS65_LL_IVX18 U3530 ( .A(n13995), .Z(addr_to_iram_22) );
  HS65_LL_IVX18 U3531 ( .A(n13965), .Z(addr_to_iram_23) );
  HS65_LL_IVX18 U3532 ( .A(n13989), .Z(addr_to_iram_20) );
  HS65_LL_IVX18 U3533 ( .A(n13963), .Z(addr_to_iram_21) );
  HS65_LL_IVX18 U3534 ( .A(n13991), .Z(addr_to_iram_18) );
  HS65_LL_IVX18 U3535 ( .A(n13961), .Z(addr_to_iram_19) );
  HS65_LL_IVX18 U3536 ( .A(n13985), .Z(addr_to_iram_16) );
  HS65_LL_IVX18 U3537 ( .A(n13959), .Z(addr_to_iram_17) );
  HS65_LL_IVX18 U3538 ( .A(n13987), .Z(addr_to_iram_14) );
  HS65_LL_IVX18 U3539 ( .A(n13957), .Z(addr_to_iram_15) );
  HS65_LL_IVX18 U3540 ( .A(n13981), .Z(addr_to_iram_12) );
  HS65_LL_IVX18 U3541 ( .A(n13955), .Z(addr_to_iram_13) );
  HS65_LL_NAND2X2 U3543 ( .A(n14244), .B(n15501), .Z(n15411) );
  HS65_LL_IVX18 U3544 ( .A(n13983), .Z(addr_to_iram_10) );
  HS65_LL_IVX18 U3545 ( .A(n13953), .Z(addr_to_iram_11) );
  HS65_LL_IVX18 U3547 ( .A(n13977), .Z(addr_to_iram_8) );
  HS65_LL_IVX18 U3548 ( .A(n13951), .Z(addr_to_iram_9) );
  HS65_LL_IVX18 U3549 ( .A(n13979), .Z(addr_to_iram_6) );
  HS65_LL_IVX18 U3550 ( .A(n13949), .Z(addr_to_iram_7) );
  HS65_LL_IVX18 U3551 ( .A(n13947), .Z(addr_to_iram_5) );
  HS65_LL_IVX18 U3552 ( .A(n13971), .Z(addr_to_iram_4) );
  HS65_LL_IVX18 U3553 ( .A(n13975), .Z(addr_to_iram_2) );
  HS65_LH_CNIVX3 U3554 ( .A(n14005), .Z(n14006) );
  HS65_LH_IVX9 U3555 ( .A(n4239), .Z(n14004) );
  HS65_LL_IVX18 U3556 ( .A(n13945), .Z(addr_to_iram_3) );
  HS65_LH_IVX9 U3557 ( .A(n4236), .Z(n14001) );
  HS65_LH_CNIVX3 U3558 ( .A(\u_DataPath/idex_rt_i [2]), .Z(n9794) );
  HS65_LH_CNIVX3 U3559 ( .A(\u_DataPath/idex_rt_i [0]), .Z(n9641) );
  HS65_LH_BFX4 U3560 ( .A(n2775), .Z(n2773) );
  HS65_LH_BFX4 U3561 ( .A(n2776), .Z(n2774) );
  HS65_LH_BFX4 U3562 ( .A(n2777), .Z(n2775) );
  HS65_LH_BFX4 U3563 ( .A(n2778), .Z(n2776) );
  HS65_LH_BFX4 U3564 ( .A(n2779), .Z(n2777) );
  HS65_LH_BFX4 U3565 ( .A(n2780), .Z(n2778) );
  HS65_LH_BFX4 U3566 ( .A(n2781), .Z(n2779) );
  HS65_LH_BFX4 U3567 ( .A(n2782), .Z(n2780) );
  HS65_LH_BFX4 U3568 ( .A(n2783), .Z(n2781) );
  HS65_LH_BFX4 U3569 ( .A(n2784), .Z(n2782) );
  HS65_LH_BFX4 U3570 ( .A(n2785), .Z(n2783) );
  HS65_LH_BFX4 U3571 ( .A(n2786), .Z(n2784) );
  HS65_LH_BFX4 U3572 ( .A(n2787), .Z(n2785) );
  HS65_LH_BFX4 U3573 ( .A(n2788), .Z(n2786) );
  HS65_LH_BFX4 U3574 ( .A(n2789), .Z(n2787) );
  HS65_LH_BFX4 U3575 ( .A(n2790), .Z(n2788) );
  HS65_LH_BFX4 U3576 ( .A(n2791), .Z(n2789) );
  HS65_LH_BFX4 U3577 ( .A(n2792), .Z(n2790) );
  HS65_LH_BFX4 U3578 ( .A(n2793), .Z(n2791) );
  HS65_LH_BFX4 U3579 ( .A(n2794), .Z(n2792) );
  HS65_LH_BFX4 U3580 ( .A(n2795), .Z(n2793) );
  HS65_LH_BFX4 U3581 ( .A(n2796), .Z(n2794) );
  HS65_LH_BFX4 U3582 ( .A(n2797), .Z(n2795) );
  HS65_LH_BFX4 U3583 ( .A(n2798), .Z(n2796) );
  HS65_LH_BFX4 U3584 ( .A(n2799), .Z(n2797) );
  HS65_LH_BFX4 U3585 ( .A(n2800), .Z(n2798) );
  HS65_LH_BFX4 U3586 ( .A(n2801), .Z(n2799) );
  HS65_LH_BFX4 U3587 ( .A(n2802), .Z(n2800) );
  HS65_LH_BFX4 U3588 ( .A(n2803), .Z(n2801) );
  HS65_LH_BFX4 U3589 ( .A(n2804), .Z(n2802) );
  HS65_LH_BFX4 U3590 ( .A(n2805), .Z(n2803) );
  HS65_LH_BFX4 U3591 ( .A(n2806), .Z(n2804) );
  HS65_LH_BFX4 U3592 ( .A(n2807), .Z(n2805) );
  HS65_LH_BFX4 U3593 ( .A(n2808), .Z(n2806) );
  HS65_LH_BFX4 U3594 ( .A(n2809), .Z(n2807) );
  HS65_LH_BFX4 U3595 ( .A(n2810), .Z(n2808) );
  HS65_LH_BFX4 U3596 ( .A(n2811), .Z(n2809) );
  HS65_LH_BFX4 U3597 ( .A(n2812), .Z(n2810) );
  HS65_LH_BFX4 U3598 ( .A(n2813), .Z(n2811) );
  HS65_LH_BFX4 U3599 ( .A(n2814), .Z(n2812) );
  HS65_LH_BFX4 U3600 ( .A(n2815), .Z(n2813) );
  HS65_LH_BFX4 U3601 ( .A(n2816), .Z(n2814) );
  HS65_LH_BFX4 U3602 ( .A(n2817), .Z(n2815) );
  HS65_LH_BFX4 U3603 ( .A(n2818), .Z(n2816) );
  HS65_LH_BFX4 U3604 ( .A(n2819), .Z(n2817) );
  HS65_LH_BFX4 U3605 ( .A(n2820), .Z(n2818) );
  HS65_LH_BFX4 U3606 ( .A(\u_DataPath/jump_address_i [0]), .Z(n2819) );
  HS65_LH_BFX4 U3607 ( .A(\u_DataPath/branch_target_i [0]), .Z(n2820) );
  HS65_LH_BFX4 U3608 ( .A(n2823), .Z(n2821) );
  HS65_LH_BFX4 U3609 ( .A(n2824), .Z(n2822) );
  HS65_LH_BFX4 U3610 ( .A(n2825), .Z(n2823) );
  HS65_LH_BFX4 U3611 ( .A(n2826), .Z(n2824) );
  HS65_LH_BFX4 U3612 ( .A(n2827), .Z(n2825) );
  HS65_LH_BFX4 U3613 ( .A(n2828), .Z(n2826) );
  HS65_LH_BFX4 U3614 ( .A(n2829), .Z(n2827) );
  HS65_LH_BFX4 U3615 ( .A(n2830), .Z(n2828) );
  HS65_LH_BFX4 U3616 ( .A(n2831), .Z(n2829) );
  HS65_LH_BFX4 U3617 ( .A(n2832), .Z(n2830) );
  HS65_LH_BFX4 U3618 ( .A(n2833), .Z(n2831) );
  HS65_LH_BFX4 U3619 ( .A(n2834), .Z(n2832) );
  HS65_LH_BFX4 U3620 ( .A(n2835), .Z(n2833) );
  HS65_LH_BFX4 U3621 ( .A(n2836), .Z(n2834) );
  HS65_LH_BFX4 U3622 ( .A(n2837), .Z(n2835) );
  HS65_LH_BFX4 U3623 ( .A(n2838), .Z(n2836) );
  HS65_LH_BFX4 U3624 ( .A(n2839), .Z(n2837) );
  HS65_LH_BFX4 U3625 ( .A(n2840), .Z(n2838) );
  HS65_LH_BFX4 U3626 ( .A(n2841), .Z(n2839) );
  HS65_LH_BFX4 U3627 ( .A(n2842), .Z(n2840) );
  HS65_LH_BFX4 U3628 ( .A(n2843), .Z(n2841) );
  HS65_LH_BFX4 U3629 ( .A(n2844), .Z(n2842) );
  HS65_LH_BFX4 U3630 ( .A(n2845), .Z(n2843) );
  HS65_LH_BFX4 U3631 ( .A(n2846), .Z(n2844) );
  HS65_LH_BFX4 U3632 ( .A(n2847), .Z(n2845) );
  HS65_LH_BFX4 U3633 ( .A(n2848), .Z(n2846) );
  HS65_LH_BFX4 U3634 ( .A(n2849), .Z(n2847) );
  HS65_LH_BFX4 U3635 ( .A(n2850), .Z(n2848) );
  HS65_LH_BFX4 U3636 ( .A(n2851), .Z(n2849) );
  HS65_LH_BFX4 U3637 ( .A(n2852), .Z(n2850) );
  HS65_LH_BFX4 U3638 ( .A(n2853), .Z(n2851) );
  HS65_LH_BFX4 U3639 ( .A(n2854), .Z(n2852) );
  HS65_LH_BFX4 U3640 ( .A(n2855), .Z(n2853) );
  HS65_LH_BFX4 U3641 ( .A(n2856), .Z(n2854) );
  HS65_LH_BFX4 U3642 ( .A(n2857), .Z(n2855) );
  HS65_LH_BFX4 U3643 ( .A(n2858), .Z(n2856) );
  HS65_LH_BFX4 U3644 ( .A(n2859), .Z(n2857) );
  HS65_LH_BFX4 U3645 ( .A(n2860), .Z(n2858) );
  HS65_LH_BFX4 U3646 ( .A(n2861), .Z(n2859) );
  HS65_LH_BFX4 U3647 ( .A(n2862), .Z(n2860) );
  HS65_LH_BFX4 U3648 ( .A(n2863), .Z(n2861) );
  HS65_LH_BFX4 U3649 ( .A(n2864), .Z(n2862) );
  HS65_LH_BFX4 U3650 ( .A(n2865), .Z(n2863) );
  HS65_LH_BFX4 U3651 ( .A(n2866), .Z(n2864) );
  HS65_LH_BFX4 U3652 ( .A(n2867), .Z(n2865) );
  HS65_LH_BFX4 U3653 ( .A(n2868), .Z(n2866) );
  HS65_LH_BFX4 U3654 ( .A(\u_DataPath/branch_target_i [1]), .Z(n2867) );
  HS65_LH_BFX4 U3655 ( .A(\u_DataPath/jump_address_i [1]), .Z(n2868) );
  HS65_LH_BFX4 U3656 ( .A(n2872), .Z(n2869) );
  HS65_LH_BFX4 U3657 ( .A(n2873), .Z(n2870) );
  HS65_LH_BFX4 U3658 ( .A(n12764), .Z(n2871) );
  HS65_LH_BFX4 U3659 ( .A(n2874), .Z(n2872) );
  HS65_LH_BFX4 U3660 ( .A(n2875), .Z(n2873) );
  HS65_LH_BFX4 U3661 ( .A(n2876), .Z(n2874) );
  HS65_LH_BFX4 U3662 ( .A(n2877), .Z(n2875) );
  HS65_LH_BFX4 U3663 ( .A(n2878), .Z(n2876) );
  HS65_LH_BFX4 U3664 ( .A(n2879), .Z(n2877) );
  HS65_LH_BFX4 U3665 ( .A(n2880), .Z(n2878) );
  HS65_LH_BFX4 U3666 ( .A(n2881), .Z(n2879) );
  HS65_LH_BFX4 U3667 ( .A(n2882), .Z(n2880) );
  HS65_LH_BFX4 U3668 ( .A(n2883), .Z(n2881) );
  HS65_LH_BFX4 U3669 ( .A(n2884), .Z(n2882) );
  HS65_LH_BFX4 U3670 ( .A(n2885), .Z(n2883) );
  HS65_LH_BFX4 U3671 ( .A(n2886), .Z(n2884) );
  HS65_LH_BFX4 U3672 ( .A(n2887), .Z(n2885) );
  HS65_LH_BFX4 U3673 ( .A(n2888), .Z(n2886) );
  HS65_LH_BFX4 U3674 ( .A(n2889), .Z(n2887) );
  HS65_LH_BFX4 U3675 ( .A(n2890), .Z(n2888) );
  HS65_LH_BFX4 U3676 ( .A(n2891), .Z(n2889) );
  HS65_LH_BFX4 U3677 ( .A(n2892), .Z(n2890) );
  HS65_LH_BFX4 U3678 ( .A(n2893), .Z(n2891) );
  HS65_LH_BFX4 U3679 ( .A(n2894), .Z(n2892) );
  HS65_LH_BFX4 U3680 ( .A(n2895), .Z(n2893) );
  HS65_LH_BFX4 U3681 ( .A(n2896), .Z(n2894) );
  HS65_LH_BFX4 U3682 ( .A(n2897), .Z(n2895) );
  HS65_LH_BFX4 U3683 ( .A(n2898), .Z(n2896) );
  HS65_LH_BFX4 U3684 ( .A(n2899), .Z(n2897) );
  HS65_LH_BFX4 U3685 ( .A(n2900), .Z(n2898) );
  HS65_LH_BFX4 U3686 ( .A(n2901), .Z(n2899) );
  HS65_LH_BFX4 U3687 ( .A(n2902), .Z(n2900) );
  HS65_LH_BFX4 U3688 ( .A(n2903), .Z(n2901) );
  HS65_LH_BFX4 U3689 ( .A(n2904), .Z(n2902) );
  HS65_LH_BFX4 U3690 ( .A(n2905), .Z(n2903) );
  HS65_LH_BFX4 U3691 ( .A(n2906), .Z(n2904) );
  HS65_LH_BFX4 U3692 ( .A(n2907), .Z(n2905) );
  HS65_LH_BFX4 U3693 ( .A(n2908), .Z(n2906) );
  HS65_LH_BFX4 U3694 ( .A(n2909), .Z(n2907) );
  HS65_LH_BFX4 U3695 ( .A(n2910), .Z(n2908) );
  HS65_LH_BFX4 U3696 ( .A(n2911), .Z(n2909) );
  HS65_LH_BFX4 U3697 ( .A(n2912), .Z(n2910) );
  HS65_LH_BFX4 U3698 ( .A(n2913), .Z(n2911) );
  HS65_LH_BFX4 U3699 ( .A(n2914), .Z(n2912) );
  HS65_LH_BFX4 U3700 ( .A(n2915), .Z(n2913) );
  HS65_LH_BFX4 U3701 ( .A(n2916), .Z(n2914) );
  HS65_LH_BFX4 U3702 ( .A(n2917), .Z(n2915) );
  HS65_LH_BFX4 U3703 ( .A(n2918), .Z(n2916) );
  HS65_LH_BFX4 U3704 ( .A(n2919), .Z(n2917) );
  HS65_LH_BFX4 U3705 ( .A(\u_DataPath/branch_target_i [6]), .Z(n2918) );
  HS65_LH_BFX4 U3706 ( .A(\u_DataPath/jump_address_i [6]), .Z(n2919) );
  HS65_LH_BFX4 U3707 ( .A(n2923), .Z(n2920) );
  HS65_LH_BFX4 U3708 ( .A(n2924), .Z(n2921) );
  HS65_LH_BFX4 U3709 ( .A(n2925), .Z(n2922) );
  HS65_LH_BFX4 U3710 ( .A(n12672), .Z(n2923) );
  HS65_LH_BFX4 U3711 ( .A(n2926), .Z(n2924) );
  HS65_LH_BFX4 U3712 ( .A(n2927), .Z(n2925) );
  HS65_LH_BFX4 U3713 ( .A(n2928), .Z(n2926) );
  HS65_LH_BFX4 U3714 ( .A(n2929), .Z(n2927) );
  HS65_LH_BFX4 U3715 ( .A(n2930), .Z(n2928) );
  HS65_LH_BFX4 U3716 ( .A(n2931), .Z(n2929) );
  HS65_LH_BFX4 U3717 ( .A(n2932), .Z(n2930) );
  HS65_LH_BFX4 U3718 ( .A(n2933), .Z(n2931) );
  HS65_LH_BFX4 U3719 ( .A(n2934), .Z(n2932) );
  HS65_LH_BFX4 U3720 ( .A(n2935), .Z(n2933) );
  HS65_LH_BFX4 U3721 ( .A(n2936), .Z(n2934) );
  HS65_LH_BFX4 U3722 ( .A(n2937), .Z(n2935) );
  HS65_LH_BFX4 U3723 ( .A(n2938), .Z(n2936) );
  HS65_LH_BFX4 U3724 ( .A(n2939), .Z(n2937) );
  HS65_LH_BFX4 U3725 ( .A(n2940), .Z(n2938) );
  HS65_LH_BFX4 U3726 ( .A(n2941), .Z(n2939) );
  HS65_LH_BFX4 U3727 ( .A(n2942), .Z(n2940) );
  HS65_LH_BFX4 U3728 ( .A(n2943), .Z(n2941) );
  HS65_LH_BFX4 U3729 ( .A(n2944), .Z(n2942) );
  HS65_LH_BFX4 U3730 ( .A(n2945), .Z(n2943) );
  HS65_LH_BFX4 U3731 ( .A(n2946), .Z(n2944) );
  HS65_LH_BFX4 U3732 ( .A(n2947), .Z(n2945) );
  HS65_LH_BFX4 U3733 ( .A(n2948), .Z(n2946) );
  HS65_LH_BFX4 U3734 ( .A(n2949), .Z(n2947) );
  HS65_LH_BFX4 U3735 ( .A(n2950), .Z(n2948) );
  HS65_LH_BFX4 U3736 ( .A(n2951), .Z(n2949) );
  HS65_LH_BFX4 U3737 ( .A(n2952), .Z(n2950) );
  HS65_LH_BFX4 U3738 ( .A(n2953), .Z(n2951) );
  HS65_LH_BFX4 U3739 ( .A(n2954), .Z(n2952) );
  HS65_LH_BFX4 U3740 ( .A(n2955), .Z(n2953) );
  HS65_LH_BFX4 U3741 ( .A(n2956), .Z(n2954) );
  HS65_LH_BFX4 U3742 ( .A(n2957), .Z(n2955) );
  HS65_LH_BFX4 U3743 ( .A(n2958), .Z(n2956) );
  HS65_LH_BFX4 U3744 ( .A(n2959), .Z(n2957) );
  HS65_LH_BFX4 U3745 ( .A(n2960), .Z(n2958) );
  HS65_LH_BFX4 U3746 ( .A(n2961), .Z(n2959) );
  HS65_LH_BFX4 U3747 ( .A(n2962), .Z(n2960) );
  HS65_LH_BFX4 U3748 ( .A(n2963), .Z(n2961) );
  HS65_LH_BFX4 U3749 ( .A(n2964), .Z(n2962) );
  HS65_LH_BFX4 U3750 ( .A(n2965), .Z(n2963) );
  HS65_LH_BFX4 U3751 ( .A(n2966), .Z(n2964) );
  HS65_LH_BFX4 U3752 ( .A(n2967), .Z(n2965) );
  HS65_LH_BFX4 U3753 ( .A(n2968), .Z(n2966) );
  HS65_LH_BFX4 U3754 ( .A(n2969), .Z(n2967) );
  HS65_LH_BFX4 U3755 ( .A(n2970), .Z(n2968) );
  HS65_LH_BFX4 U3756 ( .A(n2971), .Z(n2969) );
  HS65_LH_BFX4 U3757 ( .A(\u_DataPath/branch_target_i [4]), .Z(n2970) );
  HS65_LH_BFX4 U3758 ( .A(\u_DataPath/jump_address_i [4]), .Z(n2971) );
  HS65_LH_BFX4 U3759 ( .A(n9480), .Z(n2972) );
  HS65_LH_BFX4 U3760 ( .A(n13890), .Z(n2973) );
  HS65_LH_IVX13 U3761 ( .A(n12806), .Z(n13947) );
  HS65_LH_BFX4 U3762 ( .A(n14082), .Z(n2974) );
  HS65_LH_BFX4 U3763 ( .A(n2977), .Z(n2975) );
  HS65_LH_BFX4 U3764 ( .A(n2978), .Z(n2976) );
  HS65_LH_BFX4 U3765 ( .A(n2979), .Z(n2977) );
  HS65_LH_BFX4 U3766 ( .A(n2980), .Z(n2978) );
  HS65_LH_BFX4 U3767 ( .A(n2981), .Z(n2979) );
  HS65_LH_BFX4 U3768 ( .A(n2982), .Z(n2980) );
  HS65_LH_BFX4 U3769 ( .A(n2983), .Z(n2981) );
  HS65_LH_BFX4 U3770 ( .A(n2984), .Z(n2982) );
  HS65_LH_BFX4 U3771 ( .A(n2985), .Z(n2983) );
  HS65_LH_BFX4 U3772 ( .A(n2986), .Z(n2984) );
  HS65_LH_BFX4 U3773 ( .A(n2987), .Z(n2985) );
  HS65_LH_BFX4 U3774 ( .A(n2988), .Z(n2986) );
  HS65_LH_BFX4 U3775 ( .A(n2989), .Z(n2987) );
  HS65_LH_BFX4 U3776 ( .A(n2990), .Z(n2988) );
  HS65_LH_BFX4 U3777 ( .A(n2991), .Z(n2989) );
  HS65_LH_BFX4 U3778 ( .A(n2992), .Z(n2990) );
  HS65_LH_BFX4 U3779 ( .A(n2993), .Z(n2991) );
  HS65_LH_BFX4 U3780 ( .A(n2994), .Z(n2992) );
  HS65_LH_BFX4 U3781 ( .A(n2995), .Z(n2993) );
  HS65_LH_BFX4 U3782 ( .A(n2996), .Z(n2994) );
  HS65_LH_BFX4 U3783 ( .A(n2997), .Z(n2995) );
  HS65_LH_BFX4 U3784 ( .A(n2998), .Z(n2996) );
  HS65_LH_BFX4 U3785 ( .A(n2999), .Z(n2997) );
  HS65_LH_BFX4 U3786 ( .A(n3000), .Z(n2998) );
  HS65_LH_BFX4 U3787 ( .A(n3001), .Z(n2999) );
  HS65_LH_BFX4 U3788 ( .A(n3002), .Z(n3000) );
  HS65_LH_BFX4 U3789 ( .A(n3003), .Z(n3001) );
  HS65_LH_BFX4 U3790 ( .A(n3004), .Z(n3002) );
  HS65_LH_BFX4 U3791 ( .A(n3005), .Z(n3003) );
  HS65_LH_BFX4 U3792 ( .A(n3006), .Z(n3004) );
  HS65_LH_BFX4 U3793 ( .A(n3007), .Z(n3005) );
  HS65_LH_BFX4 U3794 ( .A(n3008), .Z(n3006) );
  HS65_LH_BFX4 U3795 ( .A(n3009), .Z(n3007) );
  HS65_LH_BFX4 U3796 ( .A(n3010), .Z(n3008) );
  HS65_LH_BFX4 U3797 ( .A(n3011), .Z(n3009) );
  HS65_LH_BFX4 U3798 ( .A(n3012), .Z(n3010) );
  HS65_LH_BFX4 U3799 ( .A(n3013), .Z(n3011) );
  HS65_LH_BFX4 U3800 ( .A(n3014), .Z(n3012) );
  HS65_LH_BFX4 U3801 ( .A(n3015), .Z(n3013) );
  HS65_LH_BFX4 U3802 ( .A(n3016), .Z(n3014) );
  HS65_LH_BFX4 U3803 ( .A(n3017), .Z(n3015) );
  HS65_LH_BFX4 U3804 ( .A(n3018), .Z(n3016) );
  HS65_LH_BFX4 U3805 ( .A(n3019), .Z(n3017) );
  HS65_LH_BFX4 U3806 ( .A(n3020), .Z(n3018) );
  HS65_LH_BFX4 U3807 ( .A(n3021), .Z(n3019) );
  HS65_LH_BFX4 U3808 ( .A(n3022), .Z(n3020) );
  HS65_LH_BFX4 U3809 ( .A(n3023), .Z(n3021) );
  HS65_LH_BFX4 U3810 ( .A(n3024), .Z(n3022) );
  HS65_LH_BFX4 U3811 ( .A(\u_DataPath/branch_target_i [7]), .Z(n3023) );
  HS65_LH_BFX4 U3812 ( .A(\u_DataPath/jump_address_i [7]), .Z(n3024) );
  HS65_LH_BFX4 U3813 ( .A(n3028), .Z(n3025) );
  HS65_LH_BFX4 U3814 ( .A(n3029), .Z(n3026) );
  HS65_LH_BFX4 U3815 ( .A(n3030), .Z(n3027) );
  HS65_LH_BFX4 U3816 ( .A(n3031), .Z(n3028) );
  HS65_LH_BFX4 U3817 ( .A(n12851), .Z(n3029) );
  HS65_LH_BFX4 U3818 ( .A(n3032), .Z(n3030) );
  HS65_LH_BFX4 U3819 ( .A(n3033), .Z(n3031) );
  HS65_LH_BFX4 U3820 ( .A(n3034), .Z(n3032) );
  HS65_LH_BFX4 U3821 ( .A(n3035), .Z(n3033) );
  HS65_LH_BFX4 U3822 ( .A(n3036), .Z(n3034) );
  HS65_LH_BFX4 U3823 ( .A(n3037), .Z(n3035) );
  HS65_LH_BFX4 U3824 ( .A(n3038), .Z(n3036) );
  HS65_LH_BFX4 U3825 ( .A(n3039), .Z(n3037) );
  HS65_LH_BFX4 U3826 ( .A(n3040), .Z(n3038) );
  HS65_LH_BFX4 U3827 ( .A(n3041), .Z(n3039) );
  HS65_LH_BFX4 U3828 ( .A(n3042), .Z(n3040) );
  HS65_LH_BFX4 U3829 ( .A(n3043), .Z(n3041) );
  HS65_LH_BFX4 U3830 ( .A(n3044), .Z(n3042) );
  HS65_LH_BFX4 U3831 ( .A(n3045), .Z(n3043) );
  HS65_LH_BFX4 U3832 ( .A(n3046), .Z(n3044) );
  HS65_LH_BFX4 U3833 ( .A(n3047), .Z(n3045) );
  HS65_LH_BFX4 U3834 ( .A(n3048), .Z(n3046) );
  HS65_LH_BFX4 U3835 ( .A(n3049), .Z(n3047) );
  HS65_LH_BFX4 U3836 ( .A(n3050), .Z(n3048) );
  HS65_LH_BFX4 U3837 ( .A(n3051), .Z(n3049) );
  HS65_LH_BFX4 U3838 ( .A(n3052), .Z(n3050) );
  HS65_LH_BFX4 U3839 ( .A(n3053), .Z(n3051) );
  HS65_LH_BFX4 U3840 ( .A(n3054), .Z(n3052) );
  HS65_LH_BFX4 U3841 ( .A(n3055), .Z(n3053) );
  HS65_LH_BFX4 U3842 ( .A(n3056), .Z(n3054) );
  HS65_LH_BFX4 U3843 ( .A(n3057), .Z(n3055) );
  HS65_LH_BFX4 U3844 ( .A(n3058), .Z(n3056) );
  HS65_LH_BFX4 U3845 ( .A(n3059), .Z(n3057) );
  HS65_LH_BFX4 U3846 ( .A(n3060), .Z(n3058) );
  HS65_LH_BFX4 U3847 ( .A(n3061), .Z(n3059) );
  HS65_LH_BFX4 U3848 ( .A(n3062), .Z(n3060) );
  HS65_LH_BFX4 U3849 ( .A(n3063), .Z(n3061) );
  HS65_LH_BFX4 U3850 ( .A(n3064), .Z(n3062) );
  HS65_LH_BFX4 U3851 ( .A(n3065), .Z(n3063) );
  HS65_LH_BFX4 U3852 ( .A(n3066), .Z(n3064) );
  HS65_LH_BFX4 U3853 ( .A(n3067), .Z(n3065) );
  HS65_LH_BFX4 U3854 ( .A(n3068), .Z(n3066) );
  HS65_LH_BFX4 U3855 ( .A(n3069), .Z(n3067) );
  HS65_LH_BFX4 U3856 ( .A(n3070), .Z(n3068) );
  HS65_LH_BFX4 U3857 ( .A(n3071), .Z(n3069) );
  HS65_LH_BFX4 U3858 ( .A(n3072), .Z(n3070) );
  HS65_LH_BFX4 U3859 ( .A(n3073), .Z(n3071) );
  HS65_LH_BFX4 U3860 ( .A(n3074), .Z(n3072) );
  HS65_LH_BFX4 U3861 ( .A(n3075), .Z(n3073) );
  HS65_LH_BFX4 U3862 ( .A(n3076), .Z(n3074) );
  HS65_LH_BFX4 U3863 ( .A(\u_DataPath/branch_target_i [8]), .Z(n3075) );
  HS65_LH_BFX4 U3864 ( .A(\u_DataPath/jump_address_i [8]), .Z(n3076) );
  HS65_LH_IVX13 U3865 ( .A(n12896), .Z(n13949) );
  HS65_LH_BFX4 U3866 ( .A(n14084), .Z(n3077) );
  HS65_LH_BFX4 U3867 ( .A(n3080), .Z(n3078) );
  HS65_LH_BFX4 U3868 ( .A(n3081), .Z(n3079) );
  HS65_LH_BFX4 U3869 ( .A(n3082), .Z(n3080) );
  HS65_LH_BFX4 U3870 ( .A(n3083), .Z(n3081) );
  HS65_LH_BFX4 U3871 ( .A(n3084), .Z(n3082) );
  HS65_LH_BFX4 U3872 ( .A(n3085), .Z(n3083) );
  HS65_LH_BFX4 U3873 ( .A(n3086), .Z(n3084) );
  HS65_LH_BFX4 U3874 ( .A(n3087), .Z(n3085) );
  HS65_LH_BFX4 U3875 ( .A(n3088), .Z(n3086) );
  HS65_LH_BFX4 U3876 ( .A(n3089), .Z(n3087) );
  HS65_LH_BFX4 U3877 ( .A(n3090), .Z(n3088) );
  HS65_LH_BFX4 U3878 ( .A(n3091), .Z(n3089) );
  HS65_LH_BFX4 U3879 ( .A(n3092), .Z(n3090) );
  HS65_LH_BFX4 U3880 ( .A(n3093), .Z(n3091) );
  HS65_LH_BFX4 U3881 ( .A(n3094), .Z(n3092) );
  HS65_LH_BFX4 U3882 ( .A(n3095), .Z(n3093) );
  HS65_LH_BFX4 U3883 ( .A(n3096), .Z(n3094) );
  HS65_LH_BFX4 U3884 ( .A(n3097), .Z(n3095) );
  HS65_LH_BFX4 U3885 ( .A(n3098), .Z(n3096) );
  HS65_LH_BFX4 U3886 ( .A(n3099), .Z(n3097) );
  HS65_LH_BFX4 U3887 ( .A(n3100), .Z(n3098) );
  HS65_LH_BFX4 U3888 ( .A(n3101), .Z(n3099) );
  HS65_LH_BFX4 U3889 ( .A(n3102), .Z(n3100) );
  HS65_LH_BFX4 U3890 ( .A(n3103), .Z(n3101) );
  HS65_LH_BFX4 U3891 ( .A(n3104), .Z(n3102) );
  HS65_LH_BFX4 U3892 ( .A(n3105), .Z(n3103) );
  HS65_LH_BFX4 U3893 ( .A(n3106), .Z(n3104) );
  HS65_LH_BFX4 U3894 ( .A(n3107), .Z(n3105) );
  HS65_LH_BFX4 U3895 ( .A(n3108), .Z(n3106) );
  HS65_LH_BFX4 U3896 ( .A(n3109), .Z(n3107) );
  HS65_LH_BFX4 U3897 ( .A(n3110), .Z(n3108) );
  HS65_LH_BFX4 U3898 ( .A(n3111), .Z(n3109) );
  HS65_LH_BFX4 U3899 ( .A(n3112), .Z(n3110) );
  HS65_LH_BFX4 U3900 ( .A(n3113), .Z(n3111) );
  HS65_LH_BFX4 U3901 ( .A(n3114), .Z(n3112) );
  HS65_LH_BFX4 U3902 ( .A(n3115), .Z(n3113) );
  HS65_LH_BFX4 U3903 ( .A(n3116), .Z(n3114) );
  HS65_LH_BFX4 U3904 ( .A(n3117), .Z(n3115) );
  HS65_LH_BFX4 U3905 ( .A(n3118), .Z(n3116) );
  HS65_LH_BFX4 U3906 ( .A(n3119), .Z(n3117) );
  HS65_LH_BFX4 U3907 ( .A(n3120), .Z(n3118) );
  HS65_LH_BFX4 U3908 ( .A(n3121), .Z(n3119) );
  HS65_LH_BFX4 U3909 ( .A(n3122), .Z(n3120) );
  HS65_LH_BFX4 U3910 ( .A(n3123), .Z(n3121) );
  HS65_LH_BFX4 U3911 ( .A(n3124), .Z(n3122) );
  HS65_LH_BFX4 U3912 ( .A(n3125), .Z(n3123) );
  HS65_LH_BFX4 U3913 ( .A(n3126), .Z(n3124) );
  HS65_LH_BFX4 U3914 ( .A(n3127), .Z(n3125) );
  HS65_LH_BFX4 U3915 ( .A(\u_DataPath/branch_target_i [9]), .Z(n3126) );
  HS65_LH_BFX4 U3916 ( .A(\u_DataPath/jump_address_i [9]), .Z(n3127) );
  HS65_LH_BFX4 U3917 ( .A(n3131), .Z(n3128) );
  HS65_LH_BFX4 U3918 ( .A(n3132), .Z(n3129) );
  HS65_LH_BFX4 U3919 ( .A(n3133), .Z(n3130) );
  HS65_LH_BFX4 U3920 ( .A(n3134), .Z(n3131) );
  HS65_LH_BFX4 U3921 ( .A(n12941), .Z(n3132) );
  HS65_LH_BFX4 U3922 ( .A(n3135), .Z(n3133) );
  HS65_LH_BFX4 U3923 ( .A(n3136), .Z(n3134) );
  HS65_LH_BFX4 U3924 ( .A(n3137), .Z(n3135) );
  HS65_LH_BFX4 U3925 ( .A(n3138), .Z(n3136) );
  HS65_LH_BFX4 U3926 ( .A(n3139), .Z(n3137) );
  HS65_LH_BFX4 U3927 ( .A(n3140), .Z(n3138) );
  HS65_LH_BFX4 U3928 ( .A(n3141), .Z(n3139) );
  HS65_LH_BFX4 U3929 ( .A(n3142), .Z(n3140) );
  HS65_LH_BFX4 U3930 ( .A(n3143), .Z(n3141) );
  HS65_LH_BFX4 U3931 ( .A(n3144), .Z(n3142) );
  HS65_LH_BFX4 U3932 ( .A(n3145), .Z(n3143) );
  HS65_LH_BFX4 U3933 ( .A(n3146), .Z(n3144) );
  HS65_LH_BFX4 U3934 ( .A(n3147), .Z(n3145) );
  HS65_LH_BFX4 U3935 ( .A(n3148), .Z(n3146) );
  HS65_LH_BFX4 U3936 ( .A(n3149), .Z(n3147) );
  HS65_LH_BFX4 U3937 ( .A(n3150), .Z(n3148) );
  HS65_LH_BFX4 U3938 ( .A(n3151), .Z(n3149) );
  HS65_LH_BFX4 U3939 ( .A(n3152), .Z(n3150) );
  HS65_LH_BFX4 U3940 ( .A(n3153), .Z(n3151) );
  HS65_LH_BFX4 U3941 ( .A(n3154), .Z(n3152) );
  HS65_LH_BFX4 U3942 ( .A(n3155), .Z(n3153) );
  HS65_LH_BFX4 U3943 ( .A(n3156), .Z(n3154) );
  HS65_LH_BFX4 U3944 ( .A(n3157), .Z(n3155) );
  HS65_LH_BFX4 U3945 ( .A(n3158), .Z(n3156) );
  HS65_LH_BFX4 U3946 ( .A(n3159), .Z(n3157) );
  HS65_LH_BFX4 U3947 ( .A(n3160), .Z(n3158) );
  HS65_LH_BFX4 U3948 ( .A(n3161), .Z(n3159) );
  HS65_LH_BFX4 U3949 ( .A(n3162), .Z(n3160) );
  HS65_LH_BFX4 U3950 ( .A(n3163), .Z(n3161) );
  HS65_LH_BFX4 U3951 ( .A(n3164), .Z(n3162) );
  HS65_LH_BFX4 U3952 ( .A(n3165), .Z(n3163) );
  HS65_LH_BFX4 U3953 ( .A(n3166), .Z(n3164) );
  HS65_LH_BFX4 U3954 ( .A(n3167), .Z(n3165) );
  HS65_LH_BFX4 U3955 ( .A(n3168), .Z(n3166) );
  HS65_LH_BFX4 U3956 ( .A(n3169), .Z(n3167) );
  HS65_LH_BFX4 U3957 ( .A(n3170), .Z(n3168) );
  HS65_LH_BFX4 U3958 ( .A(n3171), .Z(n3169) );
  HS65_LH_BFX4 U3959 ( .A(n3172), .Z(n3170) );
  HS65_LH_BFX4 U3960 ( .A(n3173), .Z(n3171) );
  HS65_LH_BFX4 U3961 ( .A(n3174), .Z(n3172) );
  HS65_LH_BFX4 U3962 ( .A(n3175), .Z(n3173) );
  HS65_LH_BFX4 U3963 ( .A(n3176), .Z(n3174) );
  HS65_LH_BFX4 U3964 ( .A(n3177), .Z(n3175) );
  HS65_LH_BFX4 U3965 ( .A(n3178), .Z(n3176) );
  HS65_LH_BFX4 U3966 ( .A(n3179), .Z(n3177) );
  HS65_LH_BFX4 U3967 ( .A(\u_DataPath/branch_target_i [10]), .Z(n3178) );
  HS65_LH_BFX4 U3968 ( .A(\u_DataPath/jump_address_i [10]), .Z(n3179) );
  HS65_LH_IVX13 U3969 ( .A(n12986), .Z(n13951) );
  HS65_LH_BFX4 U3970 ( .A(n14086), .Z(n3180) );
  HS65_LH_BFX4 U3971 ( .A(n3183), .Z(n3181) );
  HS65_LH_BFX4 U3972 ( .A(n3184), .Z(n3182) );
  HS65_LH_BFX4 U3973 ( .A(n3185), .Z(n3183) );
  HS65_LH_BFX4 U3974 ( .A(n3186), .Z(n3184) );
  HS65_LH_BFX4 U3975 ( .A(n3187), .Z(n3185) );
  HS65_LH_BFX4 U3976 ( .A(n3188), .Z(n3186) );
  HS65_LH_BFX4 U3977 ( .A(n3189), .Z(n3187) );
  HS65_LH_BFX4 U3978 ( .A(n3190), .Z(n3188) );
  HS65_LH_BFX4 U3979 ( .A(n3191), .Z(n3189) );
  HS65_LH_BFX4 U3980 ( .A(n3192), .Z(n3190) );
  HS65_LH_BFX4 U3981 ( .A(n3193), .Z(n3191) );
  HS65_LH_BFX4 U3982 ( .A(n3194), .Z(n3192) );
  HS65_LH_BFX4 U3983 ( .A(n3195), .Z(n3193) );
  HS65_LH_BFX4 U3984 ( .A(n3196), .Z(n3194) );
  HS65_LH_BFX4 U3985 ( .A(n3197), .Z(n3195) );
  HS65_LH_BFX4 U3986 ( .A(n3198), .Z(n3196) );
  HS65_LH_BFX4 U3987 ( .A(n3199), .Z(n3197) );
  HS65_LH_BFX4 U3988 ( .A(n3200), .Z(n3198) );
  HS65_LH_BFX4 U3989 ( .A(n3201), .Z(n3199) );
  HS65_LH_BFX4 U3990 ( .A(n3202), .Z(n3200) );
  HS65_LH_BFX4 U3991 ( .A(n3203), .Z(n3201) );
  HS65_LH_BFX4 U3992 ( .A(n3204), .Z(n3202) );
  HS65_LH_BFX4 U3993 ( .A(n3205), .Z(n3203) );
  HS65_LH_BFX4 U3994 ( .A(n3206), .Z(n3204) );
  HS65_LH_BFX4 U3995 ( .A(n3207), .Z(n3205) );
  HS65_LH_BFX4 U3996 ( .A(n3208), .Z(n3206) );
  HS65_LH_BFX4 U3997 ( .A(n3209), .Z(n3207) );
  HS65_LH_BFX4 U3998 ( .A(n3210), .Z(n3208) );
  HS65_LH_BFX4 U3999 ( .A(n3211), .Z(n3209) );
  HS65_LH_BFX4 U4000 ( .A(n3212), .Z(n3210) );
  HS65_LH_BFX4 U4001 ( .A(n3213), .Z(n3211) );
  HS65_LH_BFX4 U4002 ( .A(n3214), .Z(n3212) );
  HS65_LH_BFX4 U4003 ( .A(n3215), .Z(n3213) );
  HS65_LH_BFX4 U4004 ( .A(n3216), .Z(n3214) );
  HS65_LH_BFX4 U4005 ( .A(n3217), .Z(n3215) );
  HS65_LH_BFX4 U4006 ( .A(n3218), .Z(n3216) );
  HS65_LH_BFX4 U4007 ( .A(n3219), .Z(n3217) );
  HS65_LH_BFX4 U4008 ( .A(n3220), .Z(n3218) );
  HS65_LH_BFX4 U4009 ( .A(n3221), .Z(n3219) );
  HS65_LH_BFX4 U4010 ( .A(n3222), .Z(n3220) );
  HS65_LH_BFX4 U4011 ( .A(n3223), .Z(n3221) );
  HS65_LH_BFX4 U4012 ( .A(n3224), .Z(n3222) );
  HS65_LH_BFX4 U4013 ( .A(n3225), .Z(n3223) );
  HS65_LH_BFX4 U4014 ( .A(n3226), .Z(n3224) );
  HS65_LH_BFX4 U4015 ( .A(n3227), .Z(n3225) );
  HS65_LH_BFX4 U4016 ( .A(n3228), .Z(n3226) );
  HS65_LH_BFX4 U4017 ( .A(n3229), .Z(n3227) );
  HS65_LH_BFX4 U4018 ( .A(n3230), .Z(n3228) );
  HS65_LH_BFX4 U4019 ( .A(\u_DataPath/branch_target_i [11]), .Z(n3229) );
  HS65_LH_BFX4 U4020 ( .A(\u_DataPath/jump_address_i [11]), .Z(n3230) );
  HS65_LH_BFX4 U4021 ( .A(n3234), .Z(n3231) );
  HS65_LH_BFX4 U4022 ( .A(n3235), .Z(n3232) );
  HS65_LH_BFX4 U4023 ( .A(n3236), .Z(n3233) );
  HS65_LH_BFX4 U4024 ( .A(n3237), .Z(n3234) );
  HS65_LH_BFX4 U4025 ( .A(n13031), .Z(n3235) );
  HS65_LH_BFX4 U4026 ( .A(n3238), .Z(n3236) );
  HS65_LH_BFX4 U4027 ( .A(n3239), .Z(n3237) );
  HS65_LH_BFX4 U4028 ( .A(n3240), .Z(n3238) );
  HS65_LH_BFX4 U4029 ( .A(n3241), .Z(n3239) );
  HS65_LH_BFX4 U4030 ( .A(n3242), .Z(n3240) );
  HS65_LH_BFX4 U4031 ( .A(n3243), .Z(n3241) );
  HS65_LH_BFX4 U4032 ( .A(n3244), .Z(n3242) );
  HS65_LH_BFX4 U4033 ( .A(n3245), .Z(n3243) );
  HS65_LH_BFX4 U4034 ( .A(n3246), .Z(n3244) );
  HS65_LH_BFX4 U4035 ( .A(n3247), .Z(n3245) );
  HS65_LH_BFX4 U4036 ( .A(n3248), .Z(n3246) );
  HS65_LH_BFX4 U4037 ( .A(n3249), .Z(n3247) );
  HS65_LH_BFX4 U4038 ( .A(n3250), .Z(n3248) );
  HS65_LH_BFX4 U4039 ( .A(n3251), .Z(n3249) );
  HS65_LH_BFX4 U4040 ( .A(n3252), .Z(n3250) );
  HS65_LH_BFX4 U4041 ( .A(n3253), .Z(n3251) );
  HS65_LH_BFX4 U4042 ( .A(n3254), .Z(n3252) );
  HS65_LH_BFX4 U4043 ( .A(n3255), .Z(n3253) );
  HS65_LH_BFX4 U4044 ( .A(n3256), .Z(n3254) );
  HS65_LH_BFX4 U4045 ( .A(n3257), .Z(n3255) );
  HS65_LH_BFX4 U4046 ( .A(n3258), .Z(n3256) );
  HS65_LH_BFX4 U4047 ( .A(n3259), .Z(n3257) );
  HS65_LH_BFX4 U4048 ( .A(n3260), .Z(n3258) );
  HS65_LH_BFX4 U4049 ( .A(n3261), .Z(n3259) );
  HS65_LH_BFX4 U4050 ( .A(n3262), .Z(n3260) );
  HS65_LH_BFX4 U4051 ( .A(n3263), .Z(n3261) );
  HS65_LH_BFX4 U4052 ( .A(n3264), .Z(n3262) );
  HS65_LH_BFX4 U4053 ( .A(n3265), .Z(n3263) );
  HS65_LH_BFX4 U4054 ( .A(n3266), .Z(n3264) );
  HS65_LH_BFX4 U4055 ( .A(n3267), .Z(n3265) );
  HS65_LH_BFX4 U4056 ( .A(n3268), .Z(n3266) );
  HS65_LH_BFX4 U4057 ( .A(n3269), .Z(n3267) );
  HS65_LH_BFX4 U4058 ( .A(n3270), .Z(n3268) );
  HS65_LH_BFX4 U4059 ( .A(n3271), .Z(n3269) );
  HS65_LH_BFX4 U4060 ( .A(n3272), .Z(n3270) );
  HS65_LH_BFX4 U4061 ( .A(n3273), .Z(n3271) );
  HS65_LH_BFX4 U4062 ( .A(n3274), .Z(n3272) );
  HS65_LH_BFX4 U4063 ( .A(n3275), .Z(n3273) );
  HS65_LH_BFX4 U4064 ( .A(n3276), .Z(n3274) );
  HS65_LH_BFX4 U4065 ( .A(n3277), .Z(n3275) );
  HS65_LH_BFX4 U4066 ( .A(n3278), .Z(n3276) );
  HS65_LH_BFX4 U4067 ( .A(n3279), .Z(n3277) );
  HS65_LH_BFX4 U4068 ( .A(n3280), .Z(n3278) );
  HS65_LH_BFX4 U4069 ( .A(n3281), .Z(n3279) );
  HS65_LH_BFX4 U4070 ( .A(n3282), .Z(n3280) );
  HS65_LH_BFX4 U4071 ( .A(\u_DataPath/branch_target_i [12]), .Z(n3281) );
  HS65_LH_BFX4 U4072 ( .A(\u_DataPath/jump_address_i [12]), .Z(n3282) );
  HS65_LH_IVX13 U4073 ( .A(n13076), .Z(n13953) );
  HS65_LH_BFX4 U4074 ( .A(n14088), .Z(n3283) );
  HS65_LH_BFX4 U4075 ( .A(n3286), .Z(n3284) );
  HS65_LH_BFX4 U4076 ( .A(n3287), .Z(n3285) );
  HS65_LH_BFX4 U4077 ( .A(n3288), .Z(n3286) );
  HS65_LH_BFX4 U4078 ( .A(n3289), .Z(n3287) );
  HS65_LH_BFX4 U4079 ( .A(n3290), .Z(n3288) );
  HS65_LH_BFX4 U4080 ( .A(n3291), .Z(n3289) );
  HS65_LH_BFX4 U4081 ( .A(n3292), .Z(n3290) );
  HS65_LH_BFX4 U4082 ( .A(n3293), .Z(n3291) );
  HS65_LH_BFX4 U4083 ( .A(n3294), .Z(n3292) );
  HS65_LH_BFX4 U4084 ( .A(n3295), .Z(n3293) );
  HS65_LH_BFX4 U4085 ( .A(n3296), .Z(n3294) );
  HS65_LH_BFX4 U4086 ( .A(n3297), .Z(n3295) );
  HS65_LH_BFX4 U4087 ( .A(n3298), .Z(n3296) );
  HS65_LH_BFX4 U4088 ( .A(n3299), .Z(n3297) );
  HS65_LH_BFX4 U4089 ( .A(n3300), .Z(n3298) );
  HS65_LH_BFX4 U4090 ( .A(n3301), .Z(n3299) );
  HS65_LH_BFX4 U4091 ( .A(n3302), .Z(n3300) );
  HS65_LH_BFX4 U4092 ( .A(n3303), .Z(n3301) );
  HS65_LH_BFX4 U4093 ( .A(n3304), .Z(n3302) );
  HS65_LH_BFX4 U4094 ( .A(n3305), .Z(n3303) );
  HS65_LH_BFX4 U4095 ( .A(n3306), .Z(n3304) );
  HS65_LH_BFX4 U4096 ( .A(n3307), .Z(n3305) );
  HS65_LH_BFX4 U4097 ( .A(n3308), .Z(n3306) );
  HS65_LH_BFX4 U4098 ( .A(n3309), .Z(n3307) );
  HS65_LH_BFX4 U4099 ( .A(n3310), .Z(n3308) );
  HS65_LH_BFX4 U4100 ( .A(n3311), .Z(n3309) );
  HS65_LH_BFX4 U4101 ( .A(n3312), .Z(n3310) );
  HS65_LH_BFX4 U4102 ( .A(n3313), .Z(n3311) );
  HS65_LH_BFX4 U4103 ( .A(n3314), .Z(n3312) );
  HS65_LH_BFX4 U4104 ( .A(n3315), .Z(n3313) );
  HS65_LH_BFX4 U4105 ( .A(n3316), .Z(n3314) );
  HS65_LH_BFX4 U4106 ( .A(n3317), .Z(n3315) );
  HS65_LH_BFX4 U4107 ( .A(n3318), .Z(n3316) );
  HS65_LH_BFX4 U4108 ( .A(n3319), .Z(n3317) );
  HS65_LH_BFX4 U4109 ( .A(n3320), .Z(n3318) );
  HS65_LH_BFX4 U4110 ( .A(n3321), .Z(n3319) );
  HS65_LH_BFX4 U4111 ( .A(n3322), .Z(n3320) );
  HS65_LH_BFX4 U4112 ( .A(n3323), .Z(n3321) );
  HS65_LH_BFX4 U4113 ( .A(n3324), .Z(n3322) );
  HS65_LH_BFX4 U4114 ( .A(n3325), .Z(n3323) );
  HS65_LH_BFX4 U4115 ( .A(n3326), .Z(n3324) );
  HS65_LH_BFX4 U4116 ( .A(n3327), .Z(n3325) );
  HS65_LH_BFX4 U4117 ( .A(n3328), .Z(n3326) );
  HS65_LH_BFX4 U4118 ( .A(n3329), .Z(n3327) );
  HS65_LH_BFX4 U4119 ( .A(n3330), .Z(n3328) );
  HS65_LH_BFX4 U4120 ( .A(n3331), .Z(n3329) );
  HS65_LH_BFX4 U4121 ( .A(n3332), .Z(n3330) );
  HS65_LH_BFX4 U4122 ( .A(n3333), .Z(n3331) );
  HS65_LH_BFX4 U4123 ( .A(\u_DataPath/branch_target_i [13]), .Z(n3332) );
  HS65_LH_BFX4 U4124 ( .A(\u_DataPath/jump_address_i [13]), .Z(n3333) );
  HS65_LH_BFX4 U4125 ( .A(n3337), .Z(n3334) );
  HS65_LH_BFX4 U4126 ( .A(n3338), .Z(n3335) );
  HS65_LH_BFX4 U4127 ( .A(n3339), .Z(n3336) );
  HS65_LH_BFX4 U4128 ( .A(n3340), .Z(n3337) );
  HS65_LH_BFX4 U4129 ( .A(n13121), .Z(n3338) );
  HS65_LH_BFX4 U4130 ( .A(n3341), .Z(n3339) );
  HS65_LH_BFX4 U4131 ( .A(n3342), .Z(n3340) );
  HS65_LH_BFX4 U4132 ( .A(n3343), .Z(n3341) );
  HS65_LH_BFX4 U4133 ( .A(n3344), .Z(n3342) );
  HS65_LH_BFX4 U4134 ( .A(n3345), .Z(n3343) );
  HS65_LH_BFX4 U4135 ( .A(n3346), .Z(n3344) );
  HS65_LH_BFX4 U4136 ( .A(n3347), .Z(n3345) );
  HS65_LH_BFX4 U4137 ( .A(n3348), .Z(n3346) );
  HS65_LH_BFX4 U4138 ( .A(n3349), .Z(n3347) );
  HS65_LH_BFX4 U4139 ( .A(n3350), .Z(n3348) );
  HS65_LH_BFX4 U4140 ( .A(n3351), .Z(n3349) );
  HS65_LH_BFX4 U4141 ( .A(n3352), .Z(n3350) );
  HS65_LH_BFX4 U4142 ( .A(n3353), .Z(n3351) );
  HS65_LH_BFX4 U4143 ( .A(n3354), .Z(n3352) );
  HS65_LH_BFX4 U4144 ( .A(n3355), .Z(n3353) );
  HS65_LH_BFX4 U4145 ( .A(n3356), .Z(n3354) );
  HS65_LH_BFX4 U4146 ( .A(n3357), .Z(n3355) );
  HS65_LH_BFX4 U4147 ( .A(n3358), .Z(n3356) );
  HS65_LH_BFX4 U4148 ( .A(n3359), .Z(n3357) );
  HS65_LH_BFX4 U4149 ( .A(n3360), .Z(n3358) );
  HS65_LH_BFX4 U4150 ( .A(n3361), .Z(n3359) );
  HS65_LH_BFX4 U4151 ( .A(n3362), .Z(n3360) );
  HS65_LH_BFX4 U4152 ( .A(n3363), .Z(n3361) );
  HS65_LH_BFX4 U4153 ( .A(n3364), .Z(n3362) );
  HS65_LH_BFX4 U4154 ( .A(n3365), .Z(n3363) );
  HS65_LH_BFX4 U4155 ( .A(n3366), .Z(n3364) );
  HS65_LH_BFX4 U4156 ( .A(n3367), .Z(n3365) );
  HS65_LH_BFX4 U4157 ( .A(n3368), .Z(n3366) );
  HS65_LH_BFX4 U4158 ( .A(n3369), .Z(n3367) );
  HS65_LH_BFX4 U4159 ( .A(n3370), .Z(n3368) );
  HS65_LH_BFX4 U4160 ( .A(n3371), .Z(n3369) );
  HS65_LH_BFX4 U4161 ( .A(n3372), .Z(n3370) );
  HS65_LH_BFX4 U4162 ( .A(n3373), .Z(n3371) );
  HS65_LH_BFX4 U4163 ( .A(n3374), .Z(n3372) );
  HS65_LH_BFX4 U4164 ( .A(n3375), .Z(n3373) );
  HS65_LH_BFX4 U4165 ( .A(n3376), .Z(n3374) );
  HS65_LH_BFX4 U4166 ( .A(n3377), .Z(n3375) );
  HS65_LH_BFX4 U4167 ( .A(n3378), .Z(n3376) );
  HS65_LH_BFX4 U4168 ( .A(n3379), .Z(n3377) );
  HS65_LH_BFX4 U4169 ( .A(n3380), .Z(n3378) );
  HS65_LH_BFX4 U4170 ( .A(n3381), .Z(n3379) );
  HS65_LH_BFX4 U4171 ( .A(n3382), .Z(n3380) );
  HS65_LH_BFX4 U4172 ( .A(n3383), .Z(n3381) );
  HS65_LH_BFX4 U4173 ( .A(n3384), .Z(n3382) );
  HS65_LH_BFX4 U4174 ( .A(n3385), .Z(n3383) );
  HS65_LH_BFX4 U4175 ( .A(\u_DataPath/branch_target_i [14]), .Z(n3384) );
  HS65_LH_BFX4 U4176 ( .A(\u_DataPath/jump_address_i [14]), .Z(n3385) );
  HS65_LH_IVX13 U4177 ( .A(n13166), .Z(n13955) );
  HS65_LH_BFX4 U4178 ( .A(n14090), .Z(n3386) );
  HS65_LH_BFX4 U4179 ( .A(n3389), .Z(n3387) );
  HS65_LH_BFX4 U4180 ( .A(n3390), .Z(n3388) );
  HS65_LH_BFX4 U4181 ( .A(n3391), .Z(n3389) );
  HS65_LH_BFX4 U4182 ( .A(n3392), .Z(n3390) );
  HS65_LH_BFX4 U4183 ( .A(n3393), .Z(n3391) );
  HS65_LH_BFX4 U4184 ( .A(n3394), .Z(n3392) );
  HS65_LH_BFX4 U4185 ( .A(n3395), .Z(n3393) );
  HS65_LH_BFX4 U4186 ( .A(n3396), .Z(n3394) );
  HS65_LH_BFX4 U4187 ( .A(n3397), .Z(n3395) );
  HS65_LH_BFX4 U4188 ( .A(n3398), .Z(n3396) );
  HS65_LH_BFX4 U4189 ( .A(n3399), .Z(n3397) );
  HS65_LH_BFX4 U4190 ( .A(n3400), .Z(n3398) );
  HS65_LH_BFX4 U4191 ( .A(n3401), .Z(n3399) );
  HS65_LH_BFX4 U4192 ( .A(n3402), .Z(n3400) );
  HS65_LH_BFX4 U4193 ( .A(n3403), .Z(n3401) );
  HS65_LH_BFX4 U4194 ( .A(n3404), .Z(n3402) );
  HS65_LH_BFX4 U4195 ( .A(n3405), .Z(n3403) );
  HS65_LH_BFX4 U4196 ( .A(n3406), .Z(n3404) );
  HS65_LH_BFX4 U4197 ( .A(n3407), .Z(n3405) );
  HS65_LH_BFX4 U4198 ( .A(n3408), .Z(n3406) );
  HS65_LH_BFX4 U4199 ( .A(n3409), .Z(n3407) );
  HS65_LH_BFX4 U4200 ( .A(n3410), .Z(n3408) );
  HS65_LH_BFX4 U4201 ( .A(n3411), .Z(n3409) );
  HS65_LH_BFX4 U4202 ( .A(n3412), .Z(n3410) );
  HS65_LH_BFX4 U4203 ( .A(n3413), .Z(n3411) );
  HS65_LH_BFX4 U4204 ( .A(n3414), .Z(n3412) );
  HS65_LH_BFX4 U4205 ( .A(n3415), .Z(n3413) );
  HS65_LH_BFX4 U4206 ( .A(n3416), .Z(n3414) );
  HS65_LH_BFX4 U4207 ( .A(n3417), .Z(n3415) );
  HS65_LH_BFX4 U4208 ( .A(n3418), .Z(n3416) );
  HS65_LH_BFX4 U4209 ( .A(n3419), .Z(n3417) );
  HS65_LH_BFX4 U4210 ( .A(n3420), .Z(n3418) );
  HS65_LH_BFX4 U4211 ( .A(n3421), .Z(n3419) );
  HS65_LH_BFX4 U4212 ( .A(n3422), .Z(n3420) );
  HS65_LH_BFX4 U4213 ( .A(n3423), .Z(n3421) );
  HS65_LH_BFX4 U4214 ( .A(n3424), .Z(n3422) );
  HS65_LH_BFX4 U4215 ( .A(n3425), .Z(n3423) );
  HS65_LH_BFX4 U4216 ( .A(n3426), .Z(n3424) );
  HS65_LH_BFX4 U4217 ( .A(n3427), .Z(n3425) );
  HS65_LH_BFX4 U4218 ( .A(n3428), .Z(n3426) );
  HS65_LH_BFX4 U4219 ( .A(n3429), .Z(n3427) );
  HS65_LH_BFX4 U4220 ( .A(n3430), .Z(n3428) );
  HS65_LH_BFX4 U4221 ( .A(n3431), .Z(n3429) );
  HS65_LH_BFX4 U4222 ( .A(n3432), .Z(n3430) );
  HS65_LH_BFX4 U4223 ( .A(n3433), .Z(n3431) );
  HS65_LH_BFX4 U4224 ( .A(n3434), .Z(n3432) );
  HS65_LH_BFX4 U4225 ( .A(n3435), .Z(n3433) );
  HS65_LH_BFX4 U4226 ( .A(n3436), .Z(n3434) );
  HS65_LH_BFX4 U4227 ( .A(\u_DataPath/branch_target_i [15]), .Z(n3435) );
  HS65_LH_BFX4 U4228 ( .A(\u_DataPath/jump_address_i [15]), .Z(n3436) );
  HS65_LH_BFX4 U4229 ( .A(n3440), .Z(n3437) );
  HS65_LH_BFX4 U4231 ( .A(n3442), .Z(n3439) );
  HS65_LH_BFX4 U4232 ( .A(n3443), .Z(n3440) );
  HS65_LH_BFX4 U4233 ( .A(n13211), .Z(n3441) );
  HS65_LH_BFX4 U4234 ( .A(n3444), .Z(n3442) );
  HS65_LH_BFX4 U4235 ( .A(n3445), .Z(n3443) );
  HS65_LH_BFX4 U4236 ( .A(n3446), .Z(n3444) );
  HS65_LH_BFX4 U4237 ( .A(n3447), .Z(n3445) );
  HS65_LH_BFX4 U4238 ( .A(n3448), .Z(n3446) );
  HS65_LH_BFX4 U4239 ( .A(n3449), .Z(n3447) );
  HS65_LH_BFX4 U4240 ( .A(n3450), .Z(n3448) );
  HS65_LH_BFX4 U4241 ( .A(n3451), .Z(n3449) );
  HS65_LH_BFX4 U4242 ( .A(n3452), .Z(n3450) );
  HS65_LH_BFX4 U4243 ( .A(n3453), .Z(n3451) );
  HS65_LH_BFX4 U4244 ( .A(n3454), .Z(n3452) );
  HS65_LH_BFX4 U4245 ( .A(n3455), .Z(n3453) );
  HS65_LH_BFX4 U4246 ( .A(n3456), .Z(n3454) );
  HS65_LH_BFX4 U4247 ( .A(n3457), .Z(n3455) );
  HS65_LH_BFX4 U4248 ( .A(n3458), .Z(n3456) );
  HS65_LH_BFX4 U4249 ( .A(n3459), .Z(n3457) );
  HS65_LH_BFX4 U4250 ( .A(n3460), .Z(n3458) );
  HS65_LH_BFX4 U4251 ( .A(n3461), .Z(n3459) );
  HS65_LH_BFX4 U4252 ( .A(n3462), .Z(n3460) );
  HS65_LH_BFX4 U4253 ( .A(n3463), .Z(n3461) );
  HS65_LH_BFX4 U4254 ( .A(n3464), .Z(n3462) );
  HS65_LH_BFX4 U4255 ( .A(n3465), .Z(n3463) );
  HS65_LH_BFX4 U4256 ( .A(n3466), .Z(n3464) );
  HS65_LH_BFX4 U4257 ( .A(n3467), .Z(n3465) );
  HS65_LH_BFX4 U4258 ( .A(n3468), .Z(n3466) );
  HS65_LH_BFX4 U4259 ( .A(n3469), .Z(n3467) );
  HS65_LH_BFX4 U4260 ( .A(n3470), .Z(n3468) );
  HS65_LH_BFX4 U4261 ( .A(n3471), .Z(n3469) );
  HS65_LH_BFX4 U4262 ( .A(n3472), .Z(n3470) );
  HS65_LH_BFX4 U4263 ( .A(n3473), .Z(n3471) );
  HS65_LH_BFX4 U4264 ( .A(n3474), .Z(n3472) );
  HS65_LH_BFX4 U4265 ( .A(n3475), .Z(n3473) );
  HS65_LH_BFX4 U4266 ( .A(n3476), .Z(n3474) );
  HS65_LH_BFX4 U4267 ( .A(n3477), .Z(n3475) );
  HS65_LH_BFX4 U4268 ( .A(n3478), .Z(n3476) );
  HS65_LH_BFX4 U4269 ( .A(n3479), .Z(n3477) );
  HS65_LH_BFX4 U4270 ( .A(n3480), .Z(n3478) );
  HS65_LH_BFX4 U4271 ( .A(n3481), .Z(n3479) );
  HS65_LH_BFX4 U4272 ( .A(n3482), .Z(n3480) );
  HS65_LH_BFX4 U4273 ( .A(n3483), .Z(n3481) );
  HS65_LH_BFX4 U4274 ( .A(n3484), .Z(n3482) );
  HS65_LH_BFX4 U4275 ( .A(n3485), .Z(n3483) );
  HS65_LH_BFX4 U4276 ( .A(n3486), .Z(n3484) );
  HS65_LH_BFX4 U4277 ( .A(n3487), .Z(n3485) );
  HS65_LH_BFX4 U4278 ( .A(n3488), .Z(n3486) );
  HS65_LH_BFX4 U4279 ( .A(\u_DataPath/branch_target_i [16]), .Z(n3487) );
  HS65_LH_BFX4 U4280 ( .A(\u_DataPath/jump_address_i [16]), .Z(n3488) );
  HS65_LH_IVX13 U4281 ( .A(n13256), .Z(n13957) );
  HS65_LH_BFX4 U4282 ( .A(n14092), .Z(n3489) );
  HS65_LH_BFX4 U4283 ( .A(n3492), .Z(n3490) );
  HS65_LH_BFX4 U4284 ( .A(n3493), .Z(n3491) );
  HS65_LH_BFX4 U4285 ( .A(n3494), .Z(n3492) );
  HS65_LH_BFX4 U4286 ( .A(n3495), .Z(n3493) );
  HS65_LH_BFX4 U4287 ( .A(n3496), .Z(n3494) );
  HS65_LH_BFX4 U4288 ( .A(n3497), .Z(n3495) );
  HS65_LH_BFX4 U4289 ( .A(n3498), .Z(n3496) );
  HS65_LH_BFX4 U4290 ( .A(n3499), .Z(n3497) );
  HS65_LH_BFX4 U4291 ( .A(n3500), .Z(n3498) );
  HS65_LH_BFX4 U4292 ( .A(n3501), .Z(n3499) );
  HS65_LH_BFX4 U4293 ( .A(n3502), .Z(n3500) );
  HS65_LH_BFX4 U4294 ( .A(n3503), .Z(n3501) );
  HS65_LH_BFX4 U4295 ( .A(n3504), .Z(n3502) );
  HS65_LH_BFX4 U4296 ( .A(n3505), .Z(n3503) );
  HS65_LH_BFX4 U4297 ( .A(n3506), .Z(n3504) );
  HS65_LH_BFX4 U4298 ( .A(n3507), .Z(n3505) );
  HS65_LH_BFX4 U4299 ( .A(n3508), .Z(n3506) );
  HS65_LH_BFX4 U4300 ( .A(n3509), .Z(n3507) );
  HS65_LH_BFX4 U4301 ( .A(n3510), .Z(n3508) );
  HS65_LH_BFX4 U4302 ( .A(n3511), .Z(n3509) );
  HS65_LH_BFX4 U4303 ( .A(n3512), .Z(n3510) );
  HS65_LH_BFX4 U4304 ( .A(n3513), .Z(n3511) );
  HS65_LH_BFX4 U4305 ( .A(n3514), .Z(n3512) );
  HS65_LH_BFX4 U4306 ( .A(n3515), .Z(n3513) );
  HS65_LH_BFX4 U4307 ( .A(n3516), .Z(n3514) );
  HS65_LH_BFX4 U4308 ( .A(n3517), .Z(n3515) );
  HS65_LH_BFX4 U4309 ( .A(n3518), .Z(n3516) );
  HS65_LH_BFX4 U4310 ( .A(n3519), .Z(n3517) );
  HS65_LH_BFX4 U4311 ( .A(n3520), .Z(n3518) );
  HS65_LH_BFX4 U4312 ( .A(n3521), .Z(n3519) );
  HS65_LH_BFX4 U4313 ( .A(n3522), .Z(n3520) );
  HS65_LH_BFX4 U4314 ( .A(n3523), .Z(n3521) );
  HS65_LH_BFX4 U4315 ( .A(n3524), .Z(n3522) );
  HS65_LH_BFX4 U4316 ( .A(n3525), .Z(n3523) );
  HS65_LH_BFX4 U4317 ( .A(n3526), .Z(n3524) );
  HS65_LH_BFX4 U4318 ( .A(n3527), .Z(n3525) );
  HS65_LH_BFX4 U4319 ( .A(n3528), .Z(n3526) );
  HS65_LH_BFX4 U4320 ( .A(n3529), .Z(n3527) );
  HS65_LH_BFX4 U4321 ( .A(n3530), .Z(n3528) );
  HS65_LH_BFX4 U4322 ( .A(n3531), .Z(n3529) );
  HS65_LH_BFX4 U4323 ( .A(n3532), .Z(n3530) );
  HS65_LH_BFX4 U4324 ( .A(n3533), .Z(n3531) );
  HS65_LH_BFX4 U4325 ( .A(n3534), .Z(n3532) );
  HS65_LH_BFX4 U4326 ( .A(n3535), .Z(n3533) );
  HS65_LH_BFX4 U4327 ( .A(n3536), .Z(n3534) );
  HS65_LH_BFX4 U4328 ( .A(n3537), .Z(n3535) );
  HS65_LH_BFX4 U4329 ( .A(n3538), .Z(n3536) );
  HS65_LH_BFX4 U4330 ( .A(n3539), .Z(n3537) );
  HS65_LH_BFX4 U4331 ( .A(\u_DataPath/branch_target_i [17]), .Z(n3538) );
  HS65_LH_BFX4 U4332 ( .A(\u_DataPath/jump_address_i [17]), .Z(n3539) );
  HS65_LH_BFX4 U4333 ( .A(n3543), .Z(n3540) );
  HS65_LH_BFX4 U4335 ( .A(n3545), .Z(n3542) );
  HS65_LH_BFX4 U4336 ( .A(n3546), .Z(n3543) );
  HS65_LH_BFX4 U4338 ( .A(n3547), .Z(n3545) );
  HS65_LH_BFX4 U4339 ( .A(n3548), .Z(n3546) );
  HS65_LH_BFX4 U4340 ( .A(n3549), .Z(n3547) );
  HS65_LH_BFX4 U4341 ( .A(n3550), .Z(n3548) );
  HS65_LH_BFX4 U4342 ( .A(n3551), .Z(n3549) );
  HS65_LH_BFX4 U4343 ( .A(n3552), .Z(n3550) );
  HS65_LH_BFX4 U4344 ( .A(n3553), .Z(n3551) );
  HS65_LH_BFX4 U4345 ( .A(n3554), .Z(n3552) );
  HS65_LH_BFX4 U4346 ( .A(n3555), .Z(n3553) );
  HS65_LH_BFX4 U4347 ( .A(n3556), .Z(n3554) );
  HS65_LH_BFX4 U4348 ( .A(n3557), .Z(n3555) );
  HS65_LH_BFX4 U4349 ( .A(n3558), .Z(n3556) );
  HS65_LH_BFX4 U4350 ( .A(n3559), .Z(n3557) );
  HS65_LH_BFX4 U4351 ( .A(n3560), .Z(n3558) );
  HS65_LH_BFX4 U4352 ( .A(n3561), .Z(n3559) );
  HS65_LH_BFX4 U4353 ( .A(n3562), .Z(n3560) );
  HS65_LH_BFX4 U4354 ( .A(n3563), .Z(n3561) );
  HS65_LH_BFX4 U4355 ( .A(n3564), .Z(n3562) );
  HS65_LH_BFX4 U4356 ( .A(n3565), .Z(n3563) );
  HS65_LH_BFX4 U4357 ( .A(n3566), .Z(n3564) );
  HS65_LH_BFX4 U4358 ( .A(n3567), .Z(n3565) );
  HS65_LH_BFX4 U4359 ( .A(n3568), .Z(n3566) );
  HS65_LH_BFX4 U4360 ( .A(n3569), .Z(n3567) );
  HS65_LH_BFX4 U4361 ( .A(n3570), .Z(n3568) );
  HS65_LH_BFX4 U4362 ( .A(n3571), .Z(n3569) );
  HS65_LH_BFX4 U4363 ( .A(n3572), .Z(n3570) );
  HS65_LH_BFX4 U4364 ( .A(n3573), .Z(n3571) );
  HS65_LH_BFX4 U4365 ( .A(n3574), .Z(n3572) );
  HS65_LH_BFX4 U4366 ( .A(n3575), .Z(n3573) );
  HS65_LH_BFX4 U4367 ( .A(n3576), .Z(n3574) );
  HS65_LH_BFX4 U4368 ( .A(n3577), .Z(n3575) );
  HS65_LH_BFX4 U4369 ( .A(n3578), .Z(n3576) );
  HS65_LH_BFX4 U4370 ( .A(n3579), .Z(n3577) );
  HS65_LH_BFX4 U4371 ( .A(n3580), .Z(n3578) );
  HS65_LH_BFX4 U4372 ( .A(n3581), .Z(n3579) );
  HS65_LH_BFX4 U4373 ( .A(n3582), .Z(n3580) );
  HS65_LH_BFX4 U4374 ( .A(n3583), .Z(n3581) );
  HS65_LH_BFX4 U4375 ( .A(n3584), .Z(n3582) );
  HS65_LH_BFX4 U4376 ( .A(n3585), .Z(n3583) );
  HS65_LH_BFX4 U4377 ( .A(n3586), .Z(n3584) );
  HS65_LH_BFX4 U4378 ( .A(n3587), .Z(n3585) );
  HS65_LH_BFX4 U4379 ( .A(n3588), .Z(n3586) );
  HS65_LH_BFX4 U4380 ( .A(n3589), .Z(n3587) );
  HS65_LH_BFX4 U4381 ( .A(n3590), .Z(n3588) );
  HS65_LH_BFX4 U4382 ( .A(n3591), .Z(n3589) );
  HS65_LH_BFX4 U4383 ( .A(\u_DataPath/branch_target_i [18]), .Z(n3590) );
  HS65_LH_BFX4 U4384 ( .A(\u_DataPath/jump_address_i [18]), .Z(n3591) );
  HS65_LH_IVX13 U4385 ( .A(n11920), .Z(n13959) );
  HS65_LH_BFX4 U4386 ( .A(n14094), .Z(n3592) );
  HS65_LH_BFX4 U4387 ( .A(n3595), .Z(n3593) );
  HS65_LH_BFX4 U4388 ( .A(n3596), .Z(n3594) );
  HS65_LH_BFX4 U4389 ( .A(n3597), .Z(n3595) );
  HS65_LH_BFX4 U4390 ( .A(n3598), .Z(n3596) );
  HS65_LH_BFX4 U4391 ( .A(n3599), .Z(n3597) );
  HS65_LH_BFX4 U4392 ( .A(n3600), .Z(n3598) );
  HS65_LH_BFX4 U4393 ( .A(n3601), .Z(n3599) );
  HS65_LH_BFX4 U4394 ( .A(n3602), .Z(n3600) );
  HS65_LH_BFX4 U4395 ( .A(n3603), .Z(n3601) );
  HS65_LH_BFX4 U4396 ( .A(n3604), .Z(n3602) );
  HS65_LH_BFX4 U4397 ( .A(n3605), .Z(n3603) );
  HS65_LH_BFX4 U4398 ( .A(n3606), .Z(n3604) );
  HS65_LH_BFX4 U4399 ( .A(n3607), .Z(n3605) );
  HS65_LH_BFX4 U4400 ( .A(n3608), .Z(n3606) );
  HS65_LH_BFX4 U4401 ( .A(n3609), .Z(n3607) );
  HS65_LH_BFX4 U4402 ( .A(n3610), .Z(n3608) );
  HS65_LH_BFX4 U4403 ( .A(n3611), .Z(n3609) );
  HS65_LH_BFX4 U4404 ( .A(n3612), .Z(n3610) );
  HS65_LH_BFX4 U4405 ( .A(n3613), .Z(n3611) );
  HS65_LH_BFX4 U4406 ( .A(n3614), .Z(n3612) );
  HS65_LH_BFX4 U4407 ( .A(n3615), .Z(n3613) );
  HS65_LH_BFX4 U4408 ( .A(n3616), .Z(n3614) );
  HS65_LH_BFX4 U4409 ( .A(n3617), .Z(n3615) );
  HS65_LH_BFX4 U4410 ( .A(n3618), .Z(n3616) );
  HS65_LH_BFX4 U4411 ( .A(n3619), .Z(n3617) );
  HS65_LH_BFX4 U4412 ( .A(n3620), .Z(n3618) );
  HS65_LH_BFX4 U4413 ( .A(n3621), .Z(n3619) );
  HS65_LH_BFX4 U4414 ( .A(n3622), .Z(n3620) );
  HS65_LH_BFX4 U4415 ( .A(n3623), .Z(n3621) );
  HS65_LH_BFX4 U4416 ( .A(n3624), .Z(n3622) );
  HS65_LH_BFX4 U4417 ( .A(n3625), .Z(n3623) );
  HS65_LH_BFX4 U4418 ( .A(n3626), .Z(n3624) );
  HS65_LH_BFX4 U4419 ( .A(n3627), .Z(n3625) );
  HS65_LH_BFX4 U4420 ( .A(n3628), .Z(n3626) );
  HS65_LH_BFX4 U4421 ( .A(n3629), .Z(n3627) );
  HS65_LH_BFX4 U4422 ( .A(n3630), .Z(n3628) );
  HS65_LH_BFX4 U4423 ( .A(n3631), .Z(n3629) );
  HS65_LH_BFX4 U4424 ( .A(n3632), .Z(n3630) );
  HS65_LH_BFX4 U4425 ( .A(n3633), .Z(n3631) );
  HS65_LH_BFX4 U4426 ( .A(n3634), .Z(n3632) );
  HS65_LH_BFX4 U4427 ( .A(n3635), .Z(n3633) );
  HS65_LH_BFX4 U4428 ( .A(n3636), .Z(n3634) );
  HS65_LH_BFX4 U4429 ( .A(n3637), .Z(n3635) );
  HS65_LH_BFX4 U4430 ( .A(n3638), .Z(n3636) );
  HS65_LH_BFX4 U4431 ( .A(n3639), .Z(n3637) );
  HS65_LH_BFX4 U4432 ( .A(n3640), .Z(n3638) );
  HS65_LH_BFX4 U4433 ( .A(n3641), .Z(n3639) );
  HS65_LH_BFX4 U4434 ( .A(n3642), .Z(n3640) );
  HS65_LH_BFX4 U4435 ( .A(\u_DataPath/branch_target_i [19]), .Z(n3641) );
  HS65_LH_BFX4 U4436 ( .A(\u_DataPath/jump_address_i [19]), .Z(n3642) );
  HS65_LH_BFX4 U4437 ( .A(n3646), .Z(n3643) );
  HS65_LH_BFX4 U4439 ( .A(n3648), .Z(n3645) );
  HS65_LH_BFX4 U4440 ( .A(n3649), .Z(n3646) );
  HS65_LH_BFX4 U4442 ( .A(n3650), .Z(n3648) );
  HS65_LH_BFX4 U4443 ( .A(n3651), .Z(n3649) );
  HS65_LH_BFX4 U4444 ( .A(n3652), .Z(n3650) );
  HS65_LH_BFX4 U4445 ( .A(n3653), .Z(n3651) );
  HS65_LH_BFX4 U4446 ( .A(n3654), .Z(n3652) );
  HS65_LH_BFX4 U4447 ( .A(n3655), .Z(n3653) );
  HS65_LH_BFX4 U4448 ( .A(n3656), .Z(n3654) );
  HS65_LH_BFX4 U4449 ( .A(n3657), .Z(n3655) );
  HS65_LH_BFX4 U4450 ( .A(n3658), .Z(n3656) );
  HS65_LH_BFX4 U4451 ( .A(n3659), .Z(n3657) );
  HS65_LH_BFX4 U4452 ( .A(n3660), .Z(n3658) );
  HS65_LH_BFX4 U4453 ( .A(n3661), .Z(n3659) );
  HS65_LH_BFX4 U4454 ( .A(n3662), .Z(n3660) );
  HS65_LH_BFX4 U4455 ( .A(n3663), .Z(n3661) );
  HS65_LH_BFX4 U4456 ( .A(n3664), .Z(n3662) );
  HS65_LH_BFX4 U4457 ( .A(n3665), .Z(n3663) );
  HS65_LH_BFX4 U4458 ( .A(n3666), .Z(n3664) );
  HS65_LH_BFX4 U4459 ( .A(n3667), .Z(n3665) );
  HS65_LH_BFX4 U4460 ( .A(n3668), .Z(n3666) );
  HS65_LH_BFX4 U4461 ( .A(n3669), .Z(n3667) );
  HS65_LH_BFX4 U4462 ( .A(n3670), .Z(n3668) );
  HS65_LH_BFX4 U4463 ( .A(n3671), .Z(n3669) );
  HS65_LH_BFX4 U4464 ( .A(n3672), .Z(n3670) );
  HS65_LH_BFX4 U4465 ( .A(n3673), .Z(n3671) );
  HS65_LH_BFX4 U4466 ( .A(n3674), .Z(n3672) );
  HS65_LH_BFX4 U4467 ( .A(n3675), .Z(n3673) );
  HS65_LH_BFX4 U4468 ( .A(n3676), .Z(n3674) );
  HS65_LH_BFX4 U4469 ( .A(n3677), .Z(n3675) );
  HS65_LH_BFX4 U4470 ( .A(n3678), .Z(n3676) );
  HS65_LH_BFX4 U4471 ( .A(n3679), .Z(n3677) );
  HS65_LH_BFX4 U4472 ( .A(n3680), .Z(n3678) );
  HS65_LH_BFX4 U4473 ( .A(n3681), .Z(n3679) );
  HS65_LH_BFX4 U4474 ( .A(n3682), .Z(n3680) );
  HS65_LH_BFX4 U4475 ( .A(n3683), .Z(n3681) );
  HS65_LH_BFX4 U4476 ( .A(n3684), .Z(n3682) );
  HS65_LH_BFX4 U4477 ( .A(n3685), .Z(n3683) );
  HS65_LH_BFX4 U4478 ( .A(n3686), .Z(n3684) );
  HS65_LH_BFX4 U4479 ( .A(n3687), .Z(n3685) );
  HS65_LH_BFX4 U4480 ( .A(n3688), .Z(n3686) );
  HS65_LH_BFX4 U4481 ( .A(n3689), .Z(n3687) );
  HS65_LH_BFX4 U4482 ( .A(n3690), .Z(n3688) );
  HS65_LH_BFX4 U4483 ( .A(n3691), .Z(n3689) );
  HS65_LH_BFX4 U4484 ( .A(n3692), .Z(n3690) );
  HS65_LH_BFX4 U4485 ( .A(n3693), .Z(n3691) );
  HS65_LH_BFX4 U4486 ( .A(n3694), .Z(n3692) );
  HS65_LH_BFX4 U4487 ( .A(\u_DataPath/branch_target_i [20]), .Z(n3693) );
  HS65_LH_BFX4 U4488 ( .A(\u_DataPath/jump_address_i [20]), .Z(n3694) );
  HS65_LH_IVX13 U4489 ( .A(n12010), .Z(n13961) );
  HS65_LH_BFX4 U4490 ( .A(n14096), .Z(n3695) );
  HS65_LH_BFX4 U4491 ( .A(n3698), .Z(n3696) );
  HS65_LH_BFX4 U4492 ( .A(n3699), .Z(n3697) );
  HS65_LH_BFX4 U4493 ( .A(n3700), .Z(n3698) );
  HS65_LH_BFX4 U4494 ( .A(n3701), .Z(n3699) );
  HS65_LH_BFX4 U4495 ( .A(n3702), .Z(n3700) );
  HS65_LH_BFX4 U4496 ( .A(n3703), .Z(n3701) );
  HS65_LH_BFX4 U4497 ( .A(n3704), .Z(n3702) );
  HS65_LH_BFX4 U4498 ( .A(n3705), .Z(n3703) );
  HS65_LH_BFX4 U4499 ( .A(n3706), .Z(n3704) );
  HS65_LH_BFX4 U4500 ( .A(n3707), .Z(n3705) );
  HS65_LH_BFX4 U4501 ( .A(n3708), .Z(n3706) );
  HS65_LH_BFX4 U4502 ( .A(n3709), .Z(n3707) );
  HS65_LH_BFX4 U4503 ( .A(n3710), .Z(n3708) );
  HS65_LH_BFX4 U4504 ( .A(n3711), .Z(n3709) );
  HS65_LH_BFX4 U4505 ( .A(n3712), .Z(n3710) );
  HS65_LH_BFX4 U4506 ( .A(n3713), .Z(n3711) );
  HS65_LH_BFX4 U4507 ( .A(n3714), .Z(n3712) );
  HS65_LH_BFX4 U4508 ( .A(n3715), .Z(n3713) );
  HS65_LH_BFX4 U4509 ( .A(n3716), .Z(n3714) );
  HS65_LH_BFX4 U4510 ( .A(n3717), .Z(n3715) );
  HS65_LH_BFX4 U4511 ( .A(n3718), .Z(n3716) );
  HS65_LH_BFX4 U4512 ( .A(n3719), .Z(n3717) );
  HS65_LH_BFX4 U4513 ( .A(n3720), .Z(n3718) );
  HS65_LH_BFX4 U4514 ( .A(n3721), .Z(n3719) );
  HS65_LH_BFX4 U4515 ( .A(n3722), .Z(n3720) );
  HS65_LH_BFX4 U4516 ( .A(n3723), .Z(n3721) );
  HS65_LH_BFX4 U4517 ( .A(n3724), .Z(n3722) );
  HS65_LH_BFX4 U4518 ( .A(n3725), .Z(n3723) );
  HS65_LH_BFX4 U4519 ( .A(n3726), .Z(n3724) );
  HS65_LH_BFX4 U4520 ( .A(n3727), .Z(n3725) );
  HS65_LH_BFX4 U4521 ( .A(n3728), .Z(n3726) );
  HS65_LH_BFX4 U4522 ( .A(n3729), .Z(n3727) );
  HS65_LH_BFX4 U4523 ( .A(n3730), .Z(n3728) );
  HS65_LH_BFX4 U4524 ( .A(n3731), .Z(n3729) );
  HS65_LH_BFX4 U4525 ( .A(n3732), .Z(n3730) );
  HS65_LH_BFX4 U4526 ( .A(n3733), .Z(n3731) );
  HS65_LH_BFX4 U4527 ( .A(n3734), .Z(n3732) );
  HS65_LH_BFX4 U4528 ( .A(n3735), .Z(n3733) );
  HS65_LH_BFX4 U4529 ( .A(n3736), .Z(n3734) );
  HS65_LH_BFX4 U4530 ( .A(n3737), .Z(n3735) );
  HS65_LH_BFX4 U4531 ( .A(n3738), .Z(n3736) );
  HS65_LH_BFX4 U4532 ( .A(n3739), .Z(n3737) );
  HS65_LH_BFX4 U4533 ( .A(n3740), .Z(n3738) );
  HS65_LH_BFX4 U4534 ( .A(n3741), .Z(n3739) );
  HS65_LH_BFX4 U4535 ( .A(n3742), .Z(n3740) );
  HS65_LH_BFX4 U4536 ( .A(n3743), .Z(n3741) );
  HS65_LH_BFX4 U4537 ( .A(n3744), .Z(n3742) );
  HS65_LH_BFX4 U4538 ( .A(n3745), .Z(n3743) );
  HS65_LH_BFX4 U4539 ( .A(\u_DataPath/branch_target_i [21]), .Z(n3744) );
  HS65_LH_BFX4 U4540 ( .A(\u_DataPath/jump_address_i [21]), .Z(n3745) );
  HS65_LH_BFX4 U4541 ( .A(n3749), .Z(n3746) );
  HS65_LH_BFX4 U4543 ( .A(n3751), .Z(n3748) );
  HS65_LH_BFX4 U4544 ( .A(n3752), .Z(n3749) );
  HS65_LH_BFX4 U4546 ( .A(n3753), .Z(n3751) );
  HS65_LH_BFX4 U4547 ( .A(n3754), .Z(n3752) );
  HS65_LH_BFX4 U4548 ( .A(n3755), .Z(n3753) );
  HS65_LH_BFX4 U4549 ( .A(n3756), .Z(n3754) );
  HS65_LH_BFX4 U4550 ( .A(n3757), .Z(n3755) );
  HS65_LH_BFX4 U4551 ( .A(n3758), .Z(n3756) );
  HS65_LH_BFX4 U4552 ( .A(n3759), .Z(n3757) );
  HS65_LH_BFX4 U4553 ( .A(n3760), .Z(n3758) );
  HS65_LH_BFX4 U4554 ( .A(n3761), .Z(n3759) );
  HS65_LH_BFX4 U4555 ( .A(n3762), .Z(n3760) );
  HS65_LH_BFX4 U4556 ( .A(n3763), .Z(n3761) );
  HS65_LH_BFX4 U4557 ( .A(n3764), .Z(n3762) );
  HS65_LH_BFX4 U4558 ( .A(n3765), .Z(n3763) );
  HS65_LH_BFX4 U4559 ( .A(n3766), .Z(n3764) );
  HS65_LH_BFX4 U4560 ( .A(n3767), .Z(n3765) );
  HS65_LH_BFX4 U4561 ( .A(n3768), .Z(n3766) );
  HS65_LH_BFX4 U4562 ( .A(n3769), .Z(n3767) );
  HS65_LH_BFX4 U4563 ( .A(n3770), .Z(n3768) );
  HS65_LH_BFX4 U4564 ( .A(n3771), .Z(n3769) );
  HS65_LH_BFX4 U4565 ( .A(n3772), .Z(n3770) );
  HS65_LH_BFX4 U4566 ( .A(n3773), .Z(n3771) );
  HS65_LH_BFX4 U4567 ( .A(n3774), .Z(n3772) );
  HS65_LH_BFX4 U4568 ( .A(n3775), .Z(n3773) );
  HS65_LH_BFX4 U4569 ( .A(n3776), .Z(n3774) );
  HS65_LH_BFX4 U4570 ( .A(n3777), .Z(n3775) );
  HS65_LH_BFX4 U4571 ( .A(n3778), .Z(n3776) );
  HS65_LH_BFX4 U4572 ( .A(n3779), .Z(n3777) );
  HS65_LH_BFX4 U4573 ( .A(n3780), .Z(n3778) );
  HS65_LH_BFX4 U4574 ( .A(n3781), .Z(n3779) );
  HS65_LH_BFX4 U4575 ( .A(n3782), .Z(n3780) );
  HS65_LH_BFX4 U4576 ( .A(n3783), .Z(n3781) );
  HS65_LH_BFX4 U4577 ( .A(n3784), .Z(n3782) );
  HS65_LH_BFX4 U4578 ( .A(n3785), .Z(n3783) );
  HS65_LH_BFX4 U4579 ( .A(n3786), .Z(n3784) );
  HS65_LH_BFX4 U4580 ( .A(n3787), .Z(n3785) );
  HS65_LH_BFX4 U4581 ( .A(n3788), .Z(n3786) );
  HS65_LH_BFX4 U4582 ( .A(n3789), .Z(n3787) );
  HS65_LH_BFX4 U4583 ( .A(n3790), .Z(n3788) );
  HS65_LH_BFX4 U4584 ( .A(n3791), .Z(n3789) );
  HS65_LH_BFX4 U4585 ( .A(n3792), .Z(n3790) );
  HS65_LH_BFX4 U4586 ( .A(n3793), .Z(n3791) );
  HS65_LH_BFX4 U4587 ( .A(n3794), .Z(n3792) );
  HS65_LH_BFX4 U4588 ( .A(n3795), .Z(n3793) );
  HS65_LH_BFX4 U4589 ( .A(n3796), .Z(n3794) );
  HS65_LH_BFX4 U4590 ( .A(n3797), .Z(n3795) );
  HS65_LH_BFX4 U4591 ( .A(\u_DataPath/branch_target_i [22]), .Z(n3796) );
  HS65_LH_BFX4 U4592 ( .A(\u_DataPath/jump_address_i [22]), .Z(n3797) );
  HS65_LH_IVX13 U4593 ( .A(n12100), .Z(n13963) );
  HS65_LH_BFX4 U4594 ( .A(n14098), .Z(n3798) );
  HS65_LH_BFX4 U4595 ( .A(n3801), .Z(n3799) );
  HS65_LH_BFX4 U4596 ( .A(n3802), .Z(n3800) );
  HS65_LH_BFX4 U4597 ( .A(n3803), .Z(n3801) );
  HS65_LH_BFX4 U4598 ( .A(n3804), .Z(n3802) );
  HS65_LH_BFX4 U4599 ( .A(n3805), .Z(n3803) );
  HS65_LH_BFX4 U4600 ( .A(n3806), .Z(n3804) );
  HS65_LH_BFX4 U4601 ( .A(n3807), .Z(n3805) );
  HS65_LH_BFX4 U4602 ( .A(n3808), .Z(n3806) );
  HS65_LH_BFX4 U4603 ( .A(n3809), .Z(n3807) );
  HS65_LH_BFX4 U4604 ( .A(n3810), .Z(n3808) );
  HS65_LH_BFX4 U4605 ( .A(n3811), .Z(n3809) );
  HS65_LH_BFX4 U4606 ( .A(n3812), .Z(n3810) );
  HS65_LH_BFX4 U4607 ( .A(n3813), .Z(n3811) );
  HS65_LH_BFX4 U4608 ( .A(n3814), .Z(n3812) );
  HS65_LH_BFX4 U4609 ( .A(n3815), .Z(n3813) );
  HS65_LH_BFX4 U4610 ( .A(n3816), .Z(n3814) );
  HS65_LH_BFX4 U4611 ( .A(n3817), .Z(n3815) );
  HS65_LH_BFX4 U4612 ( .A(n3818), .Z(n3816) );
  HS65_LH_BFX4 U4613 ( .A(n3819), .Z(n3817) );
  HS65_LH_BFX4 U4614 ( .A(n3820), .Z(n3818) );
  HS65_LH_BFX4 U4615 ( .A(n3821), .Z(n3819) );
  HS65_LH_BFX4 U4616 ( .A(n3822), .Z(n3820) );
  HS65_LH_BFX4 U4617 ( .A(n3823), .Z(n3821) );
  HS65_LH_BFX4 U4618 ( .A(n3824), .Z(n3822) );
  HS65_LH_BFX4 U4619 ( .A(n3825), .Z(n3823) );
  HS65_LH_BFX4 U4620 ( .A(n3826), .Z(n3824) );
  HS65_LH_BFX4 U4621 ( .A(n3827), .Z(n3825) );
  HS65_LH_BFX4 U4622 ( .A(n3828), .Z(n3826) );
  HS65_LH_BFX4 U4623 ( .A(n3829), .Z(n3827) );
  HS65_LH_BFX4 U4624 ( .A(n3830), .Z(n3828) );
  HS65_LH_BFX4 U4625 ( .A(n3831), .Z(n3829) );
  HS65_LH_BFX4 U4626 ( .A(n3832), .Z(n3830) );
  HS65_LH_BFX4 U4627 ( .A(n3833), .Z(n3831) );
  HS65_LH_BFX4 U4628 ( .A(n3834), .Z(n3832) );
  HS65_LH_BFX4 U4629 ( .A(n3835), .Z(n3833) );
  HS65_LH_BFX4 U4630 ( .A(n3836), .Z(n3834) );
  HS65_LH_BFX4 U4631 ( .A(n3837), .Z(n3835) );
  HS65_LH_BFX4 U4632 ( .A(n3838), .Z(n3836) );
  HS65_LH_BFX4 U4633 ( .A(n3839), .Z(n3837) );
  HS65_LH_BFX4 U4634 ( .A(n3840), .Z(n3838) );
  HS65_LH_BFX4 U4635 ( .A(n3841), .Z(n3839) );
  HS65_LH_BFX4 U4636 ( .A(n3842), .Z(n3840) );
  HS65_LH_BFX4 U4637 ( .A(n3843), .Z(n3841) );
  HS65_LH_BFX4 U4638 ( .A(n3844), .Z(n3842) );
  HS65_LH_BFX4 U4639 ( .A(n3845), .Z(n3843) );
  HS65_LH_BFX4 U4640 ( .A(n3846), .Z(n3844) );
  HS65_LH_BFX4 U4641 ( .A(n3847), .Z(n3845) );
  HS65_LH_BFX4 U4642 ( .A(n3848), .Z(n3846) );
  HS65_LH_BFX4 U4643 ( .A(\u_DataPath/branch_target_i [23]), .Z(n3847) );
  HS65_LH_BFX4 U4644 ( .A(\u_DataPath/jump_address_i [23]), .Z(n3848) );
  HS65_LH_BFX4 U4645 ( .A(n3852), .Z(n3849) );
  HS65_LH_BFX4 U4647 ( .A(n3854), .Z(n3851) );
  HS65_LH_BFX4 U4648 ( .A(n3855), .Z(n3852) );
  HS65_LH_BFX4 U4650 ( .A(n3856), .Z(n3854) );
  HS65_LH_BFX4 U4651 ( .A(n3857), .Z(n3855) );
  HS65_LH_BFX4 U4652 ( .A(n3858), .Z(n3856) );
  HS65_LH_BFX4 U4653 ( .A(n3859), .Z(n3857) );
  HS65_LH_BFX4 U4654 ( .A(n3860), .Z(n3858) );
  HS65_LH_BFX4 U4655 ( .A(n3861), .Z(n3859) );
  HS65_LH_BFX4 U4656 ( .A(n3862), .Z(n3860) );
  HS65_LH_BFX4 U4657 ( .A(n3863), .Z(n3861) );
  HS65_LH_BFX4 U4658 ( .A(n3864), .Z(n3862) );
  HS65_LH_BFX4 U4659 ( .A(n3865), .Z(n3863) );
  HS65_LH_BFX4 U4660 ( .A(n3866), .Z(n3864) );
  HS65_LH_BFX4 U4661 ( .A(n3867), .Z(n3865) );
  HS65_LH_BFX4 U4662 ( .A(n3868), .Z(n3866) );
  HS65_LH_BFX4 U4663 ( .A(n3869), .Z(n3867) );
  HS65_LH_BFX4 U4664 ( .A(n3870), .Z(n3868) );
  HS65_LH_BFX4 U4665 ( .A(n3871), .Z(n3869) );
  HS65_LH_BFX4 U4666 ( .A(n3872), .Z(n3870) );
  HS65_LH_BFX4 U4667 ( .A(n3873), .Z(n3871) );
  HS65_LH_BFX4 U4668 ( .A(n3874), .Z(n3872) );
  HS65_LH_BFX4 U4669 ( .A(n3875), .Z(n3873) );
  HS65_LH_BFX4 U4670 ( .A(n3876), .Z(n3874) );
  HS65_LH_BFX4 U4671 ( .A(n3877), .Z(n3875) );
  HS65_LH_BFX4 U4672 ( .A(n3878), .Z(n3876) );
  HS65_LH_BFX4 U4673 ( .A(n3879), .Z(n3877) );
  HS65_LH_BFX4 U4674 ( .A(n3880), .Z(n3878) );
  HS65_LH_BFX4 U4675 ( .A(n3881), .Z(n3879) );
  HS65_LH_BFX4 U4676 ( .A(n3882), .Z(n3880) );
  HS65_LH_BFX4 U4677 ( .A(n3883), .Z(n3881) );
  HS65_LH_BFX4 U4678 ( .A(n3884), .Z(n3882) );
  HS65_LH_BFX4 U4679 ( .A(n3885), .Z(n3883) );
  HS65_LH_BFX4 U4680 ( .A(n3886), .Z(n3884) );
  HS65_LH_BFX4 U4681 ( .A(n3887), .Z(n3885) );
  HS65_LH_BFX4 U4682 ( .A(n3888), .Z(n3886) );
  HS65_LH_BFX4 U4683 ( .A(n3889), .Z(n3887) );
  HS65_LH_BFX4 U4684 ( .A(n3890), .Z(n3888) );
  HS65_LH_BFX4 U4685 ( .A(n3891), .Z(n3889) );
  HS65_LH_BFX4 U4686 ( .A(n3892), .Z(n3890) );
  HS65_LH_BFX4 U4687 ( .A(n3893), .Z(n3891) );
  HS65_LH_BFX4 U4688 ( .A(n3894), .Z(n3892) );
  HS65_LH_BFX4 U4689 ( .A(n3895), .Z(n3893) );
  HS65_LH_BFX4 U4690 ( .A(n3896), .Z(n3894) );
  HS65_LH_BFX4 U4691 ( .A(n3897), .Z(n3895) );
  HS65_LH_BFX4 U4692 ( .A(n3898), .Z(n3896) );
  HS65_LH_BFX4 U4693 ( .A(n3899), .Z(n3897) );
  HS65_LH_BFX4 U4694 ( .A(n3900), .Z(n3898) );
  HS65_LH_BFX4 U4695 ( .A(\u_DataPath/branch_target_i [24]), .Z(n3899) );
  HS65_LH_BFX4 U4696 ( .A(\u_DataPath/jump_address_i [24]), .Z(n3900) );
  HS65_LH_IVX13 U4697 ( .A(n12190), .Z(n13965) );
  HS65_LH_BFX4 U4698 ( .A(n14100), .Z(n3901) );
  HS65_LH_BFX4 U4699 ( .A(n3904), .Z(n3902) );
  HS65_LH_BFX4 U4700 ( .A(n3905), .Z(n3903) );
  HS65_LH_BFX4 U4701 ( .A(n3906), .Z(n3904) );
  HS65_LH_BFX4 U4702 ( .A(n3907), .Z(n3905) );
  HS65_LH_BFX4 U4703 ( .A(n3908), .Z(n3906) );
  HS65_LH_BFX4 U4704 ( .A(n3909), .Z(n3907) );
  HS65_LH_BFX4 U4705 ( .A(n3910), .Z(n3908) );
  HS65_LH_BFX4 U4706 ( .A(n3911), .Z(n3909) );
  HS65_LH_BFX4 U4707 ( .A(n3912), .Z(n3910) );
  HS65_LH_BFX4 U4708 ( .A(n3913), .Z(n3911) );
  HS65_LH_BFX4 U4709 ( .A(n3914), .Z(n3912) );
  HS65_LH_BFX4 U4710 ( .A(n3915), .Z(n3913) );
  HS65_LH_BFX4 U4711 ( .A(n3916), .Z(n3914) );
  HS65_LH_BFX4 U4712 ( .A(n3917), .Z(n3915) );
  HS65_LH_BFX4 U4713 ( .A(n3918), .Z(n3916) );
  HS65_LH_BFX4 U4714 ( .A(n3919), .Z(n3917) );
  HS65_LH_BFX4 U4715 ( .A(n3920), .Z(n3918) );
  HS65_LH_BFX4 U4716 ( .A(n3921), .Z(n3919) );
  HS65_LH_BFX4 U4717 ( .A(n3922), .Z(n3920) );
  HS65_LH_BFX4 U4718 ( .A(n3923), .Z(n3921) );
  HS65_LH_BFX4 U4719 ( .A(n3924), .Z(n3922) );
  HS65_LH_BFX4 U4720 ( .A(n3925), .Z(n3923) );
  HS65_LH_BFX4 U4721 ( .A(n3926), .Z(n3924) );
  HS65_LH_BFX4 U4722 ( .A(n3927), .Z(n3925) );
  HS65_LH_BFX4 U4723 ( .A(n3928), .Z(n3926) );
  HS65_LH_BFX4 U4724 ( .A(n3929), .Z(n3927) );
  HS65_LH_BFX4 U4725 ( .A(n3930), .Z(n3928) );
  HS65_LH_BFX4 U4726 ( .A(n3931), .Z(n3929) );
  HS65_LH_BFX4 U4727 ( .A(n3932), .Z(n3930) );
  HS65_LH_BFX4 U4728 ( .A(n3933), .Z(n3931) );
  HS65_LH_BFX4 U4729 ( .A(n3934), .Z(n3932) );
  HS65_LH_BFX4 U4730 ( .A(n3935), .Z(n3933) );
  HS65_LH_BFX4 U4731 ( .A(n3936), .Z(n3934) );
  HS65_LH_BFX4 U4732 ( .A(n3937), .Z(n3935) );
  HS65_LH_BFX4 U4733 ( .A(n3938), .Z(n3936) );
  HS65_LH_BFX4 U4734 ( .A(n3939), .Z(n3937) );
  HS65_LH_BFX4 U4735 ( .A(n3940), .Z(n3938) );
  HS65_LH_BFX4 U4736 ( .A(n3941), .Z(n3939) );
  HS65_LH_BFX4 U4737 ( .A(n3942), .Z(n3940) );
  HS65_LH_BFX4 U4738 ( .A(n3943), .Z(n3941) );
  HS65_LH_BFX4 U4739 ( .A(n3944), .Z(n3942) );
  HS65_LH_BFX4 U4740 ( .A(n3945), .Z(n3943) );
  HS65_LH_BFX4 U4741 ( .A(n3946), .Z(n3944) );
  HS65_LH_BFX4 U4742 ( .A(n3947), .Z(n3945) );
  HS65_LH_BFX4 U4743 ( .A(n3948), .Z(n3946) );
  HS65_LH_BFX4 U4744 ( .A(n3949), .Z(n3947) );
  HS65_LH_BFX4 U4745 ( .A(n3950), .Z(n3948) );
  HS65_LH_BFX4 U4746 ( .A(n3951), .Z(n3949) );
  HS65_LH_BFX4 U4747 ( .A(\u_DataPath/branch_target_i [25]), .Z(n3950) );
  HS65_LH_BFX4 U4748 ( .A(\u_DataPath/jump_address_i [25]), .Z(n3951) );
  HS65_LH_BFX4 U4749 ( .A(n3955), .Z(n3952) );
  HS65_LH_BFX4 U4751 ( .A(n3957), .Z(n3954) );
  HS65_LH_BFX4 U4752 ( .A(n3958), .Z(n3955) );
  HS65_LH_BFX4 U4754 ( .A(n3959), .Z(n3957) );
  HS65_LH_BFX4 U4755 ( .A(n3960), .Z(n3958) );
  HS65_LH_BFX4 U4756 ( .A(n3961), .Z(n3959) );
  HS65_LH_BFX4 U4757 ( .A(n3962), .Z(n3960) );
  HS65_LH_BFX4 U4758 ( .A(n3963), .Z(n3961) );
  HS65_LH_BFX4 U4759 ( .A(n3964), .Z(n3962) );
  HS65_LH_BFX4 U4760 ( .A(n3965), .Z(n3963) );
  HS65_LH_BFX4 U4761 ( .A(n3966), .Z(n3964) );
  HS65_LH_BFX4 U4762 ( .A(n3967), .Z(n3965) );
  HS65_LH_BFX4 U4763 ( .A(n3968), .Z(n3966) );
  HS65_LH_BFX4 U4764 ( .A(n3969), .Z(n3967) );
  HS65_LH_BFX4 U4765 ( .A(n3970), .Z(n3968) );
  HS65_LH_BFX4 U4766 ( .A(n3971), .Z(n3969) );
  HS65_LH_BFX4 U4767 ( .A(n3972), .Z(n3970) );
  HS65_LH_BFX4 U4768 ( .A(n3973), .Z(n3971) );
  HS65_LH_BFX4 U4769 ( .A(n3974), .Z(n3972) );
  HS65_LH_BFX4 U4770 ( .A(n3975), .Z(n3973) );
  HS65_LH_BFX4 U4771 ( .A(n3976), .Z(n3974) );
  HS65_LH_BFX4 U4772 ( .A(n3977), .Z(n3975) );
  HS65_LH_BFX4 U4773 ( .A(n3978), .Z(n3976) );
  HS65_LH_BFX4 U4774 ( .A(n3979), .Z(n3977) );
  HS65_LH_BFX4 U4775 ( .A(n3980), .Z(n3978) );
  HS65_LH_BFX4 U4776 ( .A(n3981), .Z(n3979) );
  HS65_LH_BFX4 U4777 ( .A(n3982), .Z(n3980) );
  HS65_LH_BFX4 U4778 ( .A(n3983), .Z(n3981) );
  HS65_LH_BFX4 U4779 ( .A(n3984), .Z(n3982) );
  HS65_LH_BFX4 U4780 ( .A(n3985), .Z(n3983) );
  HS65_LH_BFX4 U4781 ( .A(n3986), .Z(n3984) );
  HS65_LH_BFX4 U4782 ( .A(n3987), .Z(n3985) );
  HS65_LH_BFX4 U4783 ( .A(n3988), .Z(n3986) );
  HS65_LH_BFX4 U4784 ( .A(n3989), .Z(n3987) );
  HS65_LH_BFX4 U4785 ( .A(n3990), .Z(n3988) );
  HS65_LH_BFX4 U4786 ( .A(n3991), .Z(n3989) );
  HS65_LH_BFX4 U4787 ( .A(n3992), .Z(n3990) );
  HS65_LH_BFX4 U4788 ( .A(n3993), .Z(n3991) );
  HS65_LH_BFX4 U4789 ( .A(n3994), .Z(n3992) );
  HS65_LH_BFX4 U4790 ( .A(n3995), .Z(n3993) );
  HS65_LH_BFX4 U4791 ( .A(n3996), .Z(n3994) );
  HS65_LH_BFX4 U4792 ( .A(n3997), .Z(n3995) );
  HS65_LH_BFX4 U4793 ( .A(n3998), .Z(n3996) );
  HS65_LH_BFX4 U4794 ( .A(n3999), .Z(n3997) );
  HS65_LH_BFX4 U4795 ( .A(n4000), .Z(n3998) );
  HS65_LH_BFX4 U4796 ( .A(n4001), .Z(n3999) );
  HS65_LH_BFX4 U4797 ( .A(n4002), .Z(n4000) );
  HS65_LH_BFX4 U4798 ( .A(n4003), .Z(n4001) );
  HS65_LH_BFX4 U4799 ( .A(\u_DataPath/branch_target_i [26]), .Z(n4002) );
  HS65_LH_BFX4 U4800 ( .A(\u_DataPath/jump_address_i [26]), .Z(n4003) );
  HS65_LH_IVX13 U4801 ( .A(n13346), .Z(n13967) );
  HS65_LH_BFX4 U4802 ( .A(n14102), .Z(n4004) );
  HS65_LH_BFX4 U4803 ( .A(n4007), .Z(n4005) );
  HS65_LH_BFX4 U4804 ( .A(n4008), .Z(n4006) );
  HS65_LH_BFX4 U4805 ( .A(n4009), .Z(n4007) );
  HS65_LH_BFX4 U4806 ( .A(n4010), .Z(n4008) );
  HS65_LH_BFX4 U4807 ( .A(n4011), .Z(n4009) );
  HS65_LH_BFX4 U4808 ( .A(n4012), .Z(n4010) );
  HS65_LH_BFX4 U4809 ( .A(n4013), .Z(n4011) );
  HS65_LH_BFX4 U4810 ( .A(n4014), .Z(n4012) );
  HS65_LH_BFX4 U4811 ( .A(n4015), .Z(n4013) );
  HS65_LH_BFX4 U4812 ( .A(n4016), .Z(n4014) );
  HS65_LH_BFX4 U4813 ( .A(n4017), .Z(n4015) );
  HS65_LH_BFX4 U4814 ( .A(n4018), .Z(n4016) );
  HS65_LH_BFX4 U4815 ( .A(n4019), .Z(n4017) );
  HS65_LH_BFX4 U4816 ( .A(n4020), .Z(n4018) );
  HS65_LH_BFX4 U4817 ( .A(n4021), .Z(n4019) );
  HS65_LH_BFX4 U4818 ( .A(n4022), .Z(n4020) );
  HS65_LH_BFX4 U4819 ( .A(n4023), .Z(n4021) );
  HS65_LH_BFX4 U4820 ( .A(n4024), .Z(n4022) );
  HS65_LH_BFX4 U4821 ( .A(n4025), .Z(n4023) );
  HS65_LH_BFX4 U4822 ( .A(n4026), .Z(n4024) );
  HS65_LH_BFX4 U4823 ( .A(n4027), .Z(n4025) );
  HS65_LH_BFX4 U4824 ( .A(n4028), .Z(n4026) );
  HS65_LH_BFX4 U4825 ( .A(n4029), .Z(n4027) );
  HS65_LH_BFX4 U4826 ( .A(n4030), .Z(n4028) );
  HS65_LH_BFX4 U4827 ( .A(n4031), .Z(n4029) );
  HS65_LH_BFX4 U4828 ( .A(n4032), .Z(n4030) );
  HS65_LH_BFX4 U4829 ( .A(n4033), .Z(n4031) );
  HS65_LH_BFX4 U4830 ( .A(n4034), .Z(n4032) );
  HS65_LH_BFX4 U4831 ( .A(n4035), .Z(n4033) );
  HS65_LH_BFX4 U4832 ( .A(n4036), .Z(n4034) );
  HS65_LH_BFX4 U4833 ( .A(n4037), .Z(n4035) );
  HS65_LH_BFX4 U4834 ( .A(n4038), .Z(n4036) );
  HS65_LH_BFX4 U4835 ( .A(n4039), .Z(n4037) );
  HS65_LH_BFX4 U4836 ( .A(n4040), .Z(n4038) );
  HS65_LH_BFX4 U4837 ( .A(n4041), .Z(n4039) );
  HS65_LH_BFX4 U4838 ( .A(n4042), .Z(n4040) );
  HS65_LH_BFX4 U4839 ( .A(n4043), .Z(n4041) );
  HS65_LH_BFX4 U4840 ( .A(n4044), .Z(n4042) );
  HS65_LH_BFX4 U4841 ( .A(n4045), .Z(n4043) );
  HS65_LH_BFX4 U4842 ( .A(n4046), .Z(n4044) );
  HS65_LH_BFX4 U4843 ( .A(n4047), .Z(n4045) );
  HS65_LH_BFX4 U4844 ( .A(n4048), .Z(n4046) );
  HS65_LH_BFX4 U4845 ( .A(n4049), .Z(n4047) );
  HS65_LH_BFX4 U4846 ( .A(n4050), .Z(n4048) );
  HS65_LH_BFX4 U4847 ( .A(n4051), .Z(n4049) );
  HS65_LH_BFX4 U4848 ( .A(n4052), .Z(n4050) );
  HS65_LH_BFX4 U4849 ( .A(n4053), .Z(n4051) );
  HS65_LH_BFX4 U4850 ( .A(n4054), .Z(n4052) );
  HS65_LH_BFX4 U4851 ( .A(\u_DataPath/branch_target_i [27]), .Z(n4053) );
  HS65_LH_BFX4 U4852 ( .A(\u_DataPath/jump_address_i [27]), .Z(n4054) );
  HS65_LH_BFX4 U4853 ( .A(n4058), .Z(n4055) );
  HS65_LH_BFX4 U4855 ( .A(n4060), .Z(n4057) );
  HS65_LH_BFX4 U4856 ( .A(n4061), .Z(n4058) );
  HS65_LH_BFX4 U4858 ( .A(n4062), .Z(n4060) );
  HS65_LH_BFX4 U4859 ( .A(n4063), .Z(n4061) );
  HS65_LH_BFX4 U4860 ( .A(n4064), .Z(n4062) );
  HS65_LH_BFX4 U4861 ( .A(n4065), .Z(n4063) );
  HS65_LH_BFX4 U4862 ( .A(n4066), .Z(n4064) );
  HS65_LH_BFX4 U4863 ( .A(n4067), .Z(n4065) );
  HS65_LH_BFX4 U4864 ( .A(n4068), .Z(n4066) );
  HS65_LH_BFX4 U4865 ( .A(n4069), .Z(n4067) );
  HS65_LH_BFX4 U4866 ( .A(n4070), .Z(n4068) );
  HS65_LH_BFX4 U4867 ( .A(n4071), .Z(n4069) );
  HS65_LH_BFX4 U4868 ( .A(n4072), .Z(n4070) );
  HS65_LH_BFX4 U4869 ( .A(n4073), .Z(n4071) );
  HS65_LH_BFX4 U4870 ( .A(n4074), .Z(n4072) );
  HS65_LH_BFX4 U4871 ( .A(n4075), .Z(n4073) );
  HS65_LH_BFX4 U4872 ( .A(n4076), .Z(n4074) );
  HS65_LH_BFX4 U4873 ( .A(n4077), .Z(n4075) );
  HS65_LH_BFX4 U4874 ( .A(n4078), .Z(n4076) );
  HS65_LH_BFX4 U4875 ( .A(n4079), .Z(n4077) );
  HS65_LH_BFX4 U4876 ( .A(n4080), .Z(n4078) );
  HS65_LH_BFX4 U4877 ( .A(n4081), .Z(n4079) );
  HS65_LH_BFX4 U4878 ( .A(n4082), .Z(n4080) );
  HS65_LH_BFX4 U4879 ( .A(n4083), .Z(n4081) );
  HS65_LH_BFX4 U4880 ( .A(n4084), .Z(n4082) );
  HS65_LH_BFX4 U4881 ( .A(n4085), .Z(n4083) );
  HS65_LH_BFX4 U4882 ( .A(n4086), .Z(n4084) );
  HS65_LH_BFX4 U4883 ( .A(n4087), .Z(n4085) );
  HS65_LH_BFX4 U4884 ( .A(n4088), .Z(n4086) );
  HS65_LH_BFX4 U4885 ( .A(n4089), .Z(n4087) );
  HS65_LH_BFX4 U4886 ( .A(n4090), .Z(n4088) );
  HS65_LH_BFX4 U4887 ( .A(n4091), .Z(n4089) );
  HS65_LH_BFX4 U4888 ( .A(n4092), .Z(n4090) );
  HS65_LH_BFX4 U4889 ( .A(n4093), .Z(n4091) );
  HS65_LH_BFX4 U4890 ( .A(n4094), .Z(n4092) );
  HS65_LH_BFX4 U4891 ( .A(n4095), .Z(n4093) );
  HS65_LH_BFX4 U4892 ( .A(n4096), .Z(n4094) );
  HS65_LH_BFX4 U4893 ( .A(n4097), .Z(n4095) );
  HS65_LH_BFX4 U4894 ( .A(n4098), .Z(n4096) );
  HS65_LH_BFX4 U4895 ( .A(n4099), .Z(n4097) );
  HS65_LH_BFX4 U4896 ( .A(n4100), .Z(n4098) );
  HS65_LH_BFX4 U4897 ( .A(n4101), .Z(n4099) );
  HS65_LH_BFX4 U4898 ( .A(n4102), .Z(n4100) );
  HS65_LH_BFX4 U4899 ( .A(n4103), .Z(n4101) );
  HS65_LH_BFX4 U4900 ( .A(n4104), .Z(n4102) );
  HS65_LH_BFX4 U4901 ( .A(n4105), .Z(n4103) );
  HS65_LH_BFX4 U4902 ( .A(n4106), .Z(n4104) );
  HS65_LH_BFX4 U4903 ( .A(\u_DataPath/branch_target_i [28]), .Z(n4105) );
  HS65_LH_BFX4 U4904 ( .A(\u_DataPath/jump_address_i [28]), .Z(n4106) );
  HS65_LH_IVX13 U4905 ( .A(n13436), .Z(n13969) );
  HS65_LH_BFX4 U4906 ( .A(n14104), .Z(n4107) );
  HS65_LH_BFX4 U4907 ( .A(n4110), .Z(n4108) );
  HS65_LH_BFX4 U4908 ( .A(n4111), .Z(n4109) );
  HS65_LH_BFX4 U4909 ( .A(n4112), .Z(n4110) );
  HS65_LH_BFX4 U4910 ( .A(n4113), .Z(n4111) );
  HS65_LH_BFX4 U4911 ( .A(n4114), .Z(n4112) );
  HS65_LH_BFX4 U4912 ( .A(n4115), .Z(n4113) );
  HS65_LH_BFX4 U4913 ( .A(n4116), .Z(n4114) );
  HS65_LH_BFX4 U4914 ( .A(n4117), .Z(n4115) );
  HS65_LH_BFX4 U4915 ( .A(n4118), .Z(n4116) );
  HS65_LH_BFX4 U4916 ( .A(n4119), .Z(n4117) );
  HS65_LH_BFX4 U4917 ( .A(n4120), .Z(n4118) );
  HS65_LH_BFX4 U4918 ( .A(n4121), .Z(n4119) );
  HS65_LH_BFX4 U4919 ( .A(n4122), .Z(n4120) );
  HS65_LH_BFX4 U4920 ( .A(n4123), .Z(n4121) );
  HS65_LH_BFX4 U4921 ( .A(n4124), .Z(n4122) );
  HS65_LH_BFX4 U4922 ( .A(n4125), .Z(n4123) );
  HS65_LH_BFX4 U4923 ( .A(n4126), .Z(n4124) );
  HS65_LH_BFX4 U4924 ( .A(n4127), .Z(n4125) );
  HS65_LH_BFX4 U4925 ( .A(n4128), .Z(n4126) );
  HS65_LH_BFX4 U4926 ( .A(n4129), .Z(n4127) );
  HS65_LH_BFX4 U4927 ( .A(n4130), .Z(n4128) );
  HS65_LH_BFX4 U4928 ( .A(n4131), .Z(n4129) );
  HS65_LH_BFX4 U4929 ( .A(n4132), .Z(n4130) );
  HS65_LH_BFX4 U4930 ( .A(n4133), .Z(n4131) );
  HS65_LH_BFX4 U4931 ( .A(n4134), .Z(n4132) );
  HS65_LH_BFX4 U4932 ( .A(n4135), .Z(n4133) );
  HS65_LH_BFX4 U4933 ( .A(n4136), .Z(n4134) );
  HS65_LH_BFX4 U4934 ( .A(n4137), .Z(n4135) );
  HS65_LH_BFX4 U4935 ( .A(n4138), .Z(n4136) );
  HS65_LH_BFX4 U4936 ( .A(n4139), .Z(n4137) );
  HS65_LH_BFX4 U4937 ( .A(n4140), .Z(n4138) );
  HS65_LH_BFX4 U4938 ( .A(n4141), .Z(n4139) );
  HS65_LH_BFX4 U4939 ( .A(n4142), .Z(n4140) );
  HS65_LH_BFX4 U4940 ( .A(n4143), .Z(n4141) );
  HS65_LH_BFX4 U4941 ( .A(n4144), .Z(n4142) );
  HS65_LH_BFX4 U4942 ( .A(n4145), .Z(n4143) );
  HS65_LH_BFX4 U4943 ( .A(n4146), .Z(n4144) );
  HS65_LH_BFX4 U4944 ( .A(n4147), .Z(n4145) );
  HS65_LH_BFX4 U4945 ( .A(n4148), .Z(n4146) );
  HS65_LH_BFX4 U4946 ( .A(n4149), .Z(n4147) );
  HS65_LH_BFX4 U4947 ( .A(n4150), .Z(n4148) );
  HS65_LH_BFX4 U4948 ( .A(n4151), .Z(n4149) );
  HS65_LH_BFX4 U4949 ( .A(n4152), .Z(n4150) );
  HS65_LH_BFX4 U4950 ( .A(n4153), .Z(n4151) );
  HS65_LH_BFX4 U4951 ( .A(n4154), .Z(n4152) );
  HS65_LH_BFX4 U4952 ( .A(n4155), .Z(n4153) );
  HS65_LH_BFX4 U4953 ( .A(n4156), .Z(n4154) );
  HS65_LH_BFX4 U4954 ( .A(n4157), .Z(n4155) );
  HS65_LH_BFX4 U4955 ( .A(\u_DataPath/branch_target_i [29]), .Z(n4156) );
  HS65_LH_BFX4 U4956 ( .A(\u_DataPath/jump_address_i [29]), .Z(n4157) );
  HS65_LH_BFX4 U4957 ( .A(n4161), .Z(n4158) );
  HS65_LH_BFX4 U4959 ( .A(n4163), .Z(n4160) );
  HS65_LH_BFX4 U4960 ( .A(n4164), .Z(n4161) );
  HS65_LH_BFX4 U4962 ( .A(n4165), .Z(n4163) );
  HS65_LH_BFX4 U4963 ( .A(n4166), .Z(n4164) );
  HS65_LH_BFX4 U4964 ( .A(n4167), .Z(n4165) );
  HS65_LH_BFX4 U4965 ( .A(n4168), .Z(n4166) );
  HS65_LH_BFX4 U4966 ( .A(n4169), .Z(n4167) );
  HS65_LH_BFX4 U4967 ( .A(n4170), .Z(n4168) );
  HS65_LH_BFX4 U4968 ( .A(n4171), .Z(n4169) );
  HS65_LH_BFX4 U4969 ( .A(n4172), .Z(n4170) );
  HS65_LH_BFX4 U4970 ( .A(n4173), .Z(n4171) );
  HS65_LH_BFX4 U4971 ( .A(n4174), .Z(n4172) );
  HS65_LH_BFX4 U4972 ( .A(n4175), .Z(n4173) );
  HS65_LH_BFX4 U4973 ( .A(n4176), .Z(n4174) );
  HS65_LH_BFX4 U4974 ( .A(n4177), .Z(n4175) );
  HS65_LH_BFX4 U4975 ( .A(n4178), .Z(n4176) );
  HS65_LH_BFX4 U4976 ( .A(n4179), .Z(n4177) );
  HS65_LH_BFX4 U4977 ( .A(n4180), .Z(n4178) );
  HS65_LH_BFX4 U4978 ( .A(n4181), .Z(n4179) );
  HS65_LH_BFX4 U4979 ( .A(n4182), .Z(n4180) );
  HS65_LH_BFX4 U4980 ( .A(n4183), .Z(n4181) );
  HS65_LH_BFX4 U4981 ( .A(n4184), .Z(n4182) );
  HS65_LH_BFX4 U4982 ( .A(n4185), .Z(n4183) );
  HS65_LH_BFX4 U4983 ( .A(n4186), .Z(n4184) );
  HS65_LH_BFX4 U4984 ( .A(n4187), .Z(n4185) );
  HS65_LH_BFX4 U4985 ( .A(n4188), .Z(n4186) );
  HS65_LH_BFX4 U4986 ( .A(n4189), .Z(n4187) );
  HS65_LH_BFX4 U4987 ( .A(n4190), .Z(n4188) );
  HS65_LH_BFX4 U4988 ( .A(n4191), .Z(n4189) );
  HS65_LH_BFX4 U4989 ( .A(n4192), .Z(n4190) );
  HS65_LH_BFX4 U4990 ( .A(n4193), .Z(n4191) );
  HS65_LH_BFX4 U4991 ( .A(n4194), .Z(n4192) );
  HS65_LH_BFX4 U4992 ( .A(n4195), .Z(n4193) );
  HS65_LH_BFX4 U4993 ( .A(n4196), .Z(n4194) );
  HS65_LH_BFX4 U4994 ( .A(n4197), .Z(n4195) );
  HS65_LH_BFX4 U4995 ( .A(n4198), .Z(n4196) );
  HS65_LH_BFX4 U4996 ( .A(n4199), .Z(n4197) );
  HS65_LH_BFX4 U4997 ( .A(n4200), .Z(n4198) );
  HS65_LH_BFX4 U4998 ( .A(n4201), .Z(n4199) );
  HS65_LH_BFX4 U4999 ( .A(n4202), .Z(n4200) );
  HS65_LH_BFX4 U5000 ( .A(n4203), .Z(n4201) );
  HS65_LH_BFX4 U5001 ( .A(n4204), .Z(n4202) );
  HS65_LH_BFX4 U5002 ( .A(n4205), .Z(n4203) );
  HS65_LH_BFX4 U5003 ( .A(n4206), .Z(n4204) );
  HS65_LH_BFX4 U5004 ( .A(n4207), .Z(n4205) );
  HS65_LH_BFX4 U5005 ( .A(n4208), .Z(n4206) );
  HS65_LH_BFX4 U5006 ( .A(n4209), .Z(n4207) );
  HS65_LH_BFX4 U5007 ( .A(\u_DataPath/branch_target_i [30]), .Z(n4208) );
  HS65_LH_BFX4 U5008 ( .A(\u_DataPath/jump_address_i [30]), .Z(n4209) );
  HS65_LH_BFX4 U5009 ( .A(n4214), .Z(n4210) );
  HS65_LH_BFX4 U5010 ( .A(n4213), .Z(n4211) );
  HS65_LH_BFX4 U5011 ( .A(n4215), .Z(n4212) );
  HS65_LH_BFX4 U5012 ( .A(n4216), .Z(n4213) );
  HS65_LH_BFX4 U5013 ( .A(n4217), .Z(n4214) );
  HS65_LH_BFX4 U5014 ( .A(n4218), .Z(n4215) );
  HS65_LH_BFX4 U5015 ( .A(n4219), .Z(n4216) );
  HS65_LH_BFX4 U5016 ( .A(n4220), .Z(n4217) );
  HS65_LH_BFX4 U5017 ( .A(n4221), .Z(n4218) );
  HS65_LH_BFX4 U5018 ( .A(n4222), .Z(n4219) );
  HS65_LH_BFX4 U5019 ( .A(n4223), .Z(n4220) );
  HS65_LH_BFX4 U5020 ( .A(n4224), .Z(n4221) );
  HS65_LH_BFX4 U5021 ( .A(n4225), .Z(n4222) );
  HS65_LH_BFX4 U5022 ( .A(n4226), .Z(n4223) );
  HS65_LH_BFX4 U5023 ( .A(n4227), .Z(n4224) );
  HS65_LH_BFX4 U5024 ( .A(n4228), .Z(n4225) );
  HS65_LH_BFX4 U5025 ( .A(n4229), .Z(n4226) );
  HS65_LH_BFX4 U5026 ( .A(n4230), .Z(n4227) );
  HS65_LH_BFX4 U5027 ( .A(n4231), .Z(n4228) );
  HS65_LH_BFX4 U5028 ( .A(n4232), .Z(n4229) );
  HS65_LH_BFX4 U5029 ( .A(n4233), .Z(n4230) );
  HS65_LH_BFX4 U5030 ( .A(n4234), .Z(n4231) );
  HS65_LH_BFX4 U5031 ( .A(n12645), .Z(n4232) );
  HS65_LH_BFX4 U5032 ( .A(n4235), .Z(n4233) );
  HS65_LH_BFX4 U5033 ( .A(n4237), .Z(n4234) );
  HS65_LH_BFX4 U5034 ( .A(n4238), .Z(n4235) );
  HS65_LH_BFX4 U5035 ( .A(n17243), .Z(n4236) );
  HS65_LH_BFX4 U5036 ( .A(n4240), .Z(n4237) );
  HS65_LH_BFX4 U5037 ( .A(n4241), .Z(n4238) );
  HS65_LH_BFX4 U5038 ( .A(n14001), .Z(n4239) );
  HS65_LH_BFX4 U5039 ( .A(n4242), .Z(n4240) );
  HS65_LH_BFX4 U5040 ( .A(n4243), .Z(n4241) );
  HS65_LH_BFX4 U5041 ( .A(n4244), .Z(n4242) );
  HS65_LH_BFX4 U5042 ( .A(n4245), .Z(n4243) );
  HS65_LH_BFX4 U5043 ( .A(n4246), .Z(n4244) );
  HS65_LH_BFX4 U5044 ( .A(n4247), .Z(n4245) );
  HS65_LH_BFX4 U5045 ( .A(n4248), .Z(n4246) );
  HS65_LH_BFX4 U5046 ( .A(n4249), .Z(n4247) );
  HS65_LH_BFX4 U5047 ( .A(n4250), .Z(n4248) );
  HS65_LH_BFX4 U5048 ( .A(n4251), .Z(n4249) );
  HS65_LH_BFX4 U5049 ( .A(n4252), .Z(n4250) );
  HS65_LH_BFX4 U5050 ( .A(n4253), .Z(n4251) );
  HS65_LH_BFX4 U5051 ( .A(n4254), .Z(n4252) );
  HS65_LH_BFX4 U5052 ( .A(n4255), .Z(n4253) );
  HS65_LH_BFX4 U5053 ( .A(n4256), .Z(n4254) );
  HS65_LH_BFX4 U5054 ( .A(n4257), .Z(n4255) );
  HS65_LH_BFX4 U5055 ( .A(n4258), .Z(n4256) );
  HS65_LH_BFX4 U5056 ( .A(n4259), .Z(n4257) );
  HS65_LH_BFX4 U5057 ( .A(n4260), .Z(n4258) );
  HS65_LH_BFX4 U5058 ( .A(n4261), .Z(n4259) );
  HS65_LH_BFX4 U5059 ( .A(n4262), .Z(n4260) );
  HS65_LH_BFX4 U5060 ( .A(n4263), .Z(n4261) );
  HS65_LH_BFX4 U5061 ( .A(n4264), .Z(n4262) );
  HS65_LH_BFX4 U5062 ( .A(n4265), .Z(n4263) );
  HS65_LH_BFX4 U5063 ( .A(n4266), .Z(n4264) );
  HS65_LH_BFX4 U5064 ( .A(n4267), .Z(n4265) );
  HS65_LH_BFX4 U5065 ( .A(n4268), .Z(n4266) );
  HS65_LH_BFX4 U5066 ( .A(n4269), .Z(n4267) );
  HS65_LH_BFX4 U5067 ( .A(\u_DataPath/branch_target_i [3]), .Z(n4268) );
  HS65_LH_BFX4 U5068 ( .A(\u_DataPath/jump_address_i [3]), .Z(n4269) );
  HS65_LH_BFX4 U5070 ( .A(n4274), .Z(n4271) );
  HS65_LH_BFX4 U5071 ( .A(n4275), .Z(n4272) );
  HS65_LH_BFX4 U5072 ( .A(n17215), .Z(n4273) );
  HS65_LH_BFX4 U5073 ( .A(n4276), .Z(n4274) );
  HS65_LH_BFX4 U5074 ( .A(n4277), .Z(n4275) );
  HS65_LH_BFX4 U5075 ( .A(n4278), .Z(n4276) );
  HS65_LH_BFX4 U5076 ( .A(n4279), .Z(n4277) );
  HS65_LH_BFX4 U5077 ( .A(n4280), .Z(n4278) );
  HS65_LH_BFX4 U5078 ( .A(n4281), .Z(n4279) );
  HS65_LH_BFX4 U5079 ( .A(n4282), .Z(n4280) );
  HS65_LH_BFX4 U5080 ( .A(n4283), .Z(n4281) );
  HS65_LH_BFX4 U5081 ( .A(n4284), .Z(n4282) );
  HS65_LH_BFX4 U5082 ( .A(n4285), .Z(n4283) );
  HS65_LH_BFX4 U5083 ( .A(n4286), .Z(n4284) );
  HS65_LH_BFX4 U5084 ( .A(n4287), .Z(n4285) );
  HS65_LH_BFX4 U5085 ( .A(n4288), .Z(n4286) );
  HS65_LH_BFX4 U5086 ( .A(n4289), .Z(n4287) );
  HS65_LH_BFX4 U5087 ( .A(n4290), .Z(n4288) );
  HS65_LH_BFX4 U5088 ( .A(n4291), .Z(n4289) );
  HS65_LH_BFX4 U5089 ( .A(n4292), .Z(n4290) );
  HS65_LH_BFX4 U5090 ( .A(n4293), .Z(n4291) );
  HS65_LH_BFX4 U5091 ( .A(n4294), .Z(n4292) );
  HS65_LH_BFX4 U5092 ( .A(n4295), .Z(n4293) );
  HS65_LH_BFX4 U5093 ( .A(n4296), .Z(n4294) );
  HS65_LH_BFX4 U5094 ( .A(n4297), .Z(n4295) );
  HS65_LH_BFX4 U5095 ( .A(n4298), .Z(n4296) );
  HS65_LH_BFX4 U5096 ( .A(n4299), .Z(n4297) );
  HS65_LH_BFX4 U5097 ( .A(n4300), .Z(n4298) );
  HS65_LH_BFX4 U5098 ( .A(n4301), .Z(n4299) );
  HS65_LH_BFX4 U5099 ( .A(n4302), .Z(n4300) );
  HS65_LH_BFX4 U5100 ( .A(n4303), .Z(n4301) );
  HS65_LH_BFX4 U5101 ( .A(n4304), .Z(n4302) );
  HS65_LH_BFX4 U5102 ( .A(n4305), .Z(n4303) );
  HS65_LH_BFX4 U5103 ( .A(n4306), .Z(n4304) );
  HS65_LH_BFX4 U5104 ( .A(n4307), .Z(n4305) );
  HS65_LH_BFX4 U5105 ( .A(n4308), .Z(n4306) );
  HS65_LH_BFX4 U5106 ( .A(n4309), .Z(n4307) );
  HS65_LH_BFX4 U5107 ( .A(n4310), .Z(n4308) );
  HS65_LH_BFX4 U5108 ( .A(n4311), .Z(n4309) );
  HS65_LH_BFX4 U5109 ( .A(n4312), .Z(n4310) );
  HS65_LH_BFX4 U5110 ( .A(n4313), .Z(n4311) );
  HS65_LH_BFX4 U5111 ( .A(n4314), .Z(n4312) );
  HS65_LH_BFX4 U5112 ( .A(n4315), .Z(n4313) );
  HS65_LH_BFX4 U5113 ( .A(n4316), .Z(n4314) );
  HS65_LH_BFX4 U5114 ( .A(n4317), .Z(n4315) );
  HS65_LH_BFX4 U5115 ( .A(n4318), .Z(n4316) );
  HS65_LH_BFX4 U5116 ( .A(n4319), .Z(n4317) );
  HS65_LH_BFX4 U5117 ( .A(n4320), .Z(n4318) );
  HS65_LH_BFX4 U5118 ( .A(n4321), .Z(n4319) );
  HS65_LH_BFX4 U5119 ( .A(\u_DataPath/branch_target_i [31]), .Z(n4320) );
  HS65_LH_BFX4 U5120 ( .A(\u_DataPath/jump_address_i [31]), .Z(n4321) );
  HS65_LH_IVX13 U5121 ( .A(n12717), .Z(n13945) );
  HS65_LH_BFX4 U5122 ( .A(n14079), .Z(n4322) );
  HS65_LH_BFX4 U5123 ( .A(n4325), .Z(n4323) );
  HS65_LH_BFX4 U5124 ( .A(n4326), .Z(n4324) );
  HS65_LH_BFX4 U5125 ( .A(n4327), .Z(n4325) );
  HS65_LH_BFX4 U5126 ( .A(n4328), .Z(n4326) );
  HS65_LH_BFX4 U5127 ( .A(n4329), .Z(n4327) );
  HS65_LH_BFX4 U5128 ( .A(n4330), .Z(n4328) );
  HS65_LH_BFX4 U5129 ( .A(n4331), .Z(n4329) );
  HS65_LH_BFX4 U5130 ( .A(n4332), .Z(n4330) );
  HS65_LH_BFX4 U5131 ( .A(n4333), .Z(n4331) );
  HS65_LH_BFX4 U5132 ( .A(n4334), .Z(n4332) );
  HS65_LH_BFX4 U5133 ( .A(n4335), .Z(n4333) );
  HS65_LH_BFX4 U5134 ( .A(n4336), .Z(n4334) );
  HS65_LH_BFX4 U5135 ( .A(n4337), .Z(n4335) );
  HS65_LH_BFX4 U5136 ( .A(n4338), .Z(n4336) );
  HS65_LH_BFX4 U5137 ( .A(n4339), .Z(n4337) );
  HS65_LH_BFX4 U5138 ( .A(n4340), .Z(n4338) );
  HS65_LH_BFX4 U5139 ( .A(n4341), .Z(n4339) );
  HS65_LH_BFX4 U5140 ( .A(n4342), .Z(n4340) );
  HS65_LH_BFX4 U5141 ( .A(n4343), .Z(n4341) );
  HS65_LH_BFX4 U5142 ( .A(n4344), .Z(n4342) );
  HS65_LH_BFX4 U5143 ( .A(n4345), .Z(n4343) );
  HS65_LH_BFX4 U5144 ( .A(n4346), .Z(n4344) );
  HS65_LH_BFX4 U5145 ( .A(n4347), .Z(n4345) );
  HS65_LH_BFX4 U5146 ( .A(n4348), .Z(n4346) );
  HS65_LH_BFX4 U5147 ( .A(n4349), .Z(n4347) );
  HS65_LH_BFX4 U5148 ( .A(n4350), .Z(n4348) );
  HS65_LH_BFX4 U5149 ( .A(n4351), .Z(n4349) );
  HS65_LH_BFX4 U5150 ( .A(n4352), .Z(n4350) );
  HS65_LH_BFX4 U5151 ( .A(n4353), .Z(n4351) );
  HS65_LH_BFX4 U5152 ( .A(n4354), .Z(n4352) );
  HS65_LH_BFX4 U5153 ( .A(n4355), .Z(n4353) );
  HS65_LH_BFX4 U5154 ( .A(n4356), .Z(n4354) );
  HS65_LH_BFX4 U5155 ( .A(n4357), .Z(n4355) );
  HS65_LH_BFX4 U5156 ( .A(n4358), .Z(n4356) );
  HS65_LH_BFX4 U5157 ( .A(n4359), .Z(n4357) );
  HS65_LH_BFX4 U5158 ( .A(n4360), .Z(n4358) );
  HS65_LH_BFX4 U5159 ( .A(n4361), .Z(n4359) );
  HS65_LH_BFX4 U5160 ( .A(n4362), .Z(n4360) );
  HS65_LH_BFX4 U5161 ( .A(n4363), .Z(n4361) );
  HS65_LH_BFX4 U5162 ( .A(n4364), .Z(n4362) );
  HS65_LH_BFX4 U5163 ( .A(n4365), .Z(n4363) );
  HS65_LH_BFX4 U5164 ( .A(n4366), .Z(n4364) );
  HS65_LH_BFX4 U5165 ( .A(n4367), .Z(n4365) );
  HS65_LH_BFX4 U5166 ( .A(n4368), .Z(n4366) );
  HS65_LH_BFX4 U5167 ( .A(n4369), .Z(n4367) );
  HS65_LH_BFX4 U5168 ( .A(n4370), .Z(n4368) );
  HS65_LH_BFX4 U5169 ( .A(n4371), .Z(n4369) );
  HS65_LH_BFX4 U5170 ( .A(n4372), .Z(n4370) );
  HS65_LH_BFX4 U5171 ( .A(\u_DataPath/branch_target_i [5]), .Z(n4371) );
  HS65_LH_BFX4 U5172 ( .A(\u_DataPath/jump_address_i [5]), .Z(n4372) );
  HS65_LH_BFX4 U5174 ( .A(n15136), .Z(n4374) );
  HS65_LH_BFX4 U5176 ( .A(n4374), .Z(n4376) );
  HS65_LH_BFX4 U5193 ( .A(n4395), .Z(n4393) );
  HS65_LH_BFX4 U5195 ( .A(n4397), .Z(n4395) );
  HS65_LH_BFX4 U5197 ( .A(n4399), .Z(n4397) );
  HS65_LH_BFX4 U5199 ( .A(n4401), .Z(n4399) );
  HS65_LH_BFX4 U5201 ( .A(n4403), .Z(n4401) );
  HS65_LH_BFX4 U5203 ( .A(n4405), .Z(n4403) );
  HS65_LH_BFX4 U5205 ( .A(n4407), .Z(n4405) );
  HS65_LH_BFX4 U5207 ( .A(n4409), .Z(n4407) );
  HS65_LH_BFX4 U5209 ( .A(n4414), .Z(n4409) );
  HS65_LH_BFX4 U5211 ( .A(n4413), .Z(n4411) );
  HS65_LH_BFX4 U5213 ( .A(\u_DataPath/u_idexreg/N31 ), .Z(n4413) );
  HS65_LH_BFX4 U5214 ( .A(n14112), .Z(n4414) );
  HS65_LH_BFX4 U5277 ( .A(\u_DataPath/data_read_ex_1_i [18]), .Z(n4477) );
  HS65_LH_BFX4 U5343 ( .A(\u_DataPath/data_read_ex_1_i [17]), .Z(n4543) );
  HS65_LH_BFX4 U5410 ( .A(\u_DataPath/data_read_ex_1_i [16]), .Z(n4610) );
  HS65_LH_BFX4 U5536 ( .A(n4738), .Z(n4736) );
  HS65_LH_BFX4 U5537 ( .A(\u_DataPath/data_read_ex_1_i [8]), .Z(n4737) );
  HS65_LH_BFX4 U5538 ( .A(n4739), .Z(n4738) );
  HS65_LH_BFX4 U5539 ( .A(n4740), .Z(n4739) );
  HS65_LH_BFX4 U5540 ( .A(n4741), .Z(n4740) );
  HS65_LH_BFX4 U5541 ( .A(n14156), .Z(n4741) );
  HS65_LH_BFX4 U5604 ( .A(\u_DataPath/data_read_ex_1_i [22]), .Z(n4804) );
  HS65_LH_BFX4 U5668 ( .A(\u_DataPath/data_read_ex_1_i [28]), .Z(n4868) );
  HS65_LH_BFX4 U5735 ( .A(\u_DataPath/data_read_ex_1_i [24]), .Z(n4935) );
  HS65_LH_BFX4 U5801 ( .A(\u_DataPath/data_read_ex_1_i [9]), .Z(n5001) );
  HS65_LH_BFX4 U5803 ( .A(n5004), .Z(n5003) );
  HS65_LH_BFX4 U5804 ( .A(n14168), .Z(n5004) );
  HS65_LH_BFX4 U5867 ( .A(\u_DataPath/data_read_ex_1_i [25]), .Z(n5067) );
  HS65_LH_BFX4 U5916 ( .A(n5118), .Z(n5116) );
  HS65_LH_BFX4 U5918 ( .A(n5120), .Z(n5118) );
  HS65_LH_BFX4 U5920 ( .A(n5122), .Z(n5120) );
  HS65_LH_BFX4 U5922 ( .A(n5124), .Z(n5122) );
  HS65_LH_BFX4 U5924 ( .A(n5126), .Z(n5124) );
  HS65_LH_BFX4 U5926 ( .A(n5128), .Z(n5126) );
  HS65_LH_BFX4 U5928 ( .A(n5130), .Z(n5128) );
  HS65_LH_BFX4 U5930 ( .A(n5132), .Z(n5130) );
  HS65_LH_BFX4 U5932 ( .A(n5134), .Z(n5132) );
  HS65_LH_BFX4 U5933 ( .A(\u_DataPath/data_read_ex_1_i [5]), .Z(n5133) );
  HS65_LH_BFX4 U5934 ( .A(n5135), .Z(n5134) );
  HS65_LH_BFX4 U5935 ( .A(n5136), .Z(n5135) );
  HS65_LH_BFX4 U5936 ( .A(n14174), .Z(n5136) );
  HS65_LH_BFX4 U5975 ( .A(\u_DataPath/data_read_ex_1_i [21]), .Z(n5175) );
  HS65_LH_CNIVX3 U6033 ( .A(\u_DataPath/u_idexreg/N56 ), .Z(n5233) );
  HS65_LH_CNIVX3 U6034 ( .A(n5233), .Z(n5234) );
  HS65_LH_BFX4 U6108 ( .A(\u_DataPath/data_read_ex_1_i [13]), .Z(n5308) );
  HS65_LH_BFX4 U6167 ( .A(n5369), .Z(n5367) );
  HS65_LH_BFX4 U6169 ( .A(n5371), .Z(n5369) );
  HS65_LH_BFX4 U6171 ( .A(n5373), .Z(n5371) );
  HS65_LH_BFX4 U6173 ( .A(n5375), .Z(n5373) );
  HS65_LH_BFX4 U6174 ( .A(\u_DataPath/data_read_ex_1_i [7]), .Z(n5374) );
  HS65_LH_BFX4 U6175 ( .A(n5376), .Z(n5375) );
  HS65_LH_BFX4 U6176 ( .A(n5377), .Z(n5376) );
  HS65_LH_BFX4 U6177 ( .A(n14186), .Z(n5377) );
  HS65_LH_BFX4 U6307 ( .A(\u_DataPath/u_idexreg/N56 ), .Z(n5507) );
  HS65_LH_BFX4 U6371 ( .A(\u_DataPath/data_read_ex_1_i [23]), .Z(n5571) );
  HS65_LH_BFX4 U6503 ( .A(\u_DataPath/data_read_ex_1_i [10]), .Z(n5703) );
  HS65_LH_BFX4 U6569 ( .A(\u_DataPath/data_read_ex_1_i [19]), .Z(n5769) );
  HS65_LH_BFX4 U6635 ( .A(\u_DataPath/data_read_ex_1_i [11]), .Z(n5835) );
  HS65_LH_BFX4 U6701 ( .A(\u_DataPath/data_read_ex_1_i [27]), .Z(n5901) );
  HS65_LH_BFX4 U6705 ( .A(n5906), .Z(n5905) );
  HS65_LH_BFX4 U6706 ( .A(n5907), .Z(n5906) );
  HS65_LH_BFX4 U6707 ( .A(n5908), .Z(n5907) );
  HS65_LH_BFX4 U6708 ( .A(n5909), .Z(n5908) );
  HS65_LH_BFX4 U6709 ( .A(n5910), .Z(n5909) );
  HS65_LH_BFX4 U6710 ( .A(n5911), .Z(n5910) );
  HS65_LH_BFX4 U6711 ( .A(n5912), .Z(n5911) );
  HS65_LH_BFX4 U6712 ( .A(n5913), .Z(n5912) );
  HS65_LH_BFX4 U6713 ( .A(n5914), .Z(n5913) );
  HS65_LH_BFX4 U6714 ( .A(n5915), .Z(n5914) );
  HS65_LH_BFX4 U6715 ( .A(n5916), .Z(n5915) );
  HS65_LH_BFX4 U6716 ( .A(n5917), .Z(n5916) );
  HS65_LH_BFX4 U6717 ( .A(n5918), .Z(n5917) );
  HS65_LH_BFX4 U6718 ( .A(n5919), .Z(n5918) );
  HS65_LH_BFX4 U6719 ( .A(n5920), .Z(n5919) );
  HS65_LH_BFX4 U6720 ( .A(n5921), .Z(n5920) );
  HS65_LH_BFX4 U6721 ( .A(n5922), .Z(n5921) );
  HS65_LH_BFX4 U6722 ( .A(n5923), .Z(n5922) );
  HS65_LH_BFX4 U6723 ( .A(n5924), .Z(n5923) );
  HS65_LH_BFX4 U6724 ( .A(n14209), .Z(n5924) );
  HS65_LH_BFX4 U6750 ( .A(n5953), .Z(n5950) );
  HS65_LH_BFX4 U6753 ( .A(n5956), .Z(n5953) );
  HS65_LH_BFX4 U6756 ( .A(n5959), .Z(n5956) );
  HS65_LH_BFX4 U6758 ( .A(\u_DataPath/u_idexreg/N184 ), .Z(n5958) );
  HS65_LH_BFX4 U6759 ( .A(n5962), .Z(n5959) );
  HS65_LH_BFX4 U6762 ( .A(n5965), .Z(n5962) );
  HS65_LH_BFX4 U6765 ( .A(n5968), .Z(n5965) );
  HS65_LH_BFX4 U6768 ( .A(n5971), .Z(n5968) );
  HS65_LH_BFX4 U6771 ( .A(n5974), .Z(n5971) );
  HS65_LH_BFX4 U6774 ( .A(n5977), .Z(n5974) );
  HS65_LH_BFX4 U6777 ( .A(n5980), .Z(n5977) );
  HS65_LH_BFX4 U6780 ( .A(n5983), .Z(n5980) );
  HS65_LH_BFX4 U6783 ( .A(n5986), .Z(n5983) );
  HS65_LH_BFX4 U6786 ( .A(n5989), .Z(n5986) );
  HS65_LH_BFX4 U6789 ( .A(n5992), .Z(n5989) );
  HS65_LH_BFX4 U6792 ( .A(n5995), .Z(n5992) );
  HS65_LH_BFX4 U6795 ( .A(n5998), .Z(n5995) );
  HS65_LH_BFX4 U6798 ( .A(n6001), .Z(n5998) );
  HS65_LH_BFX4 U6801 ( .A(n6004), .Z(n6001) );
  HS65_LH_BFX4 U6804 ( .A(n6007), .Z(n6004) );
  HS65_LH_BFX4 U6807 ( .A(n6009), .Z(n6007) );
  HS65_LH_BFX4 U6809 ( .A(n6011), .Z(n6009) );
  HS65_LH_BFX4 U6811 ( .A(n6012), .Z(n6011) );
  HS65_LH_BFX4 U6812 ( .A(n6013), .Z(n6012) );
  HS65_LH_BFX4 U6813 ( .A(n6014), .Z(n6013) );
  HS65_LH_BFX4 U6814 ( .A(\u_DataPath/u_idexreg/N36 ), .Z(n6014) );
  HS65_LH_BFX4 U6841 ( .A(n14338), .Z(n6041) );
  HS65_LH_BFX4 U6899 ( .A(n6100), .Z(n6099) );
  HS65_LH_BFX4 U6900 ( .A(n6101), .Z(n6100) );
  HS65_LH_BFX4 U6901 ( .A(n6102), .Z(n6101) );
  HS65_LH_BFX4 U6902 ( .A(n6103), .Z(n6102) );
  HS65_LH_BFX4 U6903 ( .A(\u_DataPath/data_read_ex_2_i [14]), .Z(n6103) );
  HS65_LH_BFX4 U6931 ( .A(n6133), .Z(n6131) );
  HS65_LH_BFX4 U6933 ( .A(n6135), .Z(n6133) );
  HS65_LH_BFX4 U6935 ( .A(n6137), .Z(n6135) );
  HS65_LH_BFX4 U6937 ( .A(n6139), .Z(n6137) );
  HS65_LH_BFX4 U6939 ( .A(n6221), .Z(n6139) );
  HS65_LH_BFX4 U6945 ( .A(n6146), .Z(n6145) );
  HS65_LH_BFX4 U6946 ( .A(n6147), .Z(n6146) );
  HS65_LH_BFX4 U6947 ( .A(n6148), .Z(n6147) );
  HS65_LH_BFX4 U6948 ( .A(n6149), .Z(n6148) );
  HS65_LH_BFX4 U6949 ( .A(n6150), .Z(n6149) );
  HS65_LH_BFX4 U6950 ( .A(n6151), .Z(n6150) );
  HS65_LH_BFX4 U6951 ( .A(n6152), .Z(n6151) );
  HS65_LH_BFX4 U6952 ( .A(n6153), .Z(n6152) );
  HS65_LH_BFX4 U6953 ( .A(n6154), .Z(n6153) );
  HS65_LH_BFX4 U6954 ( .A(n6155), .Z(n6154) );
  HS65_LH_BFX4 U6955 ( .A(n6156), .Z(n6155) );
  HS65_LH_BFX4 U6956 ( .A(n6157), .Z(n6156) );
  HS65_LH_BFX4 U6957 ( .A(n6158), .Z(n6157) );
  HS65_LH_BFX4 U6958 ( .A(n6159), .Z(n6158) );
  HS65_LH_BFX4 U6959 ( .A(n6160), .Z(n6159) );
  HS65_LH_BFX4 U6960 ( .A(n6161), .Z(n6160) );
  HS65_LH_BFX4 U6961 ( .A(n6162), .Z(n6161) );
  HS65_LH_BFX4 U6962 ( .A(n6163), .Z(n6162) );
  HS65_LH_BFX4 U6963 ( .A(n6164), .Z(n6163) );
  HS65_LH_BFX4 U6964 ( .A(n14234), .Z(n6164) );
  HS65_LH_BFX4 U6965 ( .A(n6166), .Z(n6165) );
  HS65_LH_BFX4 U6966 ( .A(n6168), .Z(n6166) );
  HS65_LH_BFX4 U6967 ( .A(\u_DataPath/dataOut_exe_i [14]), .Z(n6167) );
  HS65_LH_BFX4 U6968 ( .A(n15698), .Z(n6168) );
  HS65_LH_BFX4 U6969 ( .A(n6167), .Z(n6169) );
  HS65_LH_BFX4 U6970 ( .A(n6171), .Z(n6170) );
  HS65_LH_BFX4 U6971 ( .A(n6172), .Z(n6171) );
  HS65_LH_BFX4 U6972 ( .A(n6174), .Z(n6172) );
  HS65_LH_BFX4 U6973 ( .A(n6169), .Z(n6173) );
  HS65_LH_BFX4 U6974 ( .A(n6175), .Z(n6174) );
  HS65_LH_BFX4 U6975 ( .A(n6176), .Z(n6175) );
  HS65_LH_BFX4 U6976 ( .A(n6177), .Z(n6176) );
  HS65_LH_BFX4 U6977 ( .A(n6178), .Z(n6177) );
  HS65_LH_BFX4 U6978 ( .A(n6179), .Z(n6178) );
  HS65_LH_BFX4 U6979 ( .A(n6180), .Z(n6179) );
  HS65_LH_BFX4 U6980 ( .A(n6181), .Z(n6180) );
  HS65_LH_BFX4 U6981 ( .A(n6182), .Z(n6181) );
  HS65_LH_BFX4 U6982 ( .A(n6183), .Z(n6182) );
  HS65_LH_BFX4 U6983 ( .A(n6184), .Z(n6183) );
  HS65_LH_BFX4 U6984 ( .A(n6185), .Z(n6184) );
  HS65_LH_BFX4 U6985 ( .A(n6186), .Z(n6185) );
  HS65_LH_BFX4 U6986 ( .A(n6219), .Z(n6186) );
  HS65_LH_BFX4 U6989 ( .A(\u_DataPath/pc_4_to_ex_i [14]), .Z(n6189) );
  HS65_LH_BFX4 U7017 ( .A(n6220), .Z(n6217) );
  HS65_LH_BFX4 U7019 ( .A(n6222), .Z(n6219) );
  HS65_LH_BFX4 U7020 ( .A(n6223), .Z(n6220) );
  HS65_LH_BFX4 U7021 ( .A(n6224), .Z(n6221) );
  HS65_LH_BFX4 U7022 ( .A(n6173), .Z(n6222) );
  HS65_LH_BFX4 U7023 ( .A(n6225), .Z(n6223) );
  HS65_LH_BFX4 U7024 ( .A(\u_DataPath/data_read_ex_1_i [14]), .Z(n6224) );
  HS65_LH_BFX4 U7025 ( .A(n6227), .Z(n6225) );
  HS65_LH_BFX4 U7027 ( .A(n6228), .Z(n6227) );
  HS65_LH_BFX4 U7028 ( .A(n6229), .Z(n6228) );
  HS65_LH_BFX4 U7029 ( .A(n14307), .Z(n6229) );
  HS65_LH_BFX4 U7030 ( .A(n6231), .Z(n6230) );
  HS65_LH_BFX4 U7031 ( .A(n6232), .Z(n6231) );
  HS65_LH_BFX4 U7032 ( .A(n6233), .Z(n6232) );
  HS65_LH_BFX4 U7033 ( .A(n6234), .Z(n6233) );
  HS65_LH_BFX4 U7034 ( .A(n6235), .Z(n6234) );
  HS65_LH_BFX4 U7035 ( .A(n6236), .Z(n6235) );
  HS65_LH_BFX4 U7036 ( .A(n6237), .Z(n6236) );
  HS65_LH_BFX4 U7037 ( .A(n6238), .Z(n6237) );
  HS65_LH_BFX4 U7038 ( .A(n6239), .Z(n6238) );
  HS65_LH_BFX4 U7039 ( .A(n6240), .Z(n6239) );
  HS65_LH_BFX4 U7040 ( .A(n6241), .Z(n6240) );
  HS65_LH_BFX4 U7041 ( .A(n6242), .Z(n6241) );
  HS65_LH_BFX4 U7042 ( .A(n6243), .Z(n6242) );
  HS65_LH_BFX4 U7043 ( .A(n6244), .Z(n6243) );
  HS65_LH_BFX4 U7044 ( .A(n6245), .Z(n6244) );
  HS65_LH_BFX4 U7045 ( .A(n6246), .Z(n6245) );
  HS65_LH_BFX4 U7046 ( .A(n6247), .Z(n6246) );
  HS65_LH_BFX4 U7047 ( .A(n6248), .Z(n6247) );
  HS65_LH_BFX4 U7048 ( .A(n6249), .Z(n6248) );
  HS65_LH_BFX4 U7049 ( .A(n14235), .Z(n6249) );
  HS65_LH_BFX4 U7050 ( .A(n6251), .Z(n6250) );
  HS65_LH_BFX4 U7051 ( .A(n6252), .Z(n6251) );
  HS65_LH_BFX4 U7052 ( .A(n6253), .Z(n6252) );
  HS65_LH_BFX4 U7053 ( .A(n6254), .Z(n6253) );
  HS65_LH_BFX4 U7054 ( .A(n6255), .Z(n6254) );
  HS65_LH_BFX4 U7055 ( .A(n6256), .Z(n6255) );
  HS65_LH_BFX4 U7056 ( .A(n6257), .Z(n6256) );
  HS65_LH_BFX4 U7057 ( .A(n6258), .Z(n6257) );
  HS65_LH_BFX4 U7058 ( .A(n6259), .Z(n6258) );
  HS65_LH_BFX4 U7059 ( .A(n6260), .Z(n6259) );
  HS65_LH_BFX4 U7060 ( .A(n6261), .Z(n6260) );
  HS65_LH_BFX4 U7061 ( .A(n6262), .Z(n6261) );
  HS65_LH_BFX4 U7062 ( .A(n6263), .Z(n6262) );
  HS65_LH_BFX4 U7063 ( .A(n6264), .Z(n6263) );
  HS65_LH_BFX4 U7064 ( .A(n6265), .Z(n6264) );
  HS65_LH_BFX4 U7065 ( .A(n6266), .Z(n6265) );
  HS65_LH_BFX4 U7066 ( .A(n6267), .Z(n6266) );
  HS65_LH_BFX4 U7067 ( .A(n6268), .Z(n6267) );
  HS65_LH_BFX4 U7068 ( .A(n6269), .Z(n6268) );
  HS65_LH_BFX4 U7069 ( .A(n6270), .Z(n6269) );
  HS65_LH_BFX4 U7070 ( .A(n6271), .Z(n6270) );
  HS65_LH_BFX4 U7071 ( .A(n6272), .Z(n6271) );
  HS65_LH_BFX4 U7072 ( .A(n6273), .Z(n6272) );
  HS65_LH_BFX4 U7073 ( .A(n6274), .Z(n6273) );
  HS65_LH_BFX4 U7074 ( .A(n14328), .Z(n6274) );
  HS65_LH_BFX4 U7105 ( .A(n6307), .Z(n6305) );
  HS65_LH_BFX4 U7107 ( .A(n6309), .Z(n6307) );
  HS65_LH_BFX4 U7109 ( .A(n6312), .Z(n6309) );
  HS65_LH_BFX4 U7111 ( .A(n14298), .Z(n6311) );
  HS65_LH_BFX4 U7112 ( .A(n6313), .Z(n6312) );
  HS65_LH_BFX4 U7113 ( .A(n14330), .Z(n6313) );
  HS65_LH_BFX4 U7114 ( .A(n6315), .Z(n6314) );
  HS65_LH_BFX4 U7115 ( .A(n6316), .Z(n6315) );
  HS65_LH_BFX4 U7116 ( .A(n6317), .Z(n6316) );
  HS65_LH_BFX4 U7117 ( .A(n6318), .Z(n6317) );
  HS65_LH_BFX4 U7118 ( .A(n6319), .Z(n6318) );
  HS65_LH_BFX4 U7119 ( .A(n6320), .Z(n6319) );
  HS65_LH_BFX4 U7120 ( .A(n6321), .Z(n6320) );
  HS65_LH_BFX4 U7121 ( .A(n6322), .Z(n6321) );
  HS65_LH_BFX4 U7122 ( .A(n6323), .Z(n6322) );
  HS65_LH_BFX4 U7123 ( .A(n6324), .Z(n6323) );
  HS65_LH_BFX4 U7124 ( .A(n6325), .Z(n6324) );
  HS65_LH_BFX4 U7125 ( .A(n6326), .Z(n6325) );
  HS65_LH_BFX4 U7126 ( .A(n6327), .Z(n6326) );
  HS65_LH_BFX4 U7127 ( .A(n6328), .Z(n6327) );
  HS65_LH_BFX4 U7128 ( .A(n6329), .Z(n6328) );
  HS65_LH_BFX4 U7129 ( .A(n6330), .Z(n6329) );
  HS65_LH_BFX4 U7130 ( .A(n6331), .Z(n6330) );
  HS65_LH_BFX4 U7131 ( .A(n6332), .Z(n6331) );
  HS65_LH_BFX4 U7132 ( .A(n6333), .Z(n6332) );
  HS65_LH_BFX4 U7133 ( .A(n14205), .Z(n6333) );
  HS65_LH_BFX4 U7134 ( .A(n6335), .Z(n6334) );
  HS65_LH_BFX4 U7135 ( .A(n6336), .Z(n6335) );
  HS65_LH_BFX4 U7136 ( .A(n6337), .Z(n6336) );
  HS65_LH_BFX4 U7137 ( .A(n6338), .Z(n6337) );
  HS65_LH_BFX4 U7138 ( .A(n6339), .Z(n6338) );
  HS65_LH_BFX4 U7139 ( .A(n6340), .Z(n6339) );
  HS65_LH_BFX4 U7140 ( .A(n6341), .Z(n6340) );
  HS65_LH_BFX4 U7141 ( .A(n6342), .Z(n6341) );
  HS65_LH_BFX4 U7142 ( .A(n6343), .Z(n6342) );
  HS65_LH_BFX4 U7143 ( .A(n6344), .Z(n6343) );
  HS65_LH_BFX4 U7144 ( .A(n6345), .Z(n6344) );
  HS65_LH_BFX4 U7145 ( .A(n6346), .Z(n6345) );
  HS65_LH_BFX4 U7146 ( .A(n6347), .Z(n6346) );
  HS65_LH_BFX4 U7147 ( .A(n6348), .Z(n6347) );
  HS65_LH_BFX4 U7148 ( .A(n6349), .Z(n6348) );
  HS65_LH_BFX4 U7149 ( .A(n6350), .Z(n6349) );
  HS65_LH_BFX4 U7150 ( .A(n6351), .Z(n6350) );
  HS65_LH_BFX4 U7151 ( .A(n6352), .Z(n6351) );
  HS65_LH_BFX4 U7152 ( .A(n6353), .Z(n6352) );
  HS65_LH_BFX4 U7153 ( .A(n6354), .Z(n6353) );
  HS65_LH_BFX4 U7154 ( .A(n6355), .Z(n6354) );
  HS65_LH_BFX4 U7155 ( .A(n6356), .Z(n6355) );
  HS65_LH_BFX4 U7156 ( .A(n6357), .Z(n6356) );
  HS65_LH_BFX4 U7157 ( .A(n6358), .Z(n6357) );
  HS65_LH_BFX4 U7158 ( .A(n15654), .Z(n6358) );
  HS65_LH_BFX4 U7169 ( .A(n6371), .Z(n6369) );
  HS65_LH_BFX4 U7171 ( .A(n6373), .Z(n6371) );
  HS65_LH_BFX4 U7173 ( .A(n6375), .Z(n6373) );
  HS65_LH_BFX4 U7175 ( .A(n6377), .Z(n6375) );
  HS65_LH_BFX4 U7177 ( .A(n6379), .Z(n6377) );
  HS65_LH_BFX4 U7179 ( .A(n6382), .Z(n6379) );
  HS65_LH_BFX4 U7182 ( .A(n6384), .Z(n6382) );
  HS65_LH_BFX4 U7184 ( .A(n6386), .Z(n6384) );
  HS65_LH_BFX4 U7186 ( .A(n6388), .Z(n6386) );
  HS65_LH_BFX4 U7188 ( .A(n6390), .Z(n6388) );
  HS65_LH_BFX4 U7190 ( .A(n6393), .Z(n6390) );
  HS65_LH_BFX4 U7193 ( .A(n6395), .Z(n6393) );
  HS65_LH_BFX4 U7195 ( .A(n6396), .Z(n6395) );
  HS65_LH_BFX4 U7196 ( .A(n6397), .Z(n6396) );
  HS65_LH_BFX4 U7197 ( .A(n6398), .Z(n6397) );
  HS65_LH_BFX4 U7198 ( .A(n14357), .Z(n6398) );
  HS65_LH_BFX4 U7199 ( .A(n6400), .Z(n6399) );
  HS65_LH_BFX4 U7200 ( .A(n6401), .Z(n6400) );
  HS65_LH_BFX4 U7201 ( .A(n6402), .Z(n6401) );
  HS65_LH_BFX4 U7202 ( .A(n6403), .Z(n6402) );
  HS65_LH_BFX4 U7203 ( .A(n6404), .Z(n6403) );
  HS65_LH_BFX4 U7204 ( .A(n6405), .Z(n6404) );
  HS65_LH_BFX4 U7205 ( .A(n6406), .Z(n6405) );
  HS65_LH_BFX4 U7206 ( .A(n6407), .Z(n6406) );
  HS65_LH_BFX4 U7207 ( .A(n6408), .Z(n6407) );
  HS65_LH_BFX4 U7208 ( .A(n6409), .Z(n6408) );
  HS65_LH_BFX4 U7209 ( .A(n6410), .Z(n6409) );
  HS65_LH_BFX4 U7210 ( .A(n6411), .Z(n6410) );
  HS65_LH_BFX4 U7211 ( .A(n6412), .Z(n6411) );
  HS65_LH_BFX4 U7212 ( .A(n6413), .Z(n6412) );
  HS65_LH_BFX4 U7213 ( .A(n6414), .Z(n6413) );
  HS65_LH_BFX4 U7214 ( .A(n6415), .Z(n6414) );
  HS65_LH_BFX4 U7215 ( .A(n6416), .Z(n6415) );
  HS65_LH_BFX4 U7216 ( .A(n6417), .Z(n6416) );
  HS65_LH_BFX4 U7217 ( .A(n6418), .Z(n6417) );
  HS65_LH_BFX4 U7218 ( .A(n14202), .Z(n6418) );
  HS65_LH_BFX4 U7230 ( .A(n6431), .Z(n6430) );
  HS65_LH_BFX4 U7231 ( .A(n6432), .Z(n6431) );
  HS65_LH_BFX4 U7232 ( .A(n6433), .Z(n6432) );
  HS65_LH_BFX4 U7233 ( .A(n6434), .Z(n6433) );
  HS65_LH_BFX4 U7234 ( .A(n6435), .Z(n6434) );
  HS65_LH_BFX4 U7235 ( .A(n6436), .Z(n6435) );
  HS65_LH_BFX4 U7236 ( .A(n6437), .Z(n6436) );
  HS65_LH_BFX4 U7237 ( .A(n6438), .Z(n6437) );
  HS65_LH_BFX4 U7238 ( .A(n6439), .Z(n6438) );
  HS65_LH_BFX4 U7239 ( .A(n6440), .Z(n6439) );
  HS65_LH_BFX4 U7240 ( .A(n6441), .Z(n6440) );
  HS65_LH_BFX4 U7241 ( .A(n6442), .Z(n6441) );
  HS65_LH_BFX4 U7242 ( .A(n6443), .Z(n6442) );
  HS65_LH_BFX4 U7243 ( .A(n14379), .Z(n6443) );
  HS65_LH_BFX4 U7246 ( .A(n6449), .Z(n6446) );
  HS65_LH_BFX4 U7249 ( .A(n6452), .Z(n6449) );
  HS65_LH_BFX4 U7252 ( .A(n6455), .Z(n6452) );
  HS65_LH_BFX4 U7255 ( .A(n6458), .Z(n6455) );
  HS65_LH_BFX4 U7258 ( .A(n6461), .Z(n6458) );
  HS65_LH_BFX4 U7261 ( .A(n6464), .Z(n6461) );
  HS65_LH_BFX4 U7264 ( .A(n6467), .Z(n6464) );
  HS65_LH_BFX4 U7267 ( .A(n6470), .Z(n6467) );
  HS65_LH_BFX4 U7270 ( .A(n6473), .Z(n6470) );
  HS65_LH_BFX4 U7273 ( .A(n6476), .Z(n6473) );
  HS65_LH_BFX4 U7276 ( .A(n6479), .Z(n6476) );
  HS65_LH_BFX4 U7279 ( .A(n6482), .Z(n6479) );
  HS65_LH_BFX4 U7282 ( .A(n6485), .Z(n6482) );
  HS65_LH_BFX4 U7285 ( .A(n6488), .Z(n6485) );
  HS65_LH_BFX4 U7288 ( .A(n6491), .Z(n6488) );
  HS65_LH_BFX4 U7291 ( .A(n6496), .Z(n6491) );
  HS65_LH_BFX4 U7296 ( .A(n6498), .Z(n6496) );
  HS65_LH_BFX4 U7298 ( .A(n6500), .Z(n6498) );
  HS65_LH_BFX4 U7300 ( .A(n6502), .Z(n6500) );
  HS65_LH_BFX4 U7302 ( .A(n6504), .Z(n6502) );
  HS65_LH_BFX4 U7304 ( .A(n6505), .Z(n6504) );
  HS65_LH_BFX4 U7305 ( .A(n6506), .Z(n6505) );
  HS65_LH_BFX4 U7306 ( .A(n6507), .Z(n6506) );
  HS65_LH_BFX4 U7307 ( .A(\u_DataPath/u_idexreg/N28 ), .Z(n6507) );
  HS65_LH_BFX4 U7343 ( .A(n6545), .Z(n6543) );
  HS65_LH_BFX4 U7345 ( .A(n6547), .Z(n6545) );
  HS65_LH_BFX4 U7347 ( .A(n6549), .Z(n6547) );
  HS65_LH_BFX4 U7349 ( .A(n6551), .Z(n6549) );
  HS65_LH_BFX4 U7351 ( .A(n6553), .Z(n6551) );
  HS65_LH_BFX4 U7353 ( .A(n6555), .Z(n6553) );
  HS65_LH_BFX4 U7355 ( .A(n6557), .Z(n6555) );
  HS65_LH_BFX4 U7357 ( .A(n6559), .Z(n6557) );
  HS65_LH_BFX4 U7359 ( .A(n6561), .Z(n6559) );
  HS65_LH_BFX4 U7361 ( .A(n6563), .Z(n6561) );
  HS65_LH_BFX4 U7363 ( .A(n6565), .Z(n6563) );
  HS65_LH_BFX4 U7365 ( .A(n6567), .Z(n6565) );
  HS65_LH_BFX4 U7367 ( .A(n6568), .Z(n6567) );
  HS65_LH_BFX4 U7368 ( .A(n6569), .Z(n6568) );
  HS65_LH_BFX4 U7369 ( .A(n6570), .Z(n6569) );
  HS65_LH_BFX4 U7370 ( .A(n6571), .Z(n6570) );
  HS65_LH_BFX4 U7371 ( .A(n14404), .Z(n6571) );
  HS65_LH_BFX4 U7372 ( .A(n6573), .Z(n6572) );
  HS65_LH_BFX4 U7373 ( .A(n6574), .Z(n6573) );
  HS65_LH_BFX4 U7374 ( .A(n6575), .Z(n6574) );
  HS65_LH_BFX4 U7375 ( .A(n6576), .Z(n6575) );
  HS65_LH_BFX4 U7376 ( .A(n6577), .Z(n6576) );
  HS65_LH_BFX4 U7377 ( .A(n6578), .Z(n6577) );
  HS65_LH_BFX4 U7378 ( .A(n6579), .Z(n6578) );
  HS65_LH_BFX4 U7379 ( .A(n6580), .Z(n6579) );
  HS65_LH_BFX4 U7380 ( .A(n6581), .Z(n6580) );
  HS65_LH_BFX4 U7381 ( .A(n6582), .Z(n6581) );
  HS65_LH_BFX4 U7382 ( .A(n6583), .Z(n6582) );
  HS65_LH_BFX4 U7383 ( .A(n6584), .Z(n6583) );
  HS65_LH_BFX4 U7384 ( .A(n6585), .Z(n6584) );
  HS65_LH_BFX4 U7385 ( .A(n6586), .Z(n6585) );
  HS65_LH_BFX4 U7386 ( .A(n6587), .Z(n6586) );
  HS65_LH_BFX4 U7387 ( .A(n6588), .Z(n6587) );
  HS65_LH_BFX4 U7388 ( .A(n6589), .Z(n6588) );
  HS65_LH_BFX4 U7389 ( .A(n6590), .Z(n6589) );
  HS65_LH_BFX4 U7390 ( .A(n6591), .Z(n6590) );
  HS65_LH_BFX4 U7391 ( .A(n14219), .Z(n6591) );
  HS65_LH_BFX4 U7392 ( .A(n6593), .Z(n6592) );
  HS65_LH_BFX4 U7393 ( .A(n6594), .Z(n6593) );
  HS65_LH_BFX4 U7394 ( .A(n6595), .Z(n6594) );
  HS65_LH_BFX4 U7395 ( .A(n6596), .Z(n6595) );
  HS65_LH_BFX4 U7396 ( .A(n6597), .Z(n6596) );
  HS65_LH_BFX4 U7397 ( .A(n6598), .Z(n6597) );
  HS65_LH_BFX4 U7398 ( .A(n6599), .Z(n6598) );
  HS65_LH_BFX4 U7399 ( .A(n6600), .Z(n6599) );
  HS65_LH_BFX4 U7400 ( .A(n6601), .Z(n6600) );
  HS65_LH_BFX4 U7401 ( .A(n6602), .Z(n6601) );
  HS65_LH_BFX4 U7402 ( .A(n6603), .Z(n6602) );
  HS65_LH_BFX4 U7403 ( .A(n6604), .Z(n6603) );
  HS65_LH_BFX4 U7404 ( .A(n6605), .Z(n6604) );
  HS65_LH_BFX4 U7405 ( .A(n6606), .Z(n6605) );
  HS65_LH_BFX4 U7406 ( .A(n6607), .Z(n6606) );
  HS65_LH_BFX4 U7407 ( .A(n6608), .Z(n6607) );
  HS65_LH_BFX4 U7408 ( .A(n6609), .Z(n6608) );
  HS65_LH_BFX4 U7409 ( .A(n6610), .Z(n6609) );
  HS65_LH_BFX4 U7410 ( .A(n6611), .Z(n6610) );
  HS65_LH_BFX4 U7411 ( .A(n6612), .Z(n6611) );
  HS65_LH_BFX4 U7412 ( .A(n6613), .Z(n6612) );
  HS65_LH_BFX4 U7413 ( .A(n6614), .Z(n6613) );
  HS65_LH_BFX4 U7414 ( .A(n6615), .Z(n6614) );
  HS65_LH_BFX4 U7415 ( .A(n6616), .Z(n6615) );
  HS65_LH_BFX4 U7416 ( .A(n14405), .Z(n6616) );
  HS65_LH_BFX4 U7418 ( .A(n6620), .Z(n6618) );
  HS65_LH_BFX4 U7420 ( .A(n6622), .Z(n6620) );
  HS65_LH_BFX4 U7422 ( .A(n6624), .Z(n6622) );
  HS65_LH_BFX4 U7424 ( .A(n6626), .Z(n6624) );
  HS65_LH_BFX4 U7426 ( .A(n6628), .Z(n6626) );
  HS65_LH_BFX4 U7428 ( .A(n6630), .Z(n6628) );
  HS65_LH_BFX4 U7430 ( .A(n6632), .Z(n6630) );
  HS65_LH_BFX4 U7432 ( .A(n6634), .Z(n6632) );
  HS65_LH_BFX4 U7434 ( .A(n6637), .Z(n6634) );
  HS65_LH_BFX4 U7437 ( .A(n6639), .Z(n6637) );
  HS65_LH_BFX4 U7439 ( .A(n6641), .Z(n6639) );
  HS65_LH_BFX4 U7441 ( .A(n6643), .Z(n6641) );
  HS65_LH_BFX4 U7443 ( .A(n6645), .Z(n6643) );
  HS65_LH_BFX4 U7445 ( .A(n6647), .Z(n6645) );
  HS65_LH_BFX4 U7447 ( .A(n6652), .Z(n6647) );
  HS65_LH_CNIVX3 U7449 ( .A(\u_DataPath/pc_4_to_ex_i [3]), .Z(n6649) );
  HS65_LH_CNIVX3 U7450 ( .A(n6649), .Z(n6650) );
  HS65_LH_BFX2 U7451 ( .A(n14925), .Z(n6651) );
  HS65_LH_BFX4 U7452 ( .A(n6653), .Z(n6652) );
  HS65_LH_BFX4 U7453 ( .A(n6654), .Z(n6653) );
  HS65_LH_BFX4 U7454 ( .A(n6655), .Z(n6654) );
  HS65_LH_BFX4 U7455 ( .A(n6656), .Z(n6655) );
  HS65_LH_BFX4 U7456 ( .A(n14429), .Z(n6656) );
  HS65_LH_BFX4 U7457 ( .A(n6658), .Z(n6657) );
  HS65_LH_BFX4 U7458 ( .A(n6659), .Z(n6658) );
  HS65_LH_BFX4 U7459 ( .A(n6660), .Z(n6659) );
  HS65_LH_BFX4 U7460 ( .A(n6661), .Z(n6660) );
  HS65_LH_BFX4 U7461 ( .A(n6662), .Z(n6661) );
  HS65_LH_BFX4 U7462 ( .A(n6663), .Z(n6662) );
  HS65_LH_BFX4 U7463 ( .A(n6664), .Z(n6663) );
  HS65_LH_BFX4 U7464 ( .A(n6665), .Z(n6664) );
  HS65_LH_BFX4 U7465 ( .A(n6666), .Z(n6665) );
  HS65_LH_BFX4 U7466 ( .A(n6667), .Z(n6666) );
  HS65_LH_BFX4 U7467 ( .A(n6668), .Z(n6667) );
  HS65_LH_BFX4 U7468 ( .A(n6669), .Z(n6668) );
  HS65_LH_BFX4 U7469 ( .A(n6670), .Z(n6669) );
  HS65_LH_BFX4 U7470 ( .A(n6671), .Z(n6670) );
  HS65_LH_BFX4 U7471 ( .A(n6672), .Z(n6671) );
  HS65_LH_BFX4 U7472 ( .A(n6673), .Z(n6672) );
  HS65_LH_BFX4 U7473 ( .A(n6674), .Z(n6673) );
  HS65_LH_BFX4 U7474 ( .A(n6675), .Z(n6674) );
  HS65_LH_BFX4 U7475 ( .A(n6676), .Z(n6675) );
  HS65_LH_BFX4 U7476 ( .A(n14199), .Z(n6676) );
  HS65_LH_BFX4 U7477 ( .A(n6678), .Z(n6677) );
  HS65_LH_BFX4 U7478 ( .A(n6679), .Z(n6678) );
  HS65_LH_BFX4 U7479 ( .A(n6680), .Z(n6679) );
  HS65_LH_BFX4 U7480 ( .A(n6681), .Z(n6680) );
  HS65_LH_BFX4 U7481 ( .A(n6682), .Z(n6681) );
  HS65_LH_BFX4 U7482 ( .A(n6683), .Z(n6682) );
  HS65_LH_BFX4 U7483 ( .A(n6684), .Z(n6683) );
  HS65_LH_BFX4 U7484 ( .A(n6685), .Z(n6684) );
  HS65_LH_BFX4 U7485 ( .A(n6686), .Z(n6685) );
  HS65_LH_BFX4 U7486 ( .A(n6687), .Z(n6686) );
  HS65_LH_BFX4 U7487 ( .A(n6688), .Z(n6687) );
  HS65_LH_BFX4 U7488 ( .A(n6689), .Z(n6688) );
  HS65_LH_BFX4 U7489 ( .A(n6690), .Z(n6689) );
  HS65_LH_BFX4 U7490 ( .A(n6691), .Z(n6690) );
  HS65_LH_BFX4 U7491 ( .A(n6692), .Z(n6691) );
  HS65_LH_BFX4 U7492 ( .A(n6693), .Z(n6692) );
  HS65_LH_BFX4 U7493 ( .A(n6694), .Z(n6693) );
  HS65_LH_BFX4 U7494 ( .A(n6695), .Z(n6694) );
  HS65_LH_BFX4 U7495 ( .A(n6696), .Z(n6695) );
  HS65_LH_BFX4 U7496 ( .A(n6697), .Z(n6696) );
  HS65_LH_BFX4 U7497 ( .A(n6698), .Z(n6697) );
  HS65_LH_BFX4 U7498 ( .A(n6699), .Z(n6698) );
  HS65_LH_BFX4 U7499 ( .A(n6700), .Z(n6699) );
  HS65_LH_BFX4 U7500 ( .A(n6701), .Z(n6700) );
  HS65_LH_BFX4 U7501 ( .A(n15662), .Z(n6701) );
  HS65_LH_CNIVX3 U7502 ( .A(\u_DataPath/pc_4_to_ex_i [10]), .Z(n6702) );
  HS65_LH_CNIVX3 U7503 ( .A(n6702), .Z(n6703) );
  HS65_LH_BFX4 U7508 ( .A(n6710), .Z(n6708) );
  HS65_LH_BFX4 U7510 ( .A(n6712), .Z(n6710) );
  HS65_LH_BFX4 U7512 ( .A(n6714), .Z(n6712) );
  HS65_LH_BFX4 U7514 ( .A(n6716), .Z(n6714) );
  HS65_LH_BFX4 U7516 ( .A(n6718), .Z(n6716) );
  HS65_LH_BFX4 U7518 ( .A(n6720), .Z(n6718) );
  HS65_LH_BFX4 U7520 ( .A(n6722), .Z(n6720) );
  HS65_LH_BFX4 U7522 ( .A(n6724), .Z(n6722) );
  HS65_LH_BFX4 U7524 ( .A(n6726), .Z(n6724) );
  HS65_LH_BFX4 U7526 ( .A(n6728), .Z(n6726) );
  HS65_LH_BFX4 U7528 ( .A(n6730), .Z(n6728) );
  HS65_LH_BFX4 U7530 ( .A(n6732), .Z(n6730) );
  HS65_LH_BFX4 U7532 ( .A(n6734), .Z(n6732) );
  HS65_LH_BFX4 U7534 ( .A(n6736), .Z(n6734) );
  HS65_LH_BFX4 U7536 ( .A(n6738), .Z(n6736) );
  HS65_LH_BFX4 U7538 ( .A(n6739), .Z(n6738) );
  HS65_LH_BFX4 U7539 ( .A(n6740), .Z(n6739) );
  HS65_LH_BFX4 U7540 ( .A(n6741), .Z(n6740) );
  HS65_LH_BFX4 U7541 ( .A(n14451), .Z(n6741) );
  HS65_LH_BFX4 U7542 ( .A(n6743), .Z(n6742) );
  HS65_LH_BFX4 U7543 ( .A(n6744), .Z(n6743) );
  HS65_LH_BFX4 U7544 ( .A(n6745), .Z(n6744) );
  HS65_LH_BFX4 U7545 ( .A(n6746), .Z(n6745) );
  HS65_LH_BFX4 U7546 ( .A(n6747), .Z(n6746) );
  HS65_LH_BFX4 U7547 ( .A(n6748), .Z(n6747) );
  HS65_LH_BFX4 U7548 ( .A(n6749), .Z(n6748) );
  HS65_LH_BFX4 U7549 ( .A(n6750), .Z(n6749) );
  HS65_LH_BFX4 U7550 ( .A(n6751), .Z(n6750) );
  HS65_LH_BFX4 U7551 ( .A(n6752), .Z(n6751) );
  HS65_LH_BFX4 U7552 ( .A(n6753), .Z(n6752) );
  HS65_LH_BFX4 U7553 ( .A(n6754), .Z(n6753) );
  HS65_LH_BFX4 U7554 ( .A(n6755), .Z(n6754) );
  HS65_LH_BFX4 U7555 ( .A(n6756), .Z(n6755) );
  HS65_LH_BFX4 U7556 ( .A(n6757), .Z(n6756) );
  HS65_LH_BFX4 U7557 ( .A(n6758), .Z(n6757) );
  HS65_LH_BFX4 U7558 ( .A(n6759), .Z(n6758) );
  HS65_LH_BFX4 U7559 ( .A(n6760), .Z(n6759) );
  HS65_LH_BFX4 U7560 ( .A(n6761), .Z(n6760) );
  HS65_LH_BFX4 U7561 ( .A(n14196), .Z(n6761) );
  HS65_LH_CNIVX3 U7587 ( .A(\u_DataPath/pc_4_to_ex_i [26]), .Z(n6787) );
  HS65_LH_CNIVX3 U7588 ( .A(n6787), .Z(n6788) );
  HS65_LH_BFX4 U7589 ( .A(n6791), .Z(n6789) );
  HS65_LH_BFX4 U7591 ( .A(n6794), .Z(n6791) );
  HS65_LH_BFX4 U7594 ( .A(n6797), .Z(n6794) );
  HS65_LH_BFX4 U7597 ( .A(n6800), .Z(n6797) );
  HS65_LH_BFX4 U7600 ( .A(n6803), .Z(n6800) );
  HS65_LH_BFX4 U7603 ( .A(n6806), .Z(n6803) );
  HS65_LH_BFX4 U7606 ( .A(n6809), .Z(n6806) );
  HS65_LH_BFX4 U7609 ( .A(n6812), .Z(n6809) );
  HS65_LH_BFX4 U7612 ( .A(n6815), .Z(n6812) );
  HS65_LH_BFX4 U7615 ( .A(n6818), .Z(n6815) );
  HS65_LH_BFX4 U7618 ( .A(n6821), .Z(n6818) );
  HS65_LH_BFX4 U7621 ( .A(n6824), .Z(n6821) );
  HS65_LH_BFX4 U7624 ( .A(n6827), .Z(n6824) );
  HS65_LH_BFX4 U7627 ( .A(n6830), .Z(n6827) );
  HS65_LH_BFX4 U7630 ( .A(n6833), .Z(n6830) );
  HS65_LH_BFX4 U7633 ( .A(n6836), .Z(n6833) );
  HS65_LH_BFX4 U7636 ( .A(n6839), .Z(n6836) );
  HS65_LH_BFX4 U7639 ( .A(n6842), .Z(n6839) );
  HS65_LH_BFX4 U7642 ( .A(n6845), .Z(n6842) );
  HS65_LH_BFX4 U7645 ( .A(n6847), .Z(n6845) );
  HS65_LH_BFX4 U7647 ( .A(n6849), .Z(n6847) );
  HS65_LH_BFX4 U7649 ( .A(n6850), .Z(n6849) );
  HS65_LH_BFX4 U7650 ( .A(n6851), .Z(n6850) );
  HS65_LH_BFX4 U7651 ( .A(n6852), .Z(n6851) );
  HS65_LH_BFX4 U7652 ( .A(\u_DataPath/u_idexreg/N35 ), .Z(n6852) );
  HS65_LH_BFX4 U7653 ( .A(n6854), .Z(n6853) );
  HS65_LH_BFX4 U7654 ( .A(n6855), .Z(n6854) );
  HS65_LH_BFX4 U7655 ( .A(n6856), .Z(n6855) );
  HS65_LH_BFX4 U7656 ( .A(n6857), .Z(n6856) );
  HS65_LH_BFX4 U7657 ( .A(n6858), .Z(n6857) );
  HS65_LH_BFX4 U7658 ( .A(n6859), .Z(n6858) );
  HS65_LH_BFX4 U7659 ( .A(n6860), .Z(n6859) );
  HS65_LH_BFX4 U7660 ( .A(n6861), .Z(n6860) );
  HS65_LH_BFX4 U7661 ( .A(n6862), .Z(n6861) );
  HS65_LH_BFX4 U7662 ( .A(n6863), .Z(n6862) );
  HS65_LH_BFX4 U7663 ( .A(n6864), .Z(n6863) );
  HS65_LH_BFX4 U7664 ( .A(n6865), .Z(n6864) );
  HS65_LH_BFX4 U7665 ( .A(n6866), .Z(n6865) );
  HS65_LH_BFX4 U7666 ( .A(n6867), .Z(n6866) );
  HS65_LH_BFX4 U7667 ( .A(n6868), .Z(n6867) );
  HS65_LH_BFX4 U7668 ( .A(n6869), .Z(n6868) );
  HS65_LH_BFX4 U7669 ( .A(n6870), .Z(n6869) );
  HS65_LH_BFX4 U7670 ( .A(n6871), .Z(n6870) );
  HS65_LH_BFX4 U7671 ( .A(n6872), .Z(n6871) );
  HS65_LH_BFX4 U7672 ( .A(n14193), .Z(n6872) );
  HS65_LH_BFX4 U7698 ( .A(n6901), .Z(n6898) );
  HS65_LH_BFX4 U7701 ( .A(n6904), .Z(n6901) );
  HS65_LH_BFX4 U7704 ( .A(n6907), .Z(n6904) );
  HS65_LH_BFX4 U7707 ( .A(n6910), .Z(n6907) );
  HS65_LH_BFX4 U7710 ( .A(n6913), .Z(n6910) );
  HS65_LH_BFX4 U7713 ( .A(n6916), .Z(n6913) );
  HS65_LH_BFX4 U7716 ( .A(n6919), .Z(n6916) );
  HS65_LH_BFX4 U7719 ( .A(n6922), .Z(n6919) );
  HS65_LH_BFX4 U7722 ( .A(n6925), .Z(n6922) );
  HS65_LH_BFX4 U7725 ( .A(n6928), .Z(n6925) );
  HS65_LH_BFX4 U7728 ( .A(n6931), .Z(n6928) );
  HS65_LH_BFX4 U7731 ( .A(n6934), .Z(n6931) );
  HS65_LH_BFX4 U7734 ( .A(n6937), .Z(n6934) );
  HS65_LH_BFX4 U7737 ( .A(n6940), .Z(n6937) );
  HS65_LH_BFX4 U7740 ( .A(n6943), .Z(n6940) );
  HS65_LH_BFX4 U7743 ( .A(n6946), .Z(n6943) );
  HS65_LH_BFX4 U7746 ( .A(n6949), .Z(n6946) );
  HS65_LH_BFX4 U7749 ( .A(n6952), .Z(n6949) );
  HS65_LH_BFX4 U7752 ( .A(n6954), .Z(n6952) );
  HS65_LH_BFX4 U7754 ( .A(n6956), .Z(n6954) );
  HS65_LH_BFX4 U7756 ( .A(n6958), .Z(n6956) );
  HS65_LH_BFX4 U7758 ( .A(n6959), .Z(n6958) );
  HS65_LH_BFX4 U7759 ( .A(n6960), .Z(n6959) );
  HS65_LH_BFX4 U7760 ( .A(n6961), .Z(n6960) );
  HS65_LH_BFX4 U7761 ( .A(\u_DataPath/u_idexreg/N32 ), .Z(n6961) );
  HS65_LH_BFX4 U7762 ( .A(n6963), .Z(n6962) );
  HS65_LH_BFX4 U7763 ( .A(n6964), .Z(n6963) );
  HS65_LH_BFX4 U7764 ( .A(n6965), .Z(n6964) );
  HS65_LH_BFX4 U7765 ( .A(n6966), .Z(n6965) );
  HS65_LH_BFX4 U7766 ( .A(n6967), .Z(n6966) );
  HS65_LH_BFX4 U7767 ( .A(n6968), .Z(n6967) );
  HS65_LH_BFX4 U7768 ( .A(n6969), .Z(n6968) );
  HS65_LH_BFX4 U7769 ( .A(n6970), .Z(n6969) );
  HS65_LH_BFX4 U7770 ( .A(n6971), .Z(n6970) );
  HS65_LH_BFX4 U7771 ( .A(n6972), .Z(n6971) );
  HS65_LH_BFX4 U7772 ( .A(n6973), .Z(n6972) );
  HS65_LH_BFX4 U7773 ( .A(n6974), .Z(n6973) );
  HS65_LH_BFX4 U7774 ( .A(n6975), .Z(n6974) );
  HS65_LH_BFX4 U7775 ( .A(n6976), .Z(n6975) );
  HS65_LH_BFX4 U7776 ( .A(n6977), .Z(n6976) );
  HS65_LH_BFX4 U7777 ( .A(n6978), .Z(n6977) );
  HS65_LH_BFX4 U7778 ( .A(n6979), .Z(n6978) );
  HS65_LH_BFX4 U7779 ( .A(n6980), .Z(n6979) );
  HS65_LH_BFX4 U7780 ( .A(n6981), .Z(n6980) );
  HS65_LH_BFX4 U7781 ( .A(n14190), .Z(n6981) );
  HS65_LH_BFX4 U7808 ( .A(n7011), .Z(n7008) );
  HS65_LH_BFX4 U7811 ( .A(n7014), .Z(n7011) );
  HS65_LH_BFX4 U7814 ( .A(n7017), .Z(n7014) );
  HS65_LH_BFX4 U7817 ( .A(n7020), .Z(n7017) );
  HS65_LH_BFX4 U7820 ( .A(n7023), .Z(n7020) );
  HS65_LH_BFX4 U7823 ( .A(n7026), .Z(n7023) );
  HS65_LH_BFX4 U7826 ( .A(n7029), .Z(n7026) );
  HS65_LH_BFX4 U7829 ( .A(n7032), .Z(n7029) );
  HS65_LH_BFX4 U7832 ( .A(n7035), .Z(n7032) );
  HS65_LH_BFX4 U7835 ( .A(n7038), .Z(n7035) );
  HS65_LH_BFX4 U7838 ( .A(n7041), .Z(n7038) );
  HS65_LH_BFX4 U7841 ( .A(n7044), .Z(n7041) );
  HS65_LH_BFX4 U7844 ( .A(n7047), .Z(n7044) );
  HS65_LH_BFX4 U7847 ( .A(n7050), .Z(n7047) );
  HS65_LH_BFX4 U7850 ( .A(n7053), .Z(n7050) );
  HS65_LH_BFX4 U7853 ( .A(n7056), .Z(n7053) );
  HS65_LH_BFX4 U7856 ( .A(n7059), .Z(n7056) );
  HS65_LH_BFX4 U7859 ( .A(n7061), .Z(n7059) );
  HS65_LH_BFX4 U7861 ( .A(n7063), .Z(n7061) );
  HS65_LH_BFX4 U7863 ( .A(n7065), .Z(n7063) );
  HS65_LH_BFX4 U7865 ( .A(n7067), .Z(n7065) );
  HS65_LH_BFX4 U7867 ( .A(n7068), .Z(n7067) );
  HS65_LH_BFX4 U7868 ( .A(n7069), .Z(n7068) );
  HS65_LH_BFX4 U7869 ( .A(n7070), .Z(n7069) );
  HS65_LH_BFX4 U7870 ( .A(\u_DataPath/u_idexreg/N39 ), .Z(n7070) );
  HS65_LH_BFX4 U7871 ( .A(n7072), .Z(n7071) );
  HS65_LH_BFX4 U7872 ( .A(n7073), .Z(n7072) );
  HS65_LH_BFX4 U7873 ( .A(n7074), .Z(n7073) );
  HS65_LH_BFX4 U7874 ( .A(n7075), .Z(n7074) );
  HS65_LH_BFX4 U7875 ( .A(n7076), .Z(n7075) );
  HS65_LH_BFX4 U7876 ( .A(n7077), .Z(n7076) );
  HS65_LH_BFX4 U7877 ( .A(n7078), .Z(n7077) );
  HS65_LH_BFX4 U7878 ( .A(n7079), .Z(n7078) );
  HS65_LH_BFX4 U7879 ( .A(n7080), .Z(n7079) );
  HS65_LH_BFX4 U7880 ( .A(n7081), .Z(n7080) );
  HS65_LH_BFX4 U7881 ( .A(n7082), .Z(n7081) );
  HS65_LH_BFX4 U7882 ( .A(n7083), .Z(n7082) );
  HS65_LH_BFX4 U7883 ( .A(n7084), .Z(n7083) );
  HS65_LH_BFX4 U7884 ( .A(n7085), .Z(n7084) );
  HS65_LH_BFX4 U7885 ( .A(n7086), .Z(n7085) );
  HS65_LH_BFX4 U7886 ( .A(n7087), .Z(n7086) );
  HS65_LH_BFX4 U7887 ( .A(n7088), .Z(n7087) );
  HS65_LH_BFX4 U7888 ( .A(n7089), .Z(n7088) );
  HS65_LH_BFX4 U7889 ( .A(n7090), .Z(n7089) );
  HS65_LH_BFX4 U7890 ( .A(n14187), .Z(n7090) );
  HS65_LH_BFX4 U7891 ( .A(n7092), .Z(n7091) );
  HS65_LH_BFX4 U7892 ( .A(n7093), .Z(n7092) );
  HS65_LH_BFX4 U7893 ( .A(n7094), .Z(n7093) );
  HS65_LH_BFX4 U7894 ( .A(n7095), .Z(n7094) );
  HS65_LH_BFX4 U7895 ( .A(n7096), .Z(n7095) );
  HS65_LH_BFX4 U7896 ( .A(n7097), .Z(n7096) );
  HS65_LH_BFX4 U7897 ( .A(n7098), .Z(n7097) );
  HS65_LH_BFX4 U7898 ( .A(n7099), .Z(n7098) );
  HS65_LH_BFX4 U7899 ( .A(n7100), .Z(n7099) );
  HS65_LH_BFX4 U7900 ( .A(n7101), .Z(n7100) );
  HS65_LH_BFX4 U7901 ( .A(n7102), .Z(n7101) );
  HS65_LH_BFX4 U7902 ( .A(n7103), .Z(n7102) );
  HS65_LH_BFX4 U7903 ( .A(n7104), .Z(n7103) );
  HS65_LH_BFX4 U7904 ( .A(n7105), .Z(n7104) );
  HS65_LH_BFX4 U7905 ( .A(n7106), .Z(n7105) );
  HS65_LH_BFX4 U7906 ( .A(n7107), .Z(n7106) );
  HS65_LH_BFX4 U7907 ( .A(n7108), .Z(n7107) );
  HS65_LH_BFX4 U7908 ( .A(n7109), .Z(n7108) );
  HS65_LH_BFX4 U7909 ( .A(n7110), .Z(n7109) );
  HS65_LH_BFX4 U7910 ( .A(n7111), .Z(n7110) );
  HS65_LH_BFX4 U7911 ( .A(n7112), .Z(n7111) );
  HS65_LH_BFX4 U7912 ( .A(n7113), .Z(n7112) );
  HS65_LH_BFX4 U7913 ( .A(n7114), .Z(n7113) );
  HS65_LH_BFX4 U7914 ( .A(n7115), .Z(n7114) );
  HS65_LH_BFX4 U7915 ( .A(n15660), .Z(n7115) );
  HS65_LH_BFX4 U7932 ( .A(n7134), .Z(n7132) );
  HS65_LH_BFX4 U7934 ( .A(n7136), .Z(n7134) );
  HS65_LH_BFX4 U7936 ( .A(n7138), .Z(n7136) );
  HS65_LH_BFX4 U7938 ( .A(n7140), .Z(n7138) );
  HS65_LH_BFX4 U7940 ( .A(n7142), .Z(n7140) );
  HS65_LH_BFX4 U7942 ( .A(n7144), .Z(n7142) );
  HS65_LH_BFX4 U7944 ( .A(n7146), .Z(n7144) );
  HS65_LH_BFX4 U7946 ( .A(n7148), .Z(n7146) );
  HS65_LH_BFX4 U7948 ( .A(n7150), .Z(n7148) );
  HS65_LH_BFX4 U7950 ( .A(n7151), .Z(n7150) );
  HS65_LH_BFX4 U7951 ( .A(n7152), .Z(n7151) );
  HS65_LH_BFX4 U7952 ( .A(n7153), .Z(n7152) );
  HS65_LH_BFX4 U7953 ( .A(n14543), .Z(n7153) );
  HS65_LH_BFX4 U7954 ( .A(n7155), .Z(n7154) );
  HS65_LH_BFX4 U7955 ( .A(n7156), .Z(n7155) );
  HS65_LH_BFX4 U7956 ( .A(n7157), .Z(n7156) );
  HS65_LH_BFX4 U7957 ( .A(n7158), .Z(n7157) );
  HS65_LH_BFX4 U7958 ( .A(n7159), .Z(n7158) );
  HS65_LH_BFX4 U7959 ( .A(n7160), .Z(n7159) );
  HS65_LH_BFX4 U7960 ( .A(n7161), .Z(n7160) );
  HS65_LH_BFX4 U7961 ( .A(n7162), .Z(n7161) );
  HS65_LH_BFX4 U7962 ( .A(n7163), .Z(n7162) );
  HS65_LH_BFX4 U7963 ( .A(n7164), .Z(n7163) );
  HS65_LH_BFX4 U7964 ( .A(n7165), .Z(n7164) );
  HS65_LH_BFX4 U7965 ( .A(n7166), .Z(n7165) );
  HS65_LH_BFX4 U7966 ( .A(n7167), .Z(n7166) );
  HS65_LH_BFX4 U7967 ( .A(n7168), .Z(n7167) );
  HS65_LH_BFX4 U7968 ( .A(n7169), .Z(n7168) );
  HS65_LH_BFX4 U7969 ( .A(n7170), .Z(n7169) );
  HS65_LH_BFX4 U7970 ( .A(n7171), .Z(n7170) );
  HS65_LH_BFX4 U7971 ( .A(n7172), .Z(n7171) );
  HS65_LH_BFX4 U7972 ( .A(n7173), .Z(n7172) );
  HS65_LH_BFX4 U7973 ( .A(n14184), .Z(n7173) );
  HS65_LH_BFX4 U7974 ( .A(n7175), .Z(n7174) );
  HS65_LH_BFX4 U7975 ( .A(n7176), .Z(n7175) );
  HS65_LH_BFX4 U7976 ( .A(n7177), .Z(n7176) );
  HS65_LH_BFX4 U7977 ( .A(n7178), .Z(n7177) );
  HS65_LH_BFX4 U7978 ( .A(n7179), .Z(n7178) );
  HS65_LH_BFX4 U7979 ( .A(n7180), .Z(n7179) );
  HS65_LH_BFX4 U7980 ( .A(n7181), .Z(n7180) );
  HS65_LH_BFX4 U7981 ( .A(n7182), .Z(n7181) );
  HS65_LH_BFX4 U7982 ( .A(n7183), .Z(n7182) );
  HS65_LH_BFX4 U7983 ( .A(n7184), .Z(n7183) );
  HS65_LH_BFX4 U7984 ( .A(n7185), .Z(n7184) );
  HS65_LH_BFX4 U7985 ( .A(n7186), .Z(n7185) );
  HS65_LH_BFX4 U7986 ( .A(n7187), .Z(n7186) );
  HS65_LH_BFX4 U7987 ( .A(n7188), .Z(n7187) );
  HS65_LH_BFX4 U7988 ( .A(n7189), .Z(n7188) );
  HS65_LH_BFX4 U7989 ( .A(n7190), .Z(n7189) );
  HS65_LH_BFX4 U7990 ( .A(n7191), .Z(n7190) );
  HS65_LH_BFX4 U7991 ( .A(n7192), .Z(n7191) );
  HS65_LH_BFX4 U7992 ( .A(n7193), .Z(n7192) );
  HS65_LH_BFX4 U7993 ( .A(n7194), .Z(n7193) );
  HS65_LH_BFX4 U7994 ( .A(n7195), .Z(n7194) );
  HS65_LH_BFX4 U7995 ( .A(n7196), .Z(n7195) );
  HS65_LH_BFX4 U7996 ( .A(n7197), .Z(n7196) );
  HS65_LH_BFX4 U7997 ( .A(n7198), .Z(n7197) );
  HS65_LH_BFX4 U7998 ( .A(n15648), .Z(n7198) );
  HS65_LH_BFX4 U7999 ( .A(n7201), .Z(n7199) );
  HS65_LH_BFX4 U8001 ( .A(n7203), .Z(n7201) );
  HS65_LH_BFX4 U8003 ( .A(n7205), .Z(n7203) );
  HS65_LH_BFX4 U8005 ( .A(n7207), .Z(n7205) );
  HS65_LH_BFX4 U8007 ( .A(n7209), .Z(n7207) );
  HS65_LH_BFX4 U8009 ( .A(n7211), .Z(n7209) );
  HS65_LH_BFX4 U8011 ( .A(n7213), .Z(n7211) );
  HS65_LH_BFX4 U8013 ( .A(n7215), .Z(n7213) );
  HS65_LH_BFX4 U8015 ( .A(n7217), .Z(n7215) );
  HS65_LH_BFX4 U8017 ( .A(n7219), .Z(n7217) );
  HS65_LH_BFX4 U8019 ( .A(n7221), .Z(n7219) );
  HS65_LH_BFX4 U8021 ( .A(n7223), .Z(n7221) );
  HS65_LH_BFX4 U8023 ( .A(n7225), .Z(n7223) );
  HS65_LH_BFX4 U8025 ( .A(n7227), .Z(n7225) );
  HS65_LH_BFX4 U8027 ( .A(n7229), .Z(n7227) );
  HS65_LH_BFX4 U8029 ( .A(n7231), .Z(n7229) );
  HS65_LH_BFX4 U8031 ( .A(n7233), .Z(n7231) );
  HS65_LH_BFX4 U8033 ( .A(n7234), .Z(n7233) );
  HS65_LH_BFX4 U8034 ( .A(n7235), .Z(n7234) );
  HS65_LH_BFX4 U8035 ( .A(n7236), .Z(n7235) );
  HS65_LH_BFX4 U8036 ( .A(n14577), .Z(n7236) );
  HS65_LH_BFX4 U8037 ( .A(n7238), .Z(n7237) );
  HS65_LH_BFX4 U8038 ( .A(n7239), .Z(n7238) );
  HS65_LH_BFX4 U8039 ( .A(n7240), .Z(n7239) );
  HS65_LH_BFX4 U8040 ( .A(n7241), .Z(n7240) );
  HS65_LH_BFX4 U8041 ( .A(n7242), .Z(n7241) );
  HS65_LH_BFX4 U8042 ( .A(n7243), .Z(n7242) );
  HS65_LH_BFX4 U8043 ( .A(n7244), .Z(n7243) );
  HS65_LH_BFX4 U8044 ( .A(n7245), .Z(n7244) );
  HS65_LH_BFX4 U8045 ( .A(n7246), .Z(n7245) );
  HS65_LH_BFX4 U8046 ( .A(n7247), .Z(n7246) );
  HS65_LH_BFX4 U8047 ( .A(n7248), .Z(n7247) );
  HS65_LH_BFX4 U8048 ( .A(n7249), .Z(n7248) );
  HS65_LH_BFX4 U8049 ( .A(n7250), .Z(n7249) );
  HS65_LH_BFX4 U8050 ( .A(n7251), .Z(n7250) );
  HS65_LH_BFX4 U8051 ( .A(n7252), .Z(n7251) );
  HS65_LH_BFX4 U8052 ( .A(n7253), .Z(n7252) );
  HS65_LH_BFX4 U8053 ( .A(n7254), .Z(n7253) );
  HS65_LH_BFX4 U8054 ( .A(n7255), .Z(n7254) );
  HS65_LH_BFX4 U8055 ( .A(n7256), .Z(n7255) );
  HS65_LH_BFX4 U8056 ( .A(n14181), .Z(n7256) );
  HS65_LH_BFX4 U8057 ( .A(n7258), .Z(n7257) );
  HS65_LH_BFX4 U8058 ( .A(n7259), .Z(n7258) );
  HS65_LH_BFX4 U8059 ( .A(n7260), .Z(n7259) );
  HS65_LH_BFX4 U8060 ( .A(n7261), .Z(n7260) );
  HS65_LH_BFX4 U8061 ( .A(n7262), .Z(n7261) );
  HS65_LH_BFX4 U8062 ( .A(n7263), .Z(n7262) );
  HS65_LH_BFX4 U8063 ( .A(n7264), .Z(n7263) );
  HS65_LH_BFX4 U8064 ( .A(n7265), .Z(n7264) );
  HS65_LH_BFX4 U8065 ( .A(n7266), .Z(n7265) );
  HS65_LH_BFX4 U8066 ( .A(n7267), .Z(n7266) );
  HS65_LH_BFX4 U8067 ( .A(n7268), .Z(n7267) );
  HS65_LH_BFX4 U8068 ( .A(n7269), .Z(n7268) );
  HS65_LH_BFX4 U8069 ( .A(n7270), .Z(n7269) );
  HS65_LH_BFX4 U8070 ( .A(n7271), .Z(n7270) );
  HS65_LH_BFX4 U8071 ( .A(n7272), .Z(n7271) );
  HS65_LH_BFX4 U8072 ( .A(n7273), .Z(n7272) );
  HS65_LH_BFX4 U8073 ( .A(n7274), .Z(n7273) );
  HS65_LH_BFX4 U8074 ( .A(n7275), .Z(n7274) );
  HS65_LH_BFX4 U8075 ( .A(n7276), .Z(n7275) );
  HS65_LH_BFX4 U8076 ( .A(n7277), .Z(n7276) );
  HS65_LH_BFX4 U8077 ( .A(n7278), .Z(n7277) );
  HS65_LH_BFX4 U8078 ( .A(n7279), .Z(n7278) );
  HS65_LH_BFX4 U8079 ( .A(n7280), .Z(n7279) );
  HS65_LH_BFX4 U8080 ( .A(n7281), .Z(n7280) );
  HS65_LH_BFX4 U8081 ( .A(n15644), .Z(n7281) );
  HS65_LH_BFX4 U8102 ( .A(n7304), .Z(n7302) );
  HS65_LH_BFX4 U8104 ( .A(n7306), .Z(n7304) );
  HS65_LH_BFX4 U8106 ( .A(n7308), .Z(n7306) );
  HS65_LH_BFX4 U8108 ( .A(n7310), .Z(n7308) );
  HS65_LH_BFX4 U8110 ( .A(n7312), .Z(n7310) );
  HS65_LH_BFX4 U8112 ( .A(n7314), .Z(n7312) );
  HS65_LH_BFX4 U8114 ( .A(n7316), .Z(n7314) );
  HS65_LH_BFX4 U8116 ( .A(n7317), .Z(n7316) );
  HS65_LH_BFX4 U8117 ( .A(n7318), .Z(n7317) );
  HS65_LH_BFX4 U8118 ( .A(n7319), .Z(n7318) );
  HS65_LH_BFX4 U8119 ( .A(n14607), .Z(n7319) );
  HS65_LH_BFX4 U8120 ( .A(n7321), .Z(n7320) );
  HS65_LH_BFX4 U8121 ( .A(n7322), .Z(n7321) );
  HS65_LH_BFX4 U8122 ( .A(n7323), .Z(n7322) );
  HS65_LH_BFX4 U8123 ( .A(n7324), .Z(n7323) );
  HS65_LH_BFX4 U8124 ( .A(n7325), .Z(n7324) );
  HS65_LH_BFX4 U8125 ( .A(n7326), .Z(n7325) );
  HS65_LH_BFX4 U8126 ( .A(n7327), .Z(n7326) );
  HS65_LH_BFX4 U8127 ( .A(n7328), .Z(n7327) );
  HS65_LH_BFX4 U8128 ( .A(n7329), .Z(n7328) );
  HS65_LH_BFX4 U8129 ( .A(n7330), .Z(n7329) );
  HS65_LH_BFX4 U8130 ( .A(n7331), .Z(n7330) );
  HS65_LH_BFX4 U8131 ( .A(n7332), .Z(n7331) );
  HS65_LH_BFX4 U8132 ( .A(n7333), .Z(n7332) );
  HS65_LH_BFX4 U8133 ( .A(n7334), .Z(n7333) );
  HS65_LH_BFX4 U8134 ( .A(n7335), .Z(n7334) );
  HS65_LH_BFX4 U8135 ( .A(n7336), .Z(n7335) );
  HS65_LH_BFX4 U8136 ( .A(n7337), .Z(n7336) );
  HS65_LH_BFX4 U8137 ( .A(n7338), .Z(n7337) );
  HS65_LH_BFX4 U8138 ( .A(n7339), .Z(n7338) );
  HS65_LH_BFX4 U8139 ( .A(n14178), .Z(n7339) );
  HS65_LH_BFX4 U8165 ( .A(n7368), .Z(n7365) );
  HS65_LH_BFX4 U8168 ( .A(n7371), .Z(n7368) );
  HS65_LH_BFX4 U8171 ( .A(n7374), .Z(n7371) );
  HS65_LH_BFX4 U8174 ( .A(n7377), .Z(n7374) );
  HS65_LH_BFX4 U8177 ( .A(n7380), .Z(n7377) );
  HS65_LH_BFX4 U8180 ( .A(n7383), .Z(n7380) );
  HS65_LH_BFX4 U8183 ( .A(n7386), .Z(n7383) );
  HS65_LH_BFX4 U8186 ( .A(n7389), .Z(n7386) );
  HS65_LH_BFX4 U8189 ( .A(n7392), .Z(n7389) );
  HS65_LH_BFX4 U8192 ( .A(n7395), .Z(n7392) );
  HS65_LH_BFX4 U8195 ( .A(n7398), .Z(n7395) );
  HS65_LH_BFX4 U8198 ( .A(n7401), .Z(n7398) );
  HS65_LH_BFX4 U8201 ( .A(n7404), .Z(n7401) );
  HS65_LH_BFX4 U8204 ( .A(n7407), .Z(n7404) );
  HS65_LH_BFX4 U8207 ( .A(n7410), .Z(n7407) );
  HS65_LH_BFX4 U8210 ( .A(n7413), .Z(n7410) );
  HS65_LH_BFX4 U8213 ( .A(n7416), .Z(n7413) );
  HS65_LH_BFX4 U8216 ( .A(n7418), .Z(n7416) );
  HS65_LH_BFX4 U8218 ( .A(n7420), .Z(n7418) );
  HS65_LH_BFX4 U8220 ( .A(n7422), .Z(n7420) );
  HS65_LH_BFX4 U8222 ( .A(n7424), .Z(n7422) );
  HS65_LH_BFX4 U8224 ( .A(n7425), .Z(n7424) );
  HS65_LH_BFX4 U8225 ( .A(n7426), .Z(n7425) );
  HS65_LH_BFX4 U8226 ( .A(n7427), .Z(n7426) );
  HS65_LH_BFX4 U8227 ( .A(\u_DataPath/u_idexreg/N38 ), .Z(n7427) );
  HS65_LH_BFX4 U8252 ( .A(n7453), .Z(n7452) );
  HS65_LH_BFX4 U8253 ( .A(n7454), .Z(n7453) );
  HS65_LH_BFX4 U8254 ( .A(n7455), .Z(n7454) );
  HS65_LH_BFX4 U8255 ( .A(n7456), .Z(n7455) );
  HS65_LH_BFX4 U8256 ( .A(n7457), .Z(n7456) );
  HS65_LH_BFX4 U8257 ( .A(n7458), .Z(n7457) );
  HS65_LH_BFX4 U8258 ( .A(n7459), .Z(n7458) );
  HS65_LH_BFX4 U8259 ( .A(n7460), .Z(n7459) );
  HS65_LH_BFX4 U8260 ( .A(n7461), .Z(n7460) );
  HS65_LH_BFX4 U8261 ( .A(n7462), .Z(n7461) );
  HS65_LH_BFX4 U8262 ( .A(n7463), .Z(n7462) );
  HS65_LH_BFX4 U8263 ( .A(n7464), .Z(n7463) );
  HS65_LH_BFX4 U8264 ( .A(n7465), .Z(n7464) );
  HS65_LH_BFX4 U8265 ( .A(n7466), .Z(n7465) );
  HS65_LH_BFX4 U8266 ( .A(n7467), .Z(n7466) );
  HS65_LH_BFX4 U8267 ( .A(n7468), .Z(n7467) );
  HS65_LH_BFX4 U8268 ( .A(n7469), .Z(n7468) );
  HS65_LH_BFX4 U8269 ( .A(n7470), .Z(n7469) );
  HS65_LH_BFX4 U8270 ( .A(n7471), .Z(n7470) );
  HS65_LH_BFX4 U8271 ( .A(n14175), .Z(n7471) );
  HS65_LH_BFX4 U8287 ( .A(n7488), .Z(n7487) );
  HS65_LH_BFX4 U8288 ( .A(n7489), .Z(n7488) );
  HS65_LH_BFX4 U8289 ( .A(n7490), .Z(n7489) );
  HS65_LH_BFX4 U8290 ( .A(n7491), .Z(n7490) );
  HS65_LH_BFX4 U8291 ( .A(n7492), .Z(n7491) );
  HS65_LH_BFX4 U8292 ( .A(n7493), .Z(n7492) );
  HS65_LH_BFX4 U8293 ( .A(n7494), .Z(n7493) );
  HS65_LH_BFX4 U8294 ( .A(n7495), .Z(n7494) );
  HS65_LH_BFX4 U8295 ( .A(n7496), .Z(n7495) );
  HS65_LH_BFX4 U8296 ( .A(n14695), .Z(n7496) );
  HS65_LH_BFX4 U8299 ( .A(n7502), .Z(n7499) );
  HS65_LH_BFX4 U8302 ( .A(n7505), .Z(n7502) );
  HS65_LH_BFX4 U8305 ( .A(n7508), .Z(n7505) );
  HS65_LH_BFX4 U8308 ( .A(n7511), .Z(n7508) );
  HS65_LH_BFX4 U8311 ( .A(n7514), .Z(n7511) );
  HS65_LH_BFX4 U8314 ( .A(n7517), .Z(n7514) );
  HS65_LH_BFX4 U8317 ( .A(n7519), .Z(n7517) );
  HS65_LH_BFX4 U8319 ( .A(n7522), .Z(n7519) );
  HS65_LH_BFX4 U8322 ( .A(n7525), .Z(n7522) );
  HS65_LH_BFX4 U8325 ( .A(n7528), .Z(n7525) );
  HS65_LH_BFX4 U8328 ( .A(n7531), .Z(n7528) );
  HS65_LH_BFX4 U8331 ( .A(n7534), .Z(n7531) );
  HS65_LH_BFX4 U8334 ( .A(n7537), .Z(n7534) );
  HS65_LH_BFX4 U8337 ( .A(n7540), .Z(n7537) );
  HS65_LH_BFX4 U8340 ( .A(n7543), .Z(n7540) );
  HS65_LH_BFX4 U8343 ( .A(n7546), .Z(n7543) );
  HS65_LH_BFX4 U8346 ( .A(n7549), .Z(n7546) );
  HS65_LH_BFX4 U8349 ( .A(n7551), .Z(n7549) );
  HS65_LH_BFX4 U8351 ( .A(n7553), .Z(n7551) );
  HS65_LH_BFX4 U8353 ( .A(n7555), .Z(n7553) );
  HS65_LH_BFX4 U8355 ( .A(n7556), .Z(n7555) );
  HS65_LH_BFX4 U8356 ( .A(n7557), .Z(n7556) );
  HS65_LH_BFX4 U8357 ( .A(n7558), .Z(n7557) );
  HS65_LH_BFX4 U8358 ( .A(\u_DataPath/u_idexreg/N30 ), .Z(n7558) );
  HS65_LH_BFX4 U8359 ( .A(n7560), .Z(n7559) );
  HS65_LH_BFX4 U8360 ( .A(n7561), .Z(n7560) );
  HS65_LH_BFX4 U8361 ( .A(n7562), .Z(n7561) );
  HS65_LH_BFX4 U8362 ( .A(n7563), .Z(n7562) );
  HS65_LH_BFX4 U8363 ( .A(n7564), .Z(n7563) );
  HS65_LH_BFX4 U8364 ( .A(n7565), .Z(n7564) );
  HS65_LH_BFX4 U8365 ( .A(n7566), .Z(n7565) );
  HS65_LH_BFX4 U8366 ( .A(n7567), .Z(n7566) );
  HS65_LH_BFX4 U8367 ( .A(n7568), .Z(n7567) );
  HS65_LH_BFX4 U8368 ( .A(n7569), .Z(n7568) );
  HS65_LH_BFX4 U8369 ( .A(n7570), .Z(n7569) );
  HS65_LH_BFX4 U8370 ( .A(n7571), .Z(n7570) );
  HS65_LH_BFX4 U8371 ( .A(n7572), .Z(n7571) );
  HS65_LH_BFX4 U8372 ( .A(n7573), .Z(n7572) );
  HS65_LH_BFX4 U8373 ( .A(n7574), .Z(n7573) );
  HS65_LH_BFX4 U8374 ( .A(n7575), .Z(n7574) );
  HS65_LH_BFX4 U8375 ( .A(n7576), .Z(n7575) );
  HS65_LH_BFX4 U8376 ( .A(n7577), .Z(n7576) );
  HS65_LH_BFX4 U8377 ( .A(n7578), .Z(n7577) );
  HS65_LH_BFX4 U8378 ( .A(n14172), .Z(n7578) );
  HS65_LH_BFX4 U8379 ( .A(n7580), .Z(n7579) );
  HS65_LH_BFX4 U8380 ( .A(n7581), .Z(n7580) );
  HS65_LH_BFX4 U8381 ( .A(n7582), .Z(n7581) );
  HS65_LH_BFX4 U8382 ( .A(n7583), .Z(n7582) );
  HS65_LH_BFX4 U8383 ( .A(n7584), .Z(n7583) );
  HS65_LH_BFX4 U8384 ( .A(n7585), .Z(n7584) );
  HS65_LH_BFX4 U8385 ( .A(n7586), .Z(n7585) );
  HS65_LH_BFX4 U8386 ( .A(n7587), .Z(n7586) );
  HS65_LH_BFX4 U8387 ( .A(n7588), .Z(n7587) );
  HS65_LH_BFX4 U8388 ( .A(n7589), .Z(n7588) );
  HS65_LH_BFX4 U8389 ( .A(n7590), .Z(n7589) );
  HS65_LH_BFX4 U8390 ( .A(n7591), .Z(n7590) );
  HS65_LH_BFX4 U8391 ( .A(n7592), .Z(n7591) );
  HS65_LH_BFX4 U8392 ( .A(n7593), .Z(n7592) );
  HS65_LH_BFX4 U8393 ( .A(n7594), .Z(n7593) );
  HS65_LH_BFX4 U8394 ( .A(n7595), .Z(n7594) );
  HS65_LH_BFX4 U8395 ( .A(n7596), .Z(n7595) );
  HS65_LH_BFX4 U8396 ( .A(n7597), .Z(n7596) );
  HS65_LH_BFX4 U8397 ( .A(n7598), .Z(n7597) );
  HS65_LH_BFX4 U8398 ( .A(n7599), .Z(n7598) );
  HS65_LH_BFX4 U8399 ( .A(n7600), .Z(n7599) );
  HS65_LH_BFX4 U8400 ( .A(n7601), .Z(n7600) );
  HS65_LH_BFX4 U8401 ( .A(n7602), .Z(n7601) );
  HS65_LH_BFX4 U8402 ( .A(n7603), .Z(n7602) );
  HS65_LH_BFX4 U8403 ( .A(n15650), .Z(n7603) );
  HS65_LH_BFX4 U8404 ( .A(n7606), .Z(n7604) );
  HS65_LH_BFX4 U8406 ( .A(n7608), .Z(n7606) );
  HS65_LH_BFX4 U8408 ( .A(n7610), .Z(n7608) );
  HS65_LH_BFX4 U8410 ( .A(n7612), .Z(n7610) );
  HS65_LH_BFX4 U8412 ( .A(n7614), .Z(n7612) );
  HS65_LH_BFX4 U8414 ( .A(n7616), .Z(n7614) );
  HS65_LH_BFX4 U8416 ( .A(n7618), .Z(n7616) );
  HS65_LH_BFX4 U8418 ( .A(n7620), .Z(n7618) );
  HS65_LH_BFX4 U8420 ( .A(n7622), .Z(n7620) );
  HS65_LH_BFX4 U8422 ( .A(n7624), .Z(n7622) );
  HS65_LH_BFX4 U8424 ( .A(n7626), .Z(n7624) );
  HS65_LH_BFX4 U8426 ( .A(n7628), .Z(n7626) );
  HS65_LH_BFX4 U8428 ( .A(n7630), .Z(n7628) );
  HS65_LH_BFX4 U8430 ( .A(n7632), .Z(n7630) );
  HS65_LH_BFX4 U8432 ( .A(n7634), .Z(n7632) );
  HS65_LH_BFX4 U8434 ( .A(n7636), .Z(n7634) );
  HS65_LH_BFX4 U8436 ( .A(n7638), .Z(n7636) );
  HS65_LH_BFX4 U8438 ( .A(n7639), .Z(n7638) );
  HS65_LH_BFX4 U8439 ( .A(n7640), .Z(n7639) );
  HS65_LH_BFX4 U8440 ( .A(n7641), .Z(n7640) );
  HS65_LH_BFX4 U8441 ( .A(n14721), .Z(n7641) );
  HS65_LH_BFX4 U8442 ( .A(n7643), .Z(n7642) );
  HS65_LH_BFX4 U8443 ( .A(n7644), .Z(n7643) );
  HS65_LH_BFX4 U8444 ( .A(n7645), .Z(n7644) );
  HS65_LH_BFX4 U8445 ( .A(n7646), .Z(n7645) );
  HS65_LH_BFX4 U8446 ( .A(n7647), .Z(n7646) );
  HS65_LH_BFX4 U8447 ( .A(n7648), .Z(n7647) );
  HS65_LH_BFX4 U8448 ( .A(n7649), .Z(n7648) );
  HS65_LH_BFX4 U8449 ( .A(n7650), .Z(n7649) );
  HS65_LH_BFX4 U8450 ( .A(n7651), .Z(n7650) );
  HS65_LH_BFX4 U8451 ( .A(n7652), .Z(n7651) );
  HS65_LH_BFX4 U8452 ( .A(n7653), .Z(n7652) );
  HS65_LH_BFX4 U8453 ( .A(n7654), .Z(n7653) );
  HS65_LH_BFX4 U8454 ( .A(n7655), .Z(n7654) );
  HS65_LH_BFX4 U8455 ( .A(n7656), .Z(n7655) );
  HS65_LH_BFX4 U8456 ( .A(n7657), .Z(n7656) );
  HS65_LH_BFX4 U8457 ( .A(n7658), .Z(n7657) );
  HS65_LH_BFX4 U8458 ( .A(n7659), .Z(n7658) );
  HS65_LH_BFX4 U8459 ( .A(n7660), .Z(n7659) );
  HS65_LH_BFX4 U8460 ( .A(n7661), .Z(n7660) );
  HS65_LH_BFX4 U8461 ( .A(n14169), .Z(n7661) );
  HS65_LH_BFX4 U8489 ( .A(n7692), .Z(n7689) );
  HS65_LH_BFX4 U8492 ( .A(n7695), .Z(n7692) );
  HS65_LH_BFX4 U8495 ( .A(n7698), .Z(n7695) );
  HS65_LH_BFX4 U8498 ( .A(n7701), .Z(n7698) );
  HS65_LH_BFX4 U8501 ( .A(n7704), .Z(n7701) );
  HS65_LH_BFX4 U8504 ( .A(n7706), .Z(n7704) );
  HS65_LH_BFX4 U8506 ( .A(n7709), .Z(n7706) );
  HS65_LH_BFX4 U8509 ( .A(n7712), .Z(n7709) );
  HS65_LH_BFX4 U8512 ( .A(n7715), .Z(n7712) );
  HS65_LH_BFX4 U8515 ( .A(n7718), .Z(n7715) );
  HS65_LH_BFX4 U8518 ( .A(n7721), .Z(n7718) );
  HS65_LH_BFX4 U8521 ( .A(n7724), .Z(n7721) );
  HS65_LH_BFX4 U8524 ( .A(n7727), .Z(n7724) );
  HS65_LH_BFX4 U8527 ( .A(n7730), .Z(n7727) );
  HS65_LH_BFX4 U8530 ( .A(n7733), .Z(n7730) );
  HS65_LH_BFX4 U8533 ( .A(n7736), .Z(n7733) );
  HS65_LH_BFX4 U8536 ( .A(n7739), .Z(n7736) );
  HS65_LH_BFX4 U8539 ( .A(n7742), .Z(n7739) );
  HS65_LH_BFX4 U8542 ( .A(n7744), .Z(n7742) );
  HS65_LH_BFX4 U8544 ( .A(n7746), .Z(n7744) );
  HS65_LH_BFX4 U8546 ( .A(n7747), .Z(n7746) );
  HS65_LH_BFX4 U8547 ( .A(n7748), .Z(n7747) );
  HS65_LH_BFX4 U8548 ( .A(n7749), .Z(n7748) );
  HS65_LH_BFX4 U8549 ( .A(\u_DataPath/u_idexreg/N34 ), .Z(n7749) );
  HS65_LH_BFX4 U8550 ( .A(n7751), .Z(n7750) );
  HS65_LH_BFX4 U8551 ( .A(n7752), .Z(n7751) );
  HS65_LH_BFX4 U8552 ( .A(n7753), .Z(n7752) );
  HS65_LH_BFX4 U8553 ( .A(n7754), .Z(n7753) );
  HS65_LH_BFX4 U8554 ( .A(n7755), .Z(n7754) );
  HS65_LH_BFX4 U8555 ( .A(n7756), .Z(n7755) );
  HS65_LH_BFX4 U8556 ( .A(n7757), .Z(n7756) );
  HS65_LH_BFX4 U8557 ( .A(n7758), .Z(n7757) );
  HS65_LH_BFX4 U8558 ( .A(n7759), .Z(n7758) );
  HS65_LH_BFX4 U8559 ( .A(n7760), .Z(n7759) );
  HS65_LH_BFX4 U8560 ( .A(n7761), .Z(n7760) );
  HS65_LH_BFX4 U8561 ( .A(n7762), .Z(n7761) );
  HS65_LH_BFX4 U8562 ( .A(n7763), .Z(n7762) );
  HS65_LH_BFX4 U8563 ( .A(n7764), .Z(n7763) );
  HS65_LH_BFX4 U8564 ( .A(n7765), .Z(n7764) );
  HS65_LH_BFX4 U8565 ( .A(n7766), .Z(n7765) );
  HS65_LH_BFX4 U8566 ( .A(n7767), .Z(n7766) );
  HS65_LH_BFX4 U8567 ( .A(n7768), .Z(n7767) );
  HS65_LH_BFX4 U8568 ( .A(n7769), .Z(n7768) );
  HS65_LH_BFX4 U8569 ( .A(n14166), .Z(n7769) );
  HS65_LH_BFX4 U8570 ( .A(n7771), .Z(n7770) );
  HS65_LH_BFX4 U8571 ( .A(n7772), .Z(n7771) );
  HS65_LH_BFX4 U8572 ( .A(n7773), .Z(n7772) );
  HS65_LH_BFX4 U8573 ( .A(n7774), .Z(n7773) );
  HS65_LH_BFX4 U8574 ( .A(n7775), .Z(n7774) );
  HS65_LH_BFX4 U8575 ( .A(n7776), .Z(n7775) );
  HS65_LH_BFX4 U8576 ( .A(n7777), .Z(n7776) );
  HS65_LH_BFX4 U8577 ( .A(n7778), .Z(n7777) );
  HS65_LH_BFX4 U8578 ( .A(n7779), .Z(n7778) );
  HS65_LH_BFX4 U8579 ( .A(n7780), .Z(n7779) );
  HS65_LH_BFX4 U8580 ( .A(n7781), .Z(n7780) );
  HS65_LH_BFX4 U8581 ( .A(n7782), .Z(n7781) );
  HS65_LH_BFX4 U8582 ( .A(n7783), .Z(n7782) );
  HS65_LH_BFX4 U8583 ( .A(n7784), .Z(n7783) );
  HS65_LH_BFX4 U8584 ( .A(n7785), .Z(n7784) );
  HS65_LH_BFX4 U8585 ( .A(n7786), .Z(n7785) );
  HS65_LH_BFX4 U8586 ( .A(n7787), .Z(n7786) );
  HS65_LH_BFX4 U8587 ( .A(n7788), .Z(n7787) );
  HS65_LH_BFX4 U8588 ( .A(n7789), .Z(n7788) );
  HS65_LH_BFX4 U8589 ( .A(n7790), .Z(n7789) );
  HS65_LH_BFX4 U8590 ( .A(n7791), .Z(n7790) );
  HS65_LH_BFX4 U8591 ( .A(n7792), .Z(n7791) );
  HS65_LH_BFX4 U8592 ( .A(n7793), .Z(n7792) );
  HS65_LH_BFX4 U8593 ( .A(n7794), .Z(n7793) );
  HS65_LH_BFX4 U8594 ( .A(n15656), .Z(n7794) );
  HS65_LH_BFX4 U8596 ( .A(n7798), .Z(n7796) );
  HS65_LH_BFX4 U8598 ( .A(n7800), .Z(n7798) );
  HS65_LH_BFX4 U8600 ( .A(n7802), .Z(n7800) );
  HS65_LH_BFX4 U8602 ( .A(n7804), .Z(n7802) );
  HS65_LH_BFX4 U8604 ( .A(n7806), .Z(n7804) );
  HS65_LH_BFX4 U8606 ( .A(n7808), .Z(n7806) );
  HS65_LH_BFX4 U8608 ( .A(n7810), .Z(n7808) );
  HS65_LH_BFX4 U8610 ( .A(n7812), .Z(n7810) );
  HS65_LH_BFX4 U8612 ( .A(n7814), .Z(n7812) );
  HS65_LH_BFX4 U8614 ( .A(n7816), .Z(n7814) );
  HS65_LH_BFX4 U8616 ( .A(n7818), .Z(n7816) );
  HS65_LH_BFX4 U8618 ( .A(n7820), .Z(n7818) );
  HS65_LH_BFX4 U8620 ( .A(n7822), .Z(n7820) );
  HS65_LH_BFX4 U8622 ( .A(n7824), .Z(n7822) );
  HS65_LH_BFX4 U8624 ( .A(n7826), .Z(n7824) );
  HS65_LH_BFX4 U8626 ( .A(n7828), .Z(n7826) );
  HS65_LH_BFX4 U8628 ( .A(n7830), .Z(n7828) );
  HS65_LH_BFX4 U8630 ( .A(n7832), .Z(n7830) );
  HS65_LH_BFX4 U8632 ( .A(n7833), .Z(n7832) );
  HS65_LH_BFX4 U8633 ( .A(n7834), .Z(n7833) );
  HS65_LH_BFX4 U8634 ( .A(n14801), .Z(n7834) );
  HS65_LH_BFX4 U8635 ( .A(n7836), .Z(n7835) );
  HS65_LH_BFX4 U8636 ( .A(n7837), .Z(n7836) );
  HS65_LH_BFX4 U8637 ( .A(n7838), .Z(n7837) );
  HS65_LH_BFX4 U8638 ( .A(n7839), .Z(n7838) );
  HS65_LH_BFX4 U8639 ( .A(n7840), .Z(n7839) );
  HS65_LH_BFX4 U8640 ( .A(n7841), .Z(n7840) );
  HS65_LH_BFX4 U8641 ( .A(n7842), .Z(n7841) );
  HS65_LH_BFX4 U8642 ( .A(n7843), .Z(n7842) );
  HS65_LH_BFX4 U8643 ( .A(n7844), .Z(n7843) );
  HS65_LH_BFX4 U8644 ( .A(n7845), .Z(n7844) );
  HS65_LH_BFX4 U8645 ( .A(n7846), .Z(n7845) );
  HS65_LH_BFX4 U8646 ( .A(n7847), .Z(n7846) );
  HS65_LH_BFX4 U8647 ( .A(n7848), .Z(n7847) );
  HS65_LH_BFX4 U8648 ( .A(n7849), .Z(n7848) );
  HS65_LH_BFX4 U8649 ( .A(n7850), .Z(n7849) );
  HS65_LH_BFX4 U8650 ( .A(n7851), .Z(n7850) );
  HS65_LH_BFX4 U8651 ( .A(n7852), .Z(n7851) );
  HS65_LH_BFX4 U8652 ( .A(n7853), .Z(n7852) );
  HS65_LH_BFX4 U8653 ( .A(n7854), .Z(n7853) );
  HS65_LH_BFX4 U8654 ( .A(n14163), .Z(n7854) );
  HS65_LH_BFX4 U8682 ( .A(n7885), .Z(n7882) );
  HS65_LH_BFX4 U8685 ( .A(n7888), .Z(n7885) );
  HS65_LH_BFX4 U8688 ( .A(n7891), .Z(n7888) );
  HS65_LH_BFX4 U8691 ( .A(n7894), .Z(n7891) );
  HS65_LH_BFX4 U8694 ( .A(n7897), .Z(n7894) );
  HS65_LH_BFX4 U8697 ( .A(n7900), .Z(n7897) );
  HS65_LH_BFX4 U8700 ( .A(n7903), .Z(n7900) );
  HS65_LH_BFX4 U8703 ( .A(n7906), .Z(n7903) );
  HS65_LH_BFX4 U8706 ( .A(n7909), .Z(n7906) );
  HS65_LH_BFX4 U8709 ( .A(n7912), .Z(n7909) );
  HS65_LH_BFX4 U8712 ( .A(n7915), .Z(n7912) );
  HS65_LH_BFX4 U8715 ( .A(n7918), .Z(n7915) );
  HS65_LH_BFX4 U8718 ( .A(n7921), .Z(n7918) );
  HS65_LH_BFX4 U8721 ( .A(n7924), .Z(n7921) );
  HS65_LH_BFX4 U8724 ( .A(n7926), .Z(n7924) );
  HS65_LH_BFX4 U8726 ( .A(n7929), .Z(n7926) );
  HS65_LH_BFX4 U8729 ( .A(n7932), .Z(n7929) );
  HS65_LH_BFX4 U8732 ( .A(n7934), .Z(n7932) );
  HS65_LH_BFX4 U8734 ( .A(n7936), .Z(n7934) );
  HS65_LH_BFX4 U8736 ( .A(n7938), .Z(n7936) );
  HS65_LH_BFX4 U8738 ( .A(n7939), .Z(n7938) );
  HS65_LH_BFX4 U8739 ( .A(n7940), .Z(n7939) );
  HS65_LH_BFX4 U8740 ( .A(n7941), .Z(n7940) );
  HS65_LH_BFX4 U8741 ( .A(\u_DataPath/u_idexreg/N33 ), .Z(n7941) );
  HS65_LH_BFX4 U8742 ( .A(n7943), .Z(n7942) );
  HS65_LH_BFX4 U8743 ( .A(n7944), .Z(n7943) );
  HS65_LH_BFX4 U8744 ( .A(n7945), .Z(n7944) );
  HS65_LH_BFX4 U8745 ( .A(n7946), .Z(n7945) );
  HS65_LH_BFX4 U8746 ( .A(n7947), .Z(n7946) );
  HS65_LH_BFX4 U8747 ( .A(n7948), .Z(n7947) );
  HS65_LH_BFX4 U8748 ( .A(n7949), .Z(n7948) );
  HS65_LH_BFX4 U8749 ( .A(n7950), .Z(n7949) );
  HS65_LH_BFX4 U8750 ( .A(n7951), .Z(n7950) );
  HS65_LH_BFX4 U8751 ( .A(n7952), .Z(n7951) );
  HS65_LH_BFX4 U8752 ( .A(n7953), .Z(n7952) );
  HS65_LH_BFX4 U8753 ( .A(n7954), .Z(n7953) );
  HS65_LH_BFX4 U8754 ( .A(n7955), .Z(n7954) );
  HS65_LH_BFX4 U8755 ( .A(n7956), .Z(n7955) );
  HS65_LH_BFX4 U8756 ( .A(n7957), .Z(n7956) );
  HS65_LH_BFX4 U8757 ( .A(n7958), .Z(n7957) );
  HS65_LH_BFX4 U8758 ( .A(n7959), .Z(n7958) );
  HS65_LH_BFX4 U8759 ( .A(n7960), .Z(n7959) );
  HS65_LH_BFX4 U8760 ( .A(n7961), .Z(n7960) );
  HS65_LH_BFX4 U8761 ( .A(n14160), .Z(n7961) );
  HS65_LH_CNIVX3 U8787 ( .A(\u_DataPath/pc_4_to_ex_i [28]), .Z(n7987) );
  HS65_LH_CNIVX3 U8788 ( .A(n7987), .Z(n7988) );
  HS65_LH_BFX4 U8789 ( .A(n7991), .Z(n7989) );
  HS65_LH_BFX4 U8791 ( .A(n7994), .Z(n7991) );
  HS65_LH_BFX4 U8794 ( .A(n7997), .Z(n7994) );
  HS65_LH_BFX4 U8797 ( .A(n8000), .Z(n7997) );
  HS65_LH_BFX4 U8800 ( .A(n8003), .Z(n8000) );
  HS65_LH_BFX4 U8803 ( .A(n8006), .Z(n8003) );
  HS65_LH_BFX4 U8806 ( .A(n8009), .Z(n8006) );
  HS65_LH_BFX4 U8809 ( .A(n8012), .Z(n8009) );
  HS65_LH_BFX4 U8812 ( .A(n8015), .Z(n8012) );
  HS65_LH_BFX4 U8815 ( .A(n8018), .Z(n8015) );
  HS65_LH_BFX4 U8818 ( .A(n8021), .Z(n8018) );
  HS65_LH_BFX4 U8821 ( .A(n8024), .Z(n8021) );
  HS65_LH_BFX4 U8824 ( .A(n8027), .Z(n8024) );
  HS65_LH_BFX4 U8827 ( .A(n8030), .Z(n8027) );
  HS65_LH_BFX4 U8830 ( .A(n8033), .Z(n8030) );
  HS65_LH_BFX4 U8833 ( .A(n8036), .Z(n8033) );
  HS65_LH_BFX4 U8836 ( .A(n8039), .Z(n8036) );
  HS65_LH_BFX4 U8839 ( .A(n8041), .Z(n8039) );
  HS65_LH_BFX4 U8841 ( .A(n8043), .Z(n8041) );
  HS65_LH_BFX4 U8843 ( .A(n8045), .Z(n8043) );
  HS65_LH_BFX4 U8845 ( .A(n8047), .Z(n8045) );
  HS65_LH_BFX4 U8847 ( .A(n8048), .Z(n8047) );
  HS65_LH_BFX4 U8848 ( .A(n8049), .Z(n8048) );
  HS65_LH_BFX4 U8849 ( .A(n8050), .Z(n8049) );
  HS65_LH_BFX4 U8850 ( .A(\u_DataPath/u_idexreg/N37 ), .Z(n8050) );
  HS65_LH_BFX4 U8851 ( .A(n8052), .Z(n8051) );
  HS65_LH_BFX4 U8852 ( .A(n8053), .Z(n8052) );
  HS65_LH_BFX4 U8853 ( .A(n8054), .Z(n8053) );
  HS65_LH_BFX4 U8854 ( .A(n8055), .Z(n8054) );
  HS65_LH_BFX4 U8855 ( .A(n8056), .Z(n8055) );
  HS65_LH_BFX4 U8856 ( .A(n8057), .Z(n8056) );
  HS65_LH_BFX4 U8857 ( .A(n8058), .Z(n8057) );
  HS65_LH_BFX4 U8858 ( .A(n8059), .Z(n8058) );
  HS65_LH_BFX4 U8859 ( .A(n8060), .Z(n8059) );
  HS65_LH_BFX4 U8860 ( .A(n8061), .Z(n8060) );
  HS65_LH_BFX4 U8861 ( .A(n8062), .Z(n8061) );
  HS65_LH_BFX4 U8862 ( .A(n8063), .Z(n8062) );
  HS65_LH_BFX4 U8863 ( .A(n8064), .Z(n8063) );
  HS65_LH_BFX4 U8864 ( .A(n8065), .Z(n8064) );
  HS65_LH_BFX4 U8865 ( .A(n8066), .Z(n8065) );
  HS65_LH_BFX4 U8866 ( .A(n8067), .Z(n8066) );
  HS65_LH_BFX4 U8867 ( .A(n8068), .Z(n8067) );
  HS65_LH_BFX4 U8868 ( .A(n8069), .Z(n8068) );
  HS65_LH_BFX4 U8869 ( .A(n8070), .Z(n8069) );
  HS65_LH_BFX4 U8870 ( .A(n14157), .Z(n8070) );
  HS65_LH_BFX4 U8893 ( .A(n8094), .Z(n8093) );
  HS65_LH_BFX4 U8894 ( .A(n8095), .Z(n8094) );
  HS65_LH_BFX4 U8895 ( .A(n14877), .Z(n8095) );
  HS65_LH_CNIVX3 U8896 ( .A(\u_DataPath/pc_4_to_ex_i [22]), .Z(n8096) );
  HS65_LH_CNIVX3 U8897 ( .A(n8096), .Z(n8097) );
  HS65_LH_BFX4 U8898 ( .A(n8100), .Z(n8098) );
  HS65_LH_BFX4 U8900 ( .A(n8103), .Z(n8100) );
  HS65_LH_BFX4 U8903 ( .A(n8106), .Z(n8103) );
  HS65_LH_BFX4 U8906 ( .A(n8109), .Z(n8106) );
  HS65_LH_BFX4 U8909 ( .A(n8112), .Z(n8109) );
  HS65_LH_BFX4 U8912 ( .A(n8115), .Z(n8112) );
  HS65_LH_BFX4 U8915 ( .A(n8118), .Z(n8115) );
  HS65_LH_BFX4 U8918 ( .A(n8121), .Z(n8118) );
  HS65_LH_BFX4 U8921 ( .A(n8124), .Z(n8121) );
  HS65_LH_BFX4 U8924 ( .A(n8127), .Z(n8124) );
  HS65_LH_BFX4 U8927 ( .A(n8130), .Z(n8127) );
  HS65_LH_BFX4 U8930 ( .A(n8133), .Z(n8130) );
  HS65_LH_BFX4 U8933 ( .A(n8136), .Z(n8133) );
  HS65_LH_BFX4 U8936 ( .A(n8139), .Z(n8136) );
  HS65_LH_BFX4 U8939 ( .A(n8142), .Z(n8139) );
  HS65_LH_BFX4 U8942 ( .A(n8145), .Z(n8142) );
  HS65_LH_BFX4 U8945 ( .A(n8147), .Z(n8145) );
  HS65_LH_BFX4 U8947 ( .A(n8149), .Z(n8147) );
  HS65_LH_BFX4 U8949 ( .A(n8151), .Z(n8149) );
  HS65_LH_BFX4 U8951 ( .A(n8153), .Z(n8151) );
  HS65_LH_BFX4 U8953 ( .A(n8155), .Z(n8153) );
  HS65_LH_BFX4 U8955 ( .A(n8156), .Z(n8155) );
  HS65_LH_BFX4 U8956 ( .A(n8157), .Z(n8156) );
  HS65_LH_BFX4 U8957 ( .A(n8158), .Z(n8157) );
  HS65_LH_BFX4 U8958 ( .A(\u_DataPath/u_idexreg/N31 ), .Z(n8158) );
  HS65_LH_BFX4 U8998 ( .A(n8200), .Z(n8198) );
  HS65_LH_BFX4 U9000 ( .A(n8202), .Z(n8200) );
  HS65_LH_BFX4 U9002 ( .A(n8204), .Z(n8202) );
  HS65_LH_BFX4 U9004 ( .A(n8206), .Z(n8204) );
  HS65_LH_BFX4 U9006 ( .A(n8208), .Z(n8206) );
  HS65_LH_BFX4 U9008 ( .A(n8210), .Z(n8208) );
  HS65_LH_BFX4 U9010 ( .A(n8212), .Z(n8210) );
  HS65_LH_BFX4 U9012 ( .A(n8214), .Z(n8212) );
  HS65_LH_BFX4 U9014 ( .A(n8216), .Z(n8214) );
  HS65_LH_BFX4 U9016 ( .A(n8218), .Z(n8216) );
  HS65_LH_BFX4 U9018 ( .A(n8222), .Z(n8218) );
  HS65_LH_BFX4 U9019 ( .A(\u_DataPath/data_read_ex_1_i [4]), .Z(n8219) );
  HS65_LH_BFX4 U9022 ( .A(n8223), .Z(n8222) );
  HS65_LH_BFX4 U9023 ( .A(n8224), .Z(n8223) );
  HS65_LH_BFX4 U9024 ( .A(n8225), .Z(n8224) );
  HS65_LH_BFX4 U9025 ( .A(n14909), .Z(n8225) );
  HS65_LH_BFX4 U9026 ( .A(n8227), .Z(n8226) );
  HS65_LH_BFX4 U9027 ( .A(n8228), .Z(n8227) );
  HS65_LH_BFX4 U9028 ( .A(n8229), .Z(n8228) );
  HS65_LH_BFX4 U9029 ( .A(n8230), .Z(n8229) );
  HS65_LH_BFX4 U9030 ( .A(n8231), .Z(n8230) );
  HS65_LH_BFX4 U9031 ( .A(n8232), .Z(n8231) );
  HS65_LH_BFX4 U9032 ( .A(n8233), .Z(n8232) );
  HS65_LH_BFX4 U9033 ( .A(n8234), .Z(n8233) );
  HS65_LH_BFX4 U9034 ( .A(n8235), .Z(n8234) );
  HS65_LH_BFX4 U9035 ( .A(n8236), .Z(n8235) );
  HS65_LH_BFX4 U9036 ( .A(n8237), .Z(n8236) );
  HS65_LH_BFX4 U9037 ( .A(n8238), .Z(n8237) );
  HS65_LH_BFX4 U9038 ( .A(n8239), .Z(n8238) );
  HS65_LH_BFX4 U9039 ( .A(n8240), .Z(n8239) );
  HS65_LH_BFX4 U9040 ( .A(n8241), .Z(n8240) );
  HS65_LH_BFX4 U9041 ( .A(n8242), .Z(n8241) );
  HS65_LH_BFX4 U9042 ( .A(n8243), .Z(n8242) );
  HS65_LH_BFX4 U9043 ( .A(n8244), .Z(n8243) );
  HS65_LH_BFX4 U9044 ( .A(n8245), .Z(n8244) );
  HS65_LH_BFX4 U9045 ( .A(n14223), .Z(n8245) );
  HS65_LH_BFX4 U9046 ( .A(n8247), .Z(n8246) );
  HS65_LH_BFX4 U9047 ( .A(n8248), .Z(n8247) );
  HS65_LH_BFX4 U9048 ( .A(n8249), .Z(n8248) );
  HS65_LH_BFX4 U9049 ( .A(n8250), .Z(n8249) );
  HS65_LH_BFX4 U9050 ( .A(n8251), .Z(n8250) );
  HS65_LH_BFX4 U9051 ( .A(n8252), .Z(n8251) );
  HS65_LH_BFX4 U9052 ( .A(n8253), .Z(n8252) );
  HS65_LH_BFX4 U9053 ( .A(n8254), .Z(n8253) );
  HS65_LH_BFX4 U9054 ( .A(n8255), .Z(n8254) );
  HS65_LH_BFX4 U9055 ( .A(n8256), .Z(n8255) );
  HS65_LH_BFX4 U9056 ( .A(n8257), .Z(n8256) );
  HS65_LH_BFX4 U9057 ( .A(n8258), .Z(n8257) );
  HS65_LH_BFX4 U9058 ( .A(n8259), .Z(n8258) );
  HS65_LH_BFX4 U9059 ( .A(n8260), .Z(n8259) );
  HS65_LH_BFX4 U9060 ( .A(n8261), .Z(n8260) );
  HS65_LH_BFX4 U9061 ( .A(n8262), .Z(n8261) );
  HS65_LH_BFX4 U9062 ( .A(n8263), .Z(n8262) );
  HS65_LH_BFX4 U9063 ( .A(n8264), .Z(n8263) );
  HS65_LH_BFX4 U9064 ( .A(n8265), .Z(n8264) );
  HS65_LH_BFX4 U9065 ( .A(n8266), .Z(n8265) );
  HS65_LH_BFX4 U9066 ( .A(n8267), .Z(n8266) );
  HS65_LH_BFX4 U9067 ( .A(n8268), .Z(n8267) );
  HS65_LH_BFX4 U9068 ( .A(n8269), .Z(n8268) );
  HS65_LH_BFX4 U9069 ( .A(n8270), .Z(n8269) );
  HS65_LH_BFX4 U9070 ( .A(n15658), .Z(n8270) );
  HS65_LH_BFX4 U9072 ( .A(n8274), .Z(n8272) );
  HS65_LH_BFX4 U9074 ( .A(n8276), .Z(n8274) );
  HS65_LH_BFX4 U9076 ( .A(n8278), .Z(n8276) );
  HS65_LH_BFX4 U9078 ( .A(n8280), .Z(n8278) );
  HS65_LH_BFX4 U9080 ( .A(n8282), .Z(n8280) );
  HS65_LH_BFX4 U9082 ( .A(n8284), .Z(n8282) );
  HS65_LH_BFX4 U9084 ( .A(n8286), .Z(n8284) );
  HS65_LH_BFX4 U9086 ( .A(n8288), .Z(n8286) );
  HS65_LH_BFX4 U9088 ( .A(n8290), .Z(n8288) );
  HS65_LH_BFX4 U9090 ( .A(n8292), .Z(n8290) );
  HS65_LH_BFX4 U9092 ( .A(n8294), .Z(n8292) );
  HS65_LH_BFX4 U9094 ( .A(n8296), .Z(n8294) );
  HS65_LH_BFX4 U9096 ( .A(n8298), .Z(n8296) );
  HS65_LH_BFX4 U9098 ( .A(n8300), .Z(n8298) );
  HS65_LH_BFX4 U9100 ( .A(n8302), .Z(n8300) );
  HS65_LH_BFX4 U9102 ( .A(n8304), .Z(n8302) );
  HS65_LH_BFX4 U9104 ( .A(n8305), .Z(n8304) );
  HS65_LH_BFX4 U9105 ( .A(n8306), .Z(n8305) );
  HS65_LH_BFX4 U9106 ( .A(n8307), .Z(n8306) );
  HS65_LH_BFX4 U9107 ( .A(n8308), .Z(n8307) );
  HS65_LH_BFX4 U9108 ( .A(n14942), .Z(n8308) );
  HS65_LH_BFX4 U9111 ( .A(n8313), .Z(n8311) );
  HS65_LH_BFX4 U9113 ( .A(n8315), .Z(n8313) );
  HS65_LH_BFX4 U9115 ( .A(n8316), .Z(n8315) );
  HS65_LH_BFX4 U9116 ( .A(n8318), .Z(n8316) );
  HS65_LH_BFX4 U9118 ( .A(n8320), .Z(n8318) );
  HS65_LH_BFX4 U9120 ( .A(n8322), .Z(n8320) );
  HS65_LH_BFX4 U9122 ( .A(n8324), .Z(n8322) );
  HS65_LH_BFX4 U9124 ( .A(n8325), .Z(n8324) );
  HS65_LH_BFX4 U9125 ( .A(n8326), .Z(n8325) );
  HS65_LH_BFX4 U9126 ( .A(n8327), .Z(n8326) );
  HS65_LH_BFX4 U9127 ( .A(n8328), .Z(n8327) );
  HS65_LH_BFX4 U9128 ( .A(n8329), .Z(n8328) );
  HS65_LH_BFX4 U9129 ( .A(n8330), .Z(n8329) );
  HS65_LH_BFX4 U9130 ( .A(n8331), .Z(n8330) );
  HS65_LH_BFX4 U9131 ( .A(n8332), .Z(n8331) );
  HS65_LH_BFX4 U9132 ( .A(n8333), .Z(n8332) );
  HS65_LH_BFX4 U9133 ( .A(n8334), .Z(n8333) );
  HS65_LH_BFX4 U9134 ( .A(n8335), .Z(n8334) );
  HS65_LH_BFX4 U9135 ( .A(n8336), .Z(n8335) );
  HS65_LH_BFX4 U9136 ( .A(n14154), .Z(n8336) );
  HS65_LH_BFX4 U9137 ( .A(n8338), .Z(n8337) );
  HS65_LH_BFX4 U9138 ( .A(n8339), .Z(n8338) );
  HS65_LH_BFX4 U9139 ( .A(n8340), .Z(n8339) );
  HS65_LH_BFX4 U9140 ( .A(n8341), .Z(n8340) );
  HS65_LH_BFX4 U9141 ( .A(n8342), .Z(n8341) );
  HS65_LH_BFX4 U9142 ( .A(n8343), .Z(n8342) );
  HS65_LH_BFX4 U9143 ( .A(n8344), .Z(n8343) );
  HS65_LH_BFX4 U9144 ( .A(n8345), .Z(n8344) );
  HS65_LH_BFX4 U9145 ( .A(n8346), .Z(n8345) );
  HS65_LH_BFX4 U9146 ( .A(n8347), .Z(n8346) );
  HS65_LH_BFX4 U9147 ( .A(n8348), .Z(n8347) );
  HS65_LH_BFX4 U9148 ( .A(n8349), .Z(n8348) );
  HS65_LH_BFX4 U9149 ( .A(n8350), .Z(n8349) );
  HS65_LH_BFX4 U9150 ( .A(n8351), .Z(n8350) );
  HS65_LH_BFX4 U9151 ( .A(n8352), .Z(n8351) );
  HS65_LH_BFX4 U9152 ( .A(n8353), .Z(n8352) );
  HS65_LH_BFX4 U9153 ( .A(n8354), .Z(n8353) );
  HS65_LH_BFX4 U9154 ( .A(n8355), .Z(n8354) );
  HS65_LH_BFX4 U9155 ( .A(n8356), .Z(n8355) );
  HS65_LH_BFX4 U9156 ( .A(n8357), .Z(n8356) );
  HS65_LH_BFX4 U9157 ( .A(n8358), .Z(n8357) );
  HS65_LH_BFX4 U9158 ( .A(n8359), .Z(n8358) );
  HS65_LH_BFX4 U9159 ( .A(n8360), .Z(n8359) );
  HS65_LH_BFX4 U9160 ( .A(n8361), .Z(n8360) );
  HS65_LH_BFX4 U9161 ( .A(n15646), .Z(n8361) );
  HS65_LH_CNIVX3 U9162 ( .A(\u_DataPath/pc_4_to_ex_i [8]), .Z(n8362) );
  HS65_LH_CNIVX3 U9163 ( .A(n8362), .Z(n8363) );
  HS65_LH_BFX4 U9166 ( .A(n8368), .Z(n8366) );
  HS65_LH_BFX4 U9168 ( .A(n8370), .Z(n8368) );
  HS65_LH_BFX4 U9170 ( .A(n8372), .Z(n8370) );
  HS65_LH_BFX4 U9172 ( .A(n8374), .Z(n8372) );
  HS65_LH_BFX4 U9174 ( .A(n8376), .Z(n8374) );
  HS65_LH_BFX4 U9176 ( .A(n8378), .Z(n8376) );
  HS65_LH_BFX4 U9178 ( .A(n8380), .Z(n8378) );
  HS65_LH_BFX4 U9180 ( .A(n8382), .Z(n8380) );
  HS65_LH_BFX4 U9182 ( .A(n8384), .Z(n8382) );
  HS65_LH_BFX4 U9184 ( .A(n8386), .Z(n8384) );
  HS65_LH_BFX4 U9186 ( .A(n8388), .Z(n8386) );
  HS65_LH_BFX4 U9188 ( .A(n8390), .Z(n8388) );
  HS65_LH_BFX4 U9190 ( .A(n8392), .Z(n8390) );
  HS65_LH_BFX4 U9192 ( .A(n8394), .Z(n8392) );
  HS65_LH_BFX4 U9194 ( .A(n8396), .Z(n8394) );
  HS65_LH_BFX4 U9196 ( .A(n8398), .Z(n8396) );
  HS65_LH_BFX4 U9198 ( .A(n8399), .Z(n8398) );
  HS65_LH_BFX4 U9199 ( .A(n8400), .Z(n8399) );
  HS65_LH_BFX4 U9200 ( .A(n8401), .Z(n8400) );
  HS65_LH_BFX4 U9201 ( .A(n14964), .Z(n8401) );
  HS65_LH_BFX4 U9202 ( .A(n8403), .Z(n8402) );
  HS65_LH_BFX4 U9203 ( .A(n8404), .Z(n8403) );
  HS65_LH_BFX4 U9204 ( .A(n8405), .Z(n8404) );
  HS65_LH_BFX4 U9205 ( .A(n8406), .Z(n8405) );
  HS65_LH_BFX4 U9206 ( .A(n8407), .Z(n8406) );
  HS65_LH_BFX4 U9207 ( .A(n8408), .Z(n8407) );
  HS65_LH_BFX4 U9208 ( .A(n8409), .Z(n8408) );
  HS65_LH_BFX4 U9209 ( .A(n8410), .Z(n8409) );
  HS65_LH_BFX4 U9210 ( .A(n8411), .Z(n8410) );
  HS65_LH_BFX4 U9211 ( .A(n8412), .Z(n8411) );
  HS65_LH_BFX4 U9212 ( .A(n8413), .Z(n8412) );
  HS65_LH_BFX4 U9213 ( .A(n8414), .Z(n8413) );
  HS65_LH_BFX4 U9214 ( .A(n8415), .Z(n8414) );
  HS65_LH_BFX4 U9215 ( .A(n8416), .Z(n8415) );
  HS65_LH_BFX4 U9216 ( .A(n8417), .Z(n8416) );
  HS65_LH_BFX4 U9217 ( .A(n8418), .Z(n8417) );
  HS65_LH_BFX4 U9218 ( .A(n8419), .Z(n8418) );
  HS65_LH_BFX4 U9219 ( .A(n8420), .Z(n8419) );
  HS65_LH_BFX4 U9220 ( .A(n8421), .Z(n8420) );
  HS65_LH_BFX4 U9221 ( .A(n14151), .Z(n8421) );
  HS65_LH_BFX4 U9239 ( .A(n8440), .Z(n8439) );
  HS65_LH_BFX4 U9240 ( .A(n8441), .Z(n8440) );
  HS65_LH_BFX4 U9241 ( .A(n8442), .Z(n8441) );
  HS65_LH_BFX4 U9242 ( .A(n8443), .Z(n8442) );
  HS65_LH_BFX4 U9243 ( .A(n8444), .Z(n8443) );
  HS65_LH_BFX4 U9244 ( .A(n8445), .Z(n8444) );
  HS65_LH_BFX4 U9245 ( .A(n8446), .Z(n8445) );
  HS65_LH_BFX4 U9246 ( .A(n15697), .Z(n8446) );
  HS65_LH_CNIVX3 U9247 ( .A(\u_DataPath/pc_4_to_ex_i [20]), .Z(n8447) );
  HS65_LH_CNIVX3 U9248 ( .A(n8447), .Z(n8448) );
  HS65_LH_BFX4 U9249 ( .A(n8451), .Z(n8449) );
  HS65_LH_BFX4 U9251 ( .A(n8454), .Z(n8451) );
  HS65_LH_BFX4 U9254 ( .A(n8457), .Z(n8454) );
  HS65_LH_BFX4 U9257 ( .A(n8460), .Z(n8457) );
  HS65_LH_BFX4 U9260 ( .A(n8463), .Z(n8460) );
  HS65_LH_BFX4 U9263 ( .A(n8466), .Z(n8463) );
  HS65_LH_BFX4 U9266 ( .A(n8469), .Z(n8466) );
  HS65_LH_BFX4 U9269 ( .A(n8472), .Z(n8469) );
  HS65_LH_BFX4 U9272 ( .A(n8475), .Z(n8472) );
  HS65_LH_BFX4 U9275 ( .A(n8478), .Z(n8475) );
  HS65_LH_BFX4 U9278 ( .A(n8481), .Z(n8478) );
  HS65_LH_BFX4 U9281 ( .A(n8484), .Z(n8481) );
  HS65_LH_BFX4 U9284 ( .A(n8487), .Z(n8484) );
  HS65_LH_BFX4 U9287 ( .A(n8490), .Z(n8487) );
  HS65_LH_BFX4 U9290 ( .A(n8493), .Z(n8490) );
  HS65_LH_BFX4 U9293 ( .A(n8496), .Z(n8493) );
  HS65_LH_BFX4 U9296 ( .A(n8499), .Z(n8496) );
  HS65_LH_BFX4 U9299 ( .A(n8501), .Z(n8499) );
  HS65_LH_BFX4 U9301 ( .A(n8503), .Z(n8501) );
  HS65_LH_BFX4 U9303 ( .A(n8505), .Z(n8503) );
  HS65_LH_BFX4 U9305 ( .A(n8507), .Z(n8505) );
  HS65_LH_BFX4 U9307 ( .A(n8508), .Z(n8507) );
  HS65_LH_BFX4 U9308 ( .A(n8509), .Z(n8508) );
  HS65_LH_BFX4 U9309 ( .A(n8510), .Z(n8509) );
  HS65_LH_BFX4 U9310 ( .A(\u_DataPath/u_idexreg/N29 ), .Z(n8510) );
  HS65_LH_BFX4 U9311 ( .A(n8512), .Z(n8511) );
  HS65_LH_BFX4 U9312 ( .A(n8513), .Z(n8512) );
  HS65_LH_BFX4 U9313 ( .A(n8514), .Z(n8513) );
  HS65_LH_BFX4 U9314 ( .A(n8515), .Z(n8514) );
  HS65_LH_BFX4 U9315 ( .A(n8516), .Z(n8515) );
  HS65_LH_BFX4 U9316 ( .A(n8517), .Z(n8516) );
  HS65_LH_BFX4 U9317 ( .A(n8518), .Z(n8517) );
  HS65_LH_BFX4 U9318 ( .A(n8519), .Z(n8518) );
  HS65_LH_BFX4 U9319 ( .A(n8520), .Z(n8519) );
  HS65_LH_BFX4 U9320 ( .A(n8521), .Z(n8520) );
  HS65_LH_BFX4 U9321 ( .A(n8522), .Z(n8521) );
  HS65_LH_BFX4 U9322 ( .A(n8523), .Z(n8522) );
  HS65_LH_BFX4 U9323 ( .A(n8524), .Z(n8523) );
  HS65_LH_BFX4 U9324 ( .A(n8525), .Z(n8524) );
  HS65_LH_BFX4 U9325 ( .A(n8526), .Z(n8525) );
  HS65_LH_BFX4 U9326 ( .A(n8527), .Z(n8526) );
  HS65_LH_BFX4 U9327 ( .A(n8528), .Z(n8527) );
  HS65_LH_BFX4 U9328 ( .A(n8529), .Z(n8528) );
  HS65_LH_BFX4 U9329 ( .A(n8530), .Z(n8529) );
  HS65_LH_BFX4 U9330 ( .A(n14148), .Z(n8530) );
  HS65_LH_BFX4 U9331 ( .A(n8532), .Z(n8531) );
  HS65_LH_BFX4 U9332 ( .A(n8533), .Z(n8532) );
  HS65_LH_BFX4 U9333 ( .A(n8534), .Z(n8533) );
  HS65_LH_BFX4 U9334 ( .A(n8535), .Z(n8534) );
  HS65_LH_BFX4 U9335 ( .A(n8536), .Z(n8535) );
  HS65_LH_BFX4 U9336 ( .A(n8537), .Z(n8536) );
  HS65_LH_BFX4 U9337 ( .A(n8538), .Z(n8537) );
  HS65_LH_BFX4 U9338 ( .A(n8539), .Z(n8538) );
  HS65_LH_BFX4 U9339 ( .A(n8540), .Z(n8539) );
  HS65_LH_BFX4 U9340 ( .A(n8541), .Z(n8540) );
  HS65_LH_BFX4 U9341 ( .A(n8542), .Z(n8541) );
  HS65_LH_BFX4 U9342 ( .A(n8543), .Z(n8542) );
  HS65_LH_BFX4 U9343 ( .A(n8544), .Z(n8543) );
  HS65_LH_BFX4 U9344 ( .A(n8545), .Z(n8544) );
  HS65_LH_BFX4 U9345 ( .A(n8546), .Z(n8545) );
  HS65_LH_BFX4 U9346 ( .A(n8547), .Z(n8546) );
  HS65_LH_BFX4 U9347 ( .A(n8548), .Z(n8547) );
  HS65_LH_BFX4 U9348 ( .A(n8549), .Z(n8548) );
  HS65_LH_BFX4 U9349 ( .A(n8550), .Z(n8549) );
  HS65_LH_BFX4 U9350 ( .A(n8551), .Z(n8550) );
  HS65_LH_BFX4 U9351 ( .A(n8552), .Z(n8551) );
  HS65_LH_BFX4 U9352 ( .A(n8553), .Z(n8552) );
  HS65_LH_BFX4 U9353 ( .A(n8554), .Z(n8553) );
  HS65_LH_BFX4 U9354 ( .A(n8555), .Z(n8554) );
  HS65_LH_BFX4 U9355 ( .A(n14990), .Z(n8555) );
  HS65_LH_BFX4 U9358 ( .A(n8561), .Z(n8558) );
  HS65_LH_BFX4 U9361 ( .A(n8564), .Z(n8561) );
  HS65_LH_BFX4 U9364 ( .A(n8567), .Z(n8564) );
  HS65_LH_BFX4 U9367 ( .A(n8570), .Z(n8567) );
  HS65_LH_BFX4 U9370 ( .A(n8573), .Z(n8570) );
  HS65_LH_BFX4 U9373 ( .A(n8576), .Z(n8573) );
  HS65_LH_BFX4 U9376 ( .A(n8579), .Z(n8576) );
  HS65_LH_BFX4 U9379 ( .A(n8582), .Z(n8579) );
  HS65_LH_BFX4 U9382 ( .A(n8585), .Z(n8582) );
  HS65_LH_BFX4 U9385 ( .A(n8588), .Z(n8585) );
  HS65_LH_BFX4 U9388 ( .A(n8591), .Z(n8588) );
  HS65_LH_BFX4 U9391 ( .A(n8594), .Z(n8591) );
  HS65_LH_BFX4 U9394 ( .A(n8597), .Z(n8594) );
  HS65_LH_BFX4 U9397 ( .A(n8600), .Z(n8597) );
  HS65_LH_BFX4 U9400 ( .A(n8603), .Z(n8600) );
  HS65_LH_BFX4 U9403 ( .A(n8606), .Z(n8603) );
  HS65_LH_BFX4 U9406 ( .A(n8609), .Z(n8606) );
  HS65_LH_BFX4 U9409 ( .A(n8611), .Z(n8609) );
  HS65_LH_BFX4 U9411 ( .A(n8613), .Z(n8611) );
  HS65_LH_BFX4 U9412 ( .A(n8614), .Z(n8612) );
  HS65_LH_BFX4 U9413 ( .A(n8615), .Z(n8613) );
  HS65_LH_BFX4 U9414 ( .A(n15016), .Z(n8614) );
  HS65_LH_BFX4 U9415 ( .A(n8616), .Z(n8615) );
  HS65_LH_BFX4 U9416 ( .A(n8617), .Z(n8616) );
  HS65_LH_BFX4 U9417 ( .A(n8618), .Z(n8617) );
  HS65_LH_BFX4 U9418 ( .A(\u_DataPath/u_idexreg/N25 ), .Z(n8618) );
  HS65_LH_BFX4 U9419 ( .A(n8620), .Z(n8619) );
  HS65_LH_BFX4 U9420 ( .A(n8621), .Z(n8620) );
  HS65_LH_BFX4 U9421 ( .A(n8622), .Z(n8621) );
  HS65_LH_BFX4 U9422 ( .A(n8623), .Z(n8622) );
  HS65_LH_BFX4 U9423 ( .A(n8624), .Z(n8623) );
  HS65_LH_BFX4 U9424 ( .A(n8625), .Z(n8624) );
  HS65_LH_BFX4 U9425 ( .A(n8626), .Z(n8625) );
  HS65_LH_BFX4 U9426 ( .A(n8627), .Z(n8626) );
  HS65_LH_BFX4 U9427 ( .A(n8628), .Z(n8627) );
  HS65_LH_BFX4 U9428 ( .A(n8629), .Z(n8628) );
  HS65_LH_BFX4 U9429 ( .A(n8630), .Z(n8629) );
  HS65_LH_BFX4 U9430 ( .A(n8631), .Z(n8630) );
  HS65_LH_BFX4 U9431 ( .A(n8632), .Z(n8631) );
  HS65_LH_BFX4 U9432 ( .A(n8633), .Z(n8632) );
  HS65_LH_BFX4 U9433 ( .A(n8634), .Z(n8633) );
  HS65_LH_BFX4 U9434 ( .A(n8635), .Z(n8634) );
  HS65_LH_BFX4 U9435 ( .A(n8636), .Z(n8635) );
  HS65_LH_BFX4 U9436 ( .A(n8637), .Z(n8636) );
  HS65_LH_BFX4 U9437 ( .A(n8638), .Z(n8637) );
  HS65_LH_BFX4 U9438 ( .A(n14145), .Z(n8638) );
  HS65_LH_BFX4 U9441 ( .A(n8642), .Z(n8641) );
  HS65_LH_BFX4 U9442 ( .A(n8643), .Z(n8642) );
  HS65_LH_BFX4 U9443 ( .A(n8644), .Z(n8643) );
  HS65_LH_BFX4 U9444 ( .A(n8645), .Z(n8644) );
  HS65_LH_BFX4 U9445 ( .A(n8646), .Z(n8645) );
  HS65_LH_BFX4 U9446 ( .A(n8647), .Z(n8646) );
  HS65_LH_BFX4 U9447 ( .A(n8648), .Z(n8647) );
  HS65_LH_BFX4 U9448 ( .A(n8649), .Z(n8648) );
  HS65_LH_BFX4 U9449 ( .A(n8650), .Z(n8649) );
  HS65_LH_BFX4 U9450 ( .A(n8651), .Z(n8650) );
  HS65_LH_BFX4 U9451 ( .A(n8652), .Z(n8651) );
  HS65_LH_BFX4 U9452 ( .A(n8653), .Z(n8652) );
  HS65_LH_BFX4 U9453 ( .A(n8654), .Z(n8653) );
  HS65_LH_BFX4 U9454 ( .A(n8655), .Z(n8654) );
  HS65_LH_BFX4 U9455 ( .A(n8656), .Z(n8655) );
  HS65_LH_BFX4 U9456 ( .A(n8657), .Z(n8656) );
  HS65_LH_BFX4 U9457 ( .A(n8658), .Z(n8657) );
  HS65_LH_BFX4 U9458 ( .A(n8659), .Z(n8658) );
  HS65_LH_BFX4 U9459 ( .A(n8660), .Z(n8659) );
  HS65_LH_BFX4 U9460 ( .A(n8661), .Z(n8660) );
  HS65_LH_BFX4 U9461 ( .A(n8662), .Z(n8661) );
  HS65_LH_BFX4 U9462 ( .A(n8663), .Z(n8662) );
  HS65_LH_BFX4 U9463 ( .A(n15017), .Z(n8663) );
  HS65_LH_BFX4 U9465 ( .A(n8668), .Z(n8665) );
  HS65_LH_BFX4 U9468 ( .A(n8671), .Z(n8668) );
  HS65_LH_BFX4 U9471 ( .A(n8674), .Z(n8671) );
  HS65_LH_BFX4 U9474 ( .A(n8677), .Z(n8674) );
  HS65_LH_BFX4 U9477 ( .A(n8680), .Z(n8677) );
  HS65_LH_BFX4 U9480 ( .A(n8683), .Z(n8680) );
  HS65_LH_BFX4 U9483 ( .A(n8686), .Z(n8683) );
  HS65_LH_BFX4 U9486 ( .A(n8689), .Z(n8686) );
  HS65_LH_BFX4 U9489 ( .A(n8692), .Z(n8689) );
  HS65_LH_BFX4 U9492 ( .A(n8695), .Z(n8692) );
  HS65_LH_BFX4 U9495 ( .A(n8698), .Z(n8695) );
  HS65_LH_BFX4 U9498 ( .A(n8701), .Z(n8698) );
  HS65_LH_BFX4 U9501 ( .A(n8704), .Z(n8701) );
  HS65_LH_BFX4 U9504 ( .A(n8707), .Z(n8704) );
  HS65_LH_BFX4 U9507 ( .A(n8710), .Z(n8707) );
  HS65_LH_BFX4 U9510 ( .A(n8713), .Z(n8710) );
  HS65_LH_BFX4 U9513 ( .A(n8715), .Z(n8713) );
  HS65_LH_BFX4 U9515 ( .A(n8717), .Z(n8715) );
  HS65_LH_BFX4 U9517 ( .A(n8719), .Z(n8717) );
  HS65_LH_BFX4 U9519 ( .A(n8721), .Z(n8719) );
  HS65_LH_BFX4 U9521 ( .A(n8723), .Z(n8721) );
  HS65_LH_BFX4 U9523 ( .A(n8724), .Z(n8723) );
  HS65_LH_BFX4 U9524 ( .A(n8725), .Z(n8724) );
  HS65_LH_BFX4 U9525 ( .A(n8726), .Z(n8725) );
  HS65_LH_BFX4 U9526 ( .A(\u_DataPath/u_idexreg/N26 ), .Z(n8726) );
  HS65_LH_BFX4 U9556 ( .A(n8758), .Z(n8756) );
  HS65_LH_BFX4 U9558 ( .A(n8760), .Z(n8758) );
  HS65_LH_BFX4 U9560 ( .A(n8762), .Z(n8760) );
  HS65_LH_BFX4 U9562 ( .A(n8764), .Z(n8762) );
  HS65_LH_BFX4 U9564 ( .A(n8766), .Z(n8764) );
  HS65_LH_BFX4 U9566 ( .A(n8768), .Z(n8766) );
  HS65_LH_BFX4 U9568 ( .A(n8770), .Z(n8768) );
  HS65_LH_BFX4 U9570 ( .A(n8772), .Z(n8770) );
  HS65_LH_BFX4 U9572 ( .A(n8774), .Z(n8772) );
  HS65_LH_BFX4 U9574 ( .A(n8776), .Z(n8774) );
  HS65_LH_BFX4 U9576 ( .A(n8778), .Z(n8776) );
  HS65_LH_BFX4 U9578 ( .A(n8780), .Z(n8778) );
  HS65_LH_BFX4 U9580 ( .A(n8782), .Z(n8780) );
  HS65_LH_BFX4 U9582 ( .A(n8784), .Z(n8782) );
  HS65_LH_BFX4 U9584 ( .A(n8786), .Z(n8784) );
  HS65_LH_BFX4 U9586 ( .A(n8788), .Z(n8786) );
  HS65_LH_BFX4 U9588 ( .A(n8789), .Z(n8788) );
  HS65_LH_BFX4 U9589 ( .A(n8790), .Z(n8789) );
  HS65_LH_BFX4 U9590 ( .A(n8791), .Z(n8790) );
  HS65_LH_BFX4 U9591 ( .A(n15056), .Z(n8791) );
  HS65_LH_BFX4 U9592 ( .A(n8793), .Z(n8792) );
  HS65_LH_BFX4 U9593 ( .A(n8794), .Z(n8793) );
  HS65_LH_BFX4 U9594 ( .A(n8795), .Z(n8794) );
  HS65_LH_BFX4 U9595 ( .A(n8796), .Z(n8795) );
  HS65_LH_BFX4 U9596 ( .A(n8797), .Z(n8796) );
  HS65_LH_BFX4 U9597 ( .A(n8798), .Z(n8797) );
  HS65_LH_BFX4 U9598 ( .A(n8799), .Z(n8798) );
  HS65_LH_BFX4 U9599 ( .A(n8800), .Z(n8799) );
  HS65_LH_BFX4 U9600 ( .A(n8801), .Z(n8800) );
  HS65_LH_BFX4 U9601 ( .A(n8802), .Z(n8801) );
  HS65_LH_BFX4 U9602 ( .A(n8803), .Z(n8802) );
  HS65_LH_BFX4 U9603 ( .A(n8804), .Z(n8803) );
  HS65_LH_BFX4 U9604 ( .A(n8805), .Z(n8804) );
  HS65_LH_BFX4 U9605 ( .A(n8806), .Z(n8805) );
  HS65_LH_BFX4 U9606 ( .A(n8807), .Z(n8806) );
  HS65_LH_BFX4 U9607 ( .A(n8808), .Z(n8807) );
  HS65_LH_BFX4 U9608 ( .A(n8809), .Z(n8808) );
  HS65_LH_BFX4 U9609 ( .A(n8810), .Z(n8809) );
  HS65_LH_BFX4 U9610 ( .A(n8811), .Z(n8810) );
  HS65_LH_BFX4 U9611 ( .A(n14221), .Z(n8811) );
  HS65_LH_BFX4 U9612 ( .A(n8813), .Z(n8812) );
  HS65_LH_BFX4 U9613 ( .A(n8814), .Z(n8813) );
  HS65_LH_BFX4 U9614 ( .A(n8815), .Z(n8814) );
  HS65_LH_BFX4 U9615 ( .A(n8816), .Z(n8815) );
  HS65_LH_BFX4 U9616 ( .A(n8817), .Z(n8816) );
  HS65_LH_BFX4 U9617 ( .A(n8818), .Z(n8817) );
  HS65_LH_BFX4 U9618 ( .A(n8819), .Z(n8818) );
  HS65_LH_BFX4 U9619 ( .A(n8820), .Z(n8819) );
  HS65_LH_BFX4 U9620 ( .A(n8821), .Z(n8820) );
  HS65_LH_BFX4 U9621 ( .A(n8822), .Z(n8821) );
  HS65_LH_BFX4 U9622 ( .A(n8823), .Z(n8822) );
  HS65_LH_BFX4 U9623 ( .A(n8824), .Z(n8823) );
  HS65_LH_BFX4 U9624 ( .A(n8825), .Z(n8824) );
  HS65_LH_BFX4 U9625 ( .A(n8826), .Z(n8825) );
  HS65_LH_BFX4 U9626 ( .A(n8827), .Z(n8826) );
  HS65_LH_BFX4 U9627 ( .A(n8828), .Z(n8827) );
  HS65_LH_BFX4 U9628 ( .A(n8829), .Z(n8828) );
  HS65_LH_BFX4 U9629 ( .A(n8830), .Z(n8829) );
  HS65_LH_BFX4 U9630 ( .A(n8831), .Z(n8830) );
  HS65_LH_BFX4 U9631 ( .A(n8832), .Z(n8831) );
  HS65_LH_BFX4 U9632 ( .A(n8833), .Z(n8832) );
  HS65_LH_BFX4 U9633 ( .A(n8834), .Z(n8833) );
  HS65_LH_BFX4 U9634 ( .A(n8835), .Z(n8834) );
  HS65_LH_BFX4 U9635 ( .A(n8836), .Z(n8835) );
  HS65_LH_BFX4 U9636 ( .A(n15699), .Z(n8836) );
  HS65_LH_BFX4 U9637 ( .A(n10755), .Z(n8837) );
  HS65_LH_BFX4 U9638 ( .A(n8855), .Z(n8838) );
  HS65_LH_BFX4 U9640 ( .A(\u_DataPath/pc_4_to_ex_i [2]), .Z(n8840) );
  HS65_LH_BFX4 U9642 ( .A(n8840), .Z(n8842) );
  HS65_LH_BFX4 U9644 ( .A(n8842), .Z(n8844) );
  HS65_LH_BFX4 U9646 ( .A(n8844), .Z(n8846) );
  HS65_LH_BFX4 U9648 ( .A(n8846), .Z(n8848) );
  HS65_LH_BFX4 U9650 ( .A(n8848), .Z(n8850) );
  HS65_LH_BFX4 U9652 ( .A(n8850), .Z(n8852) );
  HS65_LH_CNIVX3 U9654 ( .A(n8858), .Z(n8854) );
  HS65_LH_CNIVX3 U9655 ( .A(n8854), .Z(n8855) );
  HS65_LH_BFX4 U9658 ( .A(n8862), .Z(n8858) );
  HS65_LH_CNIVX3 U9659 ( .A(n8875), .Z(n8859) );
  HS65_LH_CNIVX3 U9660 ( .A(n8859), .Z(n8860) );
  HS65_LH_BFX4 U9662 ( .A(n8864), .Z(n8862) );
  HS65_LH_BFX4 U9664 ( .A(n8866), .Z(n8864) );
  HS65_LH_BFX4 U9666 ( .A(n8868), .Z(n8866) );
  HS65_LH_BFX4 U9668 ( .A(n8870), .Z(n8868) );
  HS65_LH_BFX4 U9670 ( .A(n8872), .Z(n8870) );
  HS65_LH_BFX4 U9672 ( .A(n8874), .Z(n8872) );
  HS65_LH_BFX4 U9674 ( .A(n14110), .Z(n8874) );
  HS65_LH_BFX4 U9675 ( .A(n8876), .Z(n8875) );
  HS65_LH_BFX4 U9676 ( .A(n8877), .Z(n8876) );
  HS65_LH_BFX4 U9677 ( .A(n8852), .Z(n8877) );
  HS65_LH_BFX4 U9678 ( .A(n8879), .Z(n8878) );
  HS65_LH_BFX4 U9679 ( .A(n8880), .Z(n8879) );
  HS65_LH_BFX4 U9680 ( .A(n8881), .Z(n8880) );
  HS65_LH_BFX4 U9681 ( .A(n8882), .Z(n8881) );
  HS65_LH_BFX4 U9682 ( .A(n8883), .Z(n8882) );
  HS65_LH_BFX4 U9683 ( .A(n8884), .Z(n8883) );
  HS65_LH_BFX4 U9684 ( .A(n8885), .Z(n8884) );
  HS65_LH_BFX4 U9685 ( .A(n8886), .Z(n8885) );
  HS65_LH_BFX4 U9686 ( .A(n8887), .Z(n8886) );
  HS65_LH_BFX4 U9687 ( .A(n8888), .Z(n8887) );
  HS65_LH_BFX4 U9688 ( .A(n8889), .Z(n8888) );
  HS65_LH_BFX4 U9689 ( .A(n8890), .Z(n8889) );
  HS65_LH_BFX4 U9690 ( .A(n8891), .Z(n8890) );
  HS65_LH_BFX4 U9691 ( .A(n8892), .Z(n8891) );
  HS65_LH_BFX4 U9692 ( .A(n8893), .Z(n8892) );
  HS65_LH_BFX4 U9693 ( .A(n8894), .Z(n8893) );
  HS65_LH_BFX4 U9694 ( .A(n8895), .Z(n8894) );
  HS65_LH_BFX4 U9695 ( .A(n8896), .Z(n8895) );
  HS65_LH_BFX4 U9696 ( .A(n8897), .Z(n8896) );
  HS65_LH_BFX4 U9697 ( .A(n14113), .Z(n8897) );
  HS65_LH_BFX4 U9706 ( .A(n8907), .Z(n8906) );
  HS65_LH_BFX4 U9707 ( .A(n8908), .Z(n8907) );
  HS65_LH_BFX4 U9708 ( .A(n8909), .Z(n8908) );
  HS65_LH_BFX4 U9709 ( .A(n8910), .Z(n8909) );
  HS65_LH_BFX4 U9710 ( .A(n8911), .Z(n8910) );
  HS65_LH_BFX4 U9711 ( .A(n8912), .Z(n8911) );
  HS65_LH_BFX4 U9712 ( .A(n8913), .Z(n8912) );
  HS65_LH_BFX4 U9713 ( .A(n8914), .Z(n8913) );
  HS65_LH_BFX4 U9714 ( .A(n8915), .Z(n8914) );
  HS65_LH_BFX4 U9715 ( .A(n8916), .Z(n8915) );
  HS65_LH_BFX4 U9716 ( .A(n8917), .Z(n8916) );
  HS65_LH_BFX4 U9717 ( .A(n8918), .Z(n8917) );
  HS65_LH_BFX4 U9718 ( .A(n8919), .Z(n8918) );
  HS65_LH_BFX4 U9719 ( .A(n8920), .Z(n8919) );
  HS65_LH_BFX4 U9720 ( .A(n8921), .Z(n8920) );
  HS65_LH_BFX4 U9721 ( .A(n8922), .Z(n8921) );
  HS65_LH_BFX4 U9722 ( .A(n15094), .Z(n8922) );
  HS65_LH_CNIVX3 U9723 ( .A(\u_DataPath/pc_4_to_ex_i [18]), .Z(n8923) );
  HS65_LH_CNIVX3 U9724 ( .A(n8923), .Z(n8924) );
  HS65_LH_BFX4 U9726 ( .A(n8928), .Z(n8926) );
  HS65_LH_BFX4 U9728 ( .A(n8931), .Z(n8928) );
  HS65_LH_BFX4 U9731 ( .A(n8934), .Z(n8931) );
  HS65_LH_BFX4 U9734 ( .A(n8936), .Z(n8934) );
  HS65_LH_BFX4 U9736 ( .A(n8939), .Z(n8936) );
  HS65_LH_BFX4 U9739 ( .A(n8942), .Z(n8939) );
  HS65_LH_BFX4 U9742 ( .A(n8945), .Z(n8942) );
  HS65_LH_BFX4 U9745 ( .A(n8948), .Z(n8945) );
  HS65_LH_BFX4 U9748 ( .A(n8951), .Z(n8948) );
  HS65_LH_BFX4 U9751 ( .A(n8954), .Z(n8951) );
  HS65_LH_BFX4 U9754 ( .A(n8957), .Z(n8954) );
  HS65_LH_BFX4 U9757 ( .A(n8960), .Z(n8957) );
  HS65_LH_BFX4 U9760 ( .A(n8963), .Z(n8960) );
  HS65_LH_BFX4 U9763 ( .A(n8966), .Z(n8963) );
  HS65_LH_BFX4 U9766 ( .A(n8969), .Z(n8966) );
  HS65_LH_BFX4 U9769 ( .A(n8972), .Z(n8969) );
  HS65_LH_BFX4 U9772 ( .A(n8975), .Z(n8972) );
  HS65_LH_BFX4 U9775 ( .A(n8978), .Z(n8975) );
  HS65_LH_BFX4 U9778 ( .A(n8980), .Z(n8978) );
  HS65_LH_BFX4 U9780 ( .A(n8982), .Z(n8980) );
  HS65_LH_BFX4 U9782 ( .A(n8984), .Z(n8982) );
  HS65_LH_BFX4 U9784 ( .A(n8985), .Z(n8984) );
  HS65_LH_BFX4 U9785 ( .A(n8986), .Z(n8985) );
  HS65_LH_BFX4 U9786 ( .A(n8987), .Z(n8986) );
  HS65_LH_BFX4 U9787 ( .A(\u_DataPath/u_idexreg/N27 ), .Z(n8987) );
  HS65_LH_BFX4 U9788 ( .A(n8989), .Z(n8988) );
  HS65_LH_BFX4 U9789 ( .A(n8990), .Z(n8989) );
  HS65_LH_BFX4 U9790 ( .A(n8991), .Z(n8990) );
  HS65_LH_BFX4 U9791 ( .A(n8992), .Z(n8991) );
  HS65_LH_BFX4 U9792 ( .A(n8993), .Z(n8992) );
  HS65_LH_BFX4 U9793 ( .A(n8994), .Z(n8993) );
  HS65_LH_BFX4 U9794 ( .A(n8995), .Z(n8994) );
  HS65_LH_BFX4 U9795 ( .A(n8996), .Z(n8995) );
  HS65_LH_BFX4 U9796 ( .A(n8997), .Z(n8996) );
  HS65_LH_BFX4 U9797 ( .A(n8998), .Z(n8997) );
  HS65_LH_BFX4 U9798 ( .A(n8999), .Z(n8998) );
  HS65_LH_BFX4 U9799 ( .A(n9000), .Z(n8999) );
  HS65_LH_BFX4 U9800 ( .A(n9001), .Z(n9000) );
  HS65_LH_BFX4 U9801 ( .A(n9002), .Z(n9001) );
  HS65_LH_BFX4 U9802 ( .A(n9003), .Z(n9002) );
  HS65_LH_BFX4 U9803 ( .A(n9004), .Z(n9003) );
  HS65_LH_BFX4 U9804 ( .A(n9005), .Z(n9004) );
  HS65_LH_BFX4 U9805 ( .A(n9006), .Z(n9005) );
  HS65_LH_BFX4 U9806 ( .A(n9007), .Z(n9006) );
  HS65_LH_BFX4 U9807 ( .A(n9008), .Z(n9007) );
  HS65_LH_BFX4 U9808 ( .A(n9009), .Z(n9008) );
  HS65_LH_BFX4 U9809 ( .A(n9010), .Z(n9009) );
  HS65_LH_BFX4 U9810 ( .A(n9011), .Z(n9010) );
  HS65_LH_BFX4 U9811 ( .A(n9012), .Z(n9011) );
  HS65_LH_BFX4 U9812 ( .A(n15652), .Z(n9012) );
  HS65_LH_BFX4 U9814 ( .A(n9016), .Z(n9014) );
  HS65_LH_BFX4 U9816 ( .A(n9017), .Z(n9016) );
  HS65_LH_BFX4 U9817 ( .A(n9024), .Z(n9017) );
  HS65_LH_CNIVX3 U9819 ( .A(n9022), .Z(n9019) );
  HS65_LH_CNIVX3 U9820 ( .A(n9019), .Z(n9020) );
  HS65_LH_BFX4 U9822 ( .A(\u_DataPath/pc_4_to_ex_i [6]), .Z(n9022) );
  HS65_LH_BFX4 U9824 ( .A(n9026), .Z(n9024) );
  HS65_LH_BFX4 U9826 ( .A(n9028), .Z(n9026) );
  HS65_LH_BFX4 U9828 ( .A(n9030), .Z(n9028) );
  HS65_LH_BFX4 U9830 ( .A(n9032), .Z(n9030) );
  HS65_LH_BFX4 U9832 ( .A(n9034), .Z(n9032) );
  HS65_LH_BFX4 U9834 ( .A(n9036), .Z(n9034) );
  HS65_LH_BFX4 U9836 ( .A(n9038), .Z(n9036) );
  HS65_LH_BFX4 U9838 ( .A(n9040), .Z(n9038) );
  HS65_LH_BFX4 U9840 ( .A(n9042), .Z(n9040) );
  HS65_LH_BFX4 U9842 ( .A(n9044), .Z(n9042) );
  HS65_LH_BFX4 U9844 ( .A(n9046), .Z(n9044) );
  HS65_LH_BFX4 U9846 ( .A(n9048), .Z(n9046) );
  HS65_LH_BFX4 U9848 ( .A(n9050), .Z(n9048) );
  HS65_LH_BFX4 U9850 ( .A(n9051), .Z(n9050) );
  HS65_LH_BFX4 U9851 ( .A(n9052), .Z(n9051) );
  HS65_LH_BFX4 U9852 ( .A(n15161), .Z(n9052) );
  HS65_LH_BFX4 U9877 ( .A(n9078), .Z(n9077) );
  HS65_LH_BFX4 U9878 ( .A(n9079), .Z(n9078) );
  HS65_LH_BFX4 U9879 ( .A(n9080), .Z(n9079) );
  HS65_LH_BFX4 U9880 ( .A(n9081), .Z(n9080) );
  HS65_LH_BFX4 U9881 ( .A(n9082), .Z(n9081) );
  HS65_LH_BFX4 U9882 ( .A(n9083), .Z(n9082) );
  HS65_LH_BFX4 U9883 ( .A(n9084), .Z(n9083) );
  HS65_LH_BFX4 U9884 ( .A(n9085), .Z(n9084) );
  HS65_LH_BFX4 U9885 ( .A(n9086), .Z(n9085) );
  HS65_LH_BFX4 U9886 ( .A(n9087), .Z(n9086) );
  HS65_LH_BFX4 U9887 ( .A(n9088), .Z(n9087) );
  HS65_LH_BFX4 U9888 ( .A(n9089), .Z(n9088) );
  HS65_LH_BFX4 U9889 ( .A(n9090), .Z(n9089) );
  HS65_LH_BFX4 U9890 ( .A(n9091), .Z(n9090) );
  HS65_LH_BFX4 U9891 ( .A(n9092), .Z(n9091) );
  HS65_LH_BFX4 U9892 ( .A(n9093), .Z(n9092) );
  HS65_LH_BFX4 U9893 ( .A(n9094), .Z(n9093) );
  HS65_LH_BFX4 U9894 ( .A(n9095), .Z(n9094) );
  HS65_LH_BFX4 U9895 ( .A(n9096), .Z(n9095) );
  HS65_LH_BFX4 U9896 ( .A(n14233), .Z(n9096) );
  HS65_LH_BFX4 U9912 ( .A(n9113), .Z(n9112) );
  HS65_LH_BFX4 U9913 ( .A(n9114), .Z(n9113) );
  HS65_LH_BFX4 U9914 ( .A(n9115), .Z(n9114) );
  HS65_LH_BFX4 U9915 ( .A(n9116), .Z(n9115) );
  HS65_LH_BFX4 U9916 ( .A(n9117), .Z(n9116) );
  HS65_LH_BFX4 U9917 ( .A(n9118), .Z(n9117) );
  HS65_LH_BFX4 U9918 ( .A(n9119), .Z(n9118) );
  HS65_LH_BFX4 U9919 ( .A(n9120), .Z(n9119) );
  HS65_LH_BFX4 U9920 ( .A(\u_DataPath/data_read_ex_2_i [1]), .Z(n9120) );
  HS65_LH_BFX4 U9922 ( .A(n9124), .Z(n9122) );
  HS65_LH_BFX4 U9924 ( .A(n9126), .Z(n9124) );
  HS65_LH_BFX4 U9926 ( .A(n9128), .Z(n9126) );
  HS65_LH_BFX4 U9928 ( .A(n9130), .Z(n9128) );
  HS65_LH_BFX4 U9930 ( .A(n9132), .Z(n9130) );
  HS65_LH_BFX4 U9932 ( .A(n9134), .Z(n9132) );
  HS65_LH_BFX4 U9934 ( .A(n9136), .Z(n9134) );
  HS65_LH_BFX4 U9936 ( .A(n9138), .Z(n9136) );
  HS65_LH_BFX4 U9938 ( .A(n9140), .Z(n9138) );
  HS65_LH_BFX4 U9940 ( .A(n9142), .Z(n9140) );
  HS65_LH_BFX4 U9942 ( .A(n9144), .Z(n9142) );
  HS65_LH_BFX4 U9944 ( .A(n9146), .Z(n9144) );
  HS65_LH_BFX4 U9946 ( .A(n9148), .Z(n9146) );
  HS65_LH_BFX4 U9948 ( .A(n9150), .Z(n9148) );
  HS65_LH_BFX4 U9950 ( .A(n9152), .Z(n9150) );
  HS65_LH_BFX4 U9952 ( .A(n9154), .Z(n9152) );
  HS65_LH_BFX4 U9954 ( .A(n9156), .Z(n9154) );
  HS65_LH_BFX4 U9956 ( .A(n9158), .Z(n9156) );
  HS65_LH_BFX4 U9958 ( .A(n9160), .Z(n9158) );
  HS65_LH_BFX4 U9960 ( .A(n9161), .Z(n9160) );
  HS65_LH_BFX4 U9961 ( .A(n9162), .Z(n9161) );
  HS65_LH_BFX4 U9962 ( .A(n15162), .Z(n9162) );
  HS65_LH_BFX4 U9963 ( .A(n9164), .Z(n9163) );
  HS65_LH_BFX4 U9964 ( .A(n9165), .Z(n9164) );
  HS65_LH_BFX4 U9965 ( .A(n9166), .Z(n9165) );
  HS65_LH_BFX4 U9966 ( .A(n9167), .Z(n9166) );
  HS65_LH_BFX4 U9967 ( .A(n9168), .Z(n9167) );
  HS65_LH_BFX4 U9968 ( .A(n9169), .Z(n9168) );
  HS65_LH_BFX4 U9969 ( .A(n9170), .Z(n9169) );
  HS65_LH_BFX4 U9970 ( .A(n9171), .Z(n9170) );
  HS65_LH_BFX4 U9971 ( .A(n9172), .Z(n9171) );
  HS65_LH_BFX4 U9972 ( .A(n9173), .Z(n9172) );
  HS65_LH_BFX4 U9973 ( .A(n9174), .Z(n9173) );
  HS65_LH_BFX4 U9974 ( .A(n9175), .Z(n9174) );
  HS65_LH_BFX4 U9975 ( .A(n9176), .Z(n9175) );
  HS65_LH_BFX4 U9976 ( .A(n9177), .Z(n9176) );
  HS65_LH_BFX4 U9977 ( .A(n9178), .Z(n9177) );
  HS65_LH_BFX4 U9978 ( .A(n9179), .Z(n9178) );
  HS65_LH_BFX4 U9979 ( .A(n9180), .Z(n9179) );
  HS65_LH_BFX4 U9980 ( .A(n9181), .Z(n9180) );
  HS65_LH_BFX4 U9981 ( .A(n9182), .Z(n9181) );
  HS65_LH_BFX4 U9982 ( .A(n14214), .Z(n9182) );
  HS65_LH_BFX4 U10002 ( .A(n9203), .Z(n9202) );
  HS65_LH_BFX4 U10003 ( .A(n9204), .Z(n9203) );
  HS65_LH_BFX4 U10004 ( .A(n9205), .Z(n9204) );
  HS65_LH_BFX4 U10005 ( .A(n9206), .Z(n9205) );
  HS65_LH_BFX4 U10006 ( .A(\u_DataPath/data_read_ex_2_i [0]), .Z(n9206) );
  HS65_LH_BFX4 U10008 ( .A(n9210), .Z(n9208) );
  HS65_LH_BFX4 U10010 ( .A(n9212), .Z(n9210) );
  HS65_LH_BFX4 U10012 ( .A(n9214), .Z(n9212) );
  HS65_LH_BFX4 U10014 ( .A(n9216), .Z(n9214) );
  HS65_LH_BFX4 U10016 ( .A(n9218), .Z(n9216) );
  HS65_LH_BFX4 U10018 ( .A(n9220), .Z(n9218) );
  HS65_LH_BFX4 U10020 ( .A(n9222), .Z(n9220) );
  HS65_LH_BFX4 U10022 ( .A(n9224), .Z(n9222) );
  HS65_LH_BFX4 U10024 ( .A(n9226), .Z(n9224) );
  HS65_LH_BFX4 U10026 ( .A(n9228), .Z(n9226) );
  HS65_LH_BFX4 U10028 ( .A(n9230), .Z(n9228) );
  HS65_LH_BFX4 U10030 ( .A(n9233), .Z(n9230) );
  HS65_LH_BFX4 U10033 ( .A(n9235), .Z(n9233) );
  HS65_LH_BFX4 U10034 ( .A(n9236), .Z(n9234) );
  HS65_LH_BFX4 U10035 ( .A(n9237), .Z(n9235) );
  HS65_LH_BFX4 U10036 ( .A(n9238), .Z(n9236) );
  HS65_LH_BFX4 U10037 ( .A(n9239), .Z(n9237) );
  HS65_LH_BFX4 U10038 ( .A(n9240), .Z(n9238) );
  HS65_LH_BFX4 U10039 ( .A(n9241), .Z(n9239) );
  HS65_LH_BFX4 U10040 ( .A(n9242), .Z(n9240) );
  HS65_LH_BFX4 U10041 ( .A(n9243), .Z(n9241) );
  HS65_LH_BFX4 U10042 ( .A(n9244), .Z(n9242) );
  HS65_LH_BFX4 U10043 ( .A(n9245), .Z(n9243) );
  HS65_LH_BFX4 U10044 ( .A(n9246), .Z(n9244) );
  HS65_LH_BFX4 U10045 ( .A(n9247), .Z(n9245) );
  HS65_LH_BFX4 U10046 ( .A(n9248), .Z(n9246) );
  HS65_LH_BFX4 U10047 ( .A(n9249), .Z(n9247) );
  HS65_LH_BFX4 U10048 ( .A(\u_DataPath/data_read_ex_1_i [0]), .Z(n9248) );
  HS65_LH_BFX4 U10049 ( .A(n9250), .Z(n9249) );
  HS65_LH_BFX4 U10050 ( .A(n15166), .Z(n9250) );
  HS65_LH_BFX4 U10052 ( .A(n9254), .Z(n9252) );
  HS65_LH_BFX4 U10054 ( .A(n9256), .Z(n9254) );
  HS65_LH_BFX4 U10056 ( .A(n9258), .Z(n9256) );
  HS65_LH_BFX4 U10058 ( .A(n9260), .Z(n9258) );
  HS65_LH_BFX4 U10060 ( .A(n9262), .Z(n9260) );
  HS65_LH_BFX4 U10062 ( .A(n9264), .Z(n9262) );
  HS65_LH_BFX4 U10064 ( .A(n9266), .Z(n9264) );
  HS65_LH_BFX4 U10066 ( .A(n9270), .Z(n9266) );
  HS65_LH_BFX4 U10070 ( .A(n9272), .Z(n9270) );
  HS65_LH_BFX4 U10072 ( .A(n9274), .Z(n9272) );
  HS65_LH_BFX4 U10074 ( .A(n9275), .Z(n9274) );
  HS65_LH_BFX4 U10075 ( .A(n9276), .Z(n9275) );
  HS65_LH_BFX4 U10076 ( .A(n9277), .Z(n9276) );
  HS65_LH_BFX4 U10077 ( .A(n9278), .Z(n9277) );
  HS65_LH_BFX4 U10078 ( .A(n9279), .Z(n9278) );
  HS65_LH_BFX4 U10079 ( .A(n9280), .Z(n9279) );
  HS65_LH_BFX4 U10080 ( .A(n9281), .Z(n9280) );
  HS65_LH_BFX4 U10081 ( .A(n9282), .Z(n9281) );
  HS65_LH_BFX4 U10082 ( .A(n9283), .Z(n9282) );
  HS65_LH_BFX4 U10083 ( .A(n14216), .Z(n9283) );
  HS65_LH_BFX4 U10084 ( .A(n9288), .Z(n9284) );
  HS65_LL_NOR3AX2 U10085 ( .A(n10585), .B(n10589), .C(n14074), .Z(n14075) );
  HS65_LH_BFX4 U10086 ( .A(n9291), .Z(n9285) );
  HS65_LH_BFX4 U10087 ( .A(n9305), .Z(n9286) );
  HS65_LH_BFX4 U10088 ( .A(n14069), .Z(n9287) );
  HS65_LH_BFX4 U10089 ( .A(n9294), .Z(n9288) );
  HS65_LH_BFX4 U10090 ( .A(n10575), .Z(n9289) );
  HS65_LH_BFX4 U10091 ( .A(n10573), .Z(n9290) );
  HS65_LH_BFX4 U10092 ( .A(n9295), .Z(n9291) );
  HS65_LH_BFX4 U10093 ( .A(n9296), .Z(n9292) );
  HS65_LH_BFX4 U10094 ( .A(n9287), .Z(n9293) );
  HS65_LH_BFX4 U10095 ( .A(n9298), .Z(n9294) );
  HS65_LH_BFX4 U10096 ( .A(n9299), .Z(n9295) );
  HS65_LH_BFX4 U10097 ( .A(n9310), .Z(n9296) );
  HS65_LH_BFX4 U10098 ( .A(n15701), .Z(n9297) );
  HS65_LH_BFX4 U10099 ( .A(n9301), .Z(n9298) );
  HS65_LH_BFX4 U10100 ( .A(n9302), .Z(n9299) );
  HS65_LH_BFX4 U10101 ( .A(n9297), .Z(n9300) );
  HS65_LH_BFX4 U10102 ( .A(n10560), .Z(n9301) );
  HS65_LH_BFX4 U10103 ( .A(n9304), .Z(n9302) );
  HS65_LH_BFX4 U10104 ( .A(n9300), .Z(n9303) );
  HS65_LH_BFX4 U10105 ( .A(n10676), .Z(n9304) );
  HS65_LH_NAND3X2 U10106 ( .A(n14076), .B(n10710), .C(n14068), .Z(n15701) );
  HS65_LH_BFX4 U10107 ( .A(n9303), .Z(n9305) );
  HS65_LH_BFX4 U10108 ( .A(\u_DataPath/cw_tomem_i [4]), .Z(n9306) );
  HS65_LH_BFX4 U10109 ( .A(n9308), .Z(n9307) );
  HS65_LH_BFX4 U10110 ( .A(n9309), .Z(n9308) );
  HS65_LH_BFX4 U10111 ( .A(n288), .Z(n9309) );
  HS65_LH_BFX4 U10112 ( .A(n9311), .Z(n9310) );
  HS65_LH_BFX4 U10113 ( .A(n9312), .Z(n9311) );
  HS65_LH_BFX4 U10114 ( .A(n9313), .Z(n9312) );
  HS65_LH_BFX4 U10115 ( .A(n10554), .Z(n9313) );
  HS65_LH_BFX4 U10116 ( .A(n9316), .Z(n9314) );
  HS65_LH_BFX4 U10117 ( .A(\u_DataPath/dataOut_exe_i [0]), .Z(n9315) );
  HS65_LH_BFX4 U10118 ( .A(n14070), .Z(n9316) );
  HS65_LH_BFX4 U10119 ( .A(n9315), .Z(n9317) );
  HS65_LH_BFX4 U10120 ( .A(n9317), .Z(n9318) );
  HS65_LH_BFX4 U10121 ( .A(n9322), .Z(n9319) );
  HS65_LH_BFX4 U10122 ( .A(\u_DataPath/u_execute/link_value_i [0]), .Z(n9320)
         );
  HS65_LH_BFX4 U10124 ( .A(n9325), .Z(n9322) );
  HS65_LH_BFX4 U10125 ( .A(n9320), .Z(n9323) );
  HS65_LH_BFX4 U10127 ( .A(n9328), .Z(n9325) );
  HS65_LH_BFX4 U10128 ( .A(n9323), .Z(n9326) );
  HS65_LH_BFX4 U10130 ( .A(n9331), .Z(n9328) );
  HS65_LH_BFX4 U10131 ( .A(n9326), .Z(n9329) );
  HS65_LH_BFX4 U10133 ( .A(n9334), .Z(n9331) );
  HS65_LH_BFX4 U10134 ( .A(n9329), .Z(n9332) );
  HS65_LH_BFX4 U10136 ( .A(n9337), .Z(n9334) );
  HS65_LH_BFX4 U10137 ( .A(n9332), .Z(n9335) );
  HS65_LH_BFX4 U10139 ( .A(n9340), .Z(n9337) );
  HS65_LH_BFX4 U10140 ( .A(n9335), .Z(n9338) );
  HS65_LH_BFX4 U10142 ( .A(n9343), .Z(n9340) );
  HS65_LH_BFX4 U10143 ( .A(n9338), .Z(n9341) );
  HS65_LH_BFX4 U10145 ( .A(n9346), .Z(n9343) );
  HS65_LH_BFX4 U10146 ( .A(n9341), .Z(n9344) );
  HS65_LH_BFX4 U10148 ( .A(n9349), .Z(n9346) );
  HS65_LH_BFX4 U10149 ( .A(n9344), .Z(n9347) );
  HS65_LH_BFX4 U10151 ( .A(n9352), .Z(n9349) );
  HS65_LH_BFX4 U10152 ( .A(n9347), .Z(n9350) );
  HS65_LH_BFX4 U10154 ( .A(n9355), .Z(n9352) );
  HS65_LH_BFX4 U10155 ( .A(n9350), .Z(n9353) );
  HS65_LH_BFX4 U10157 ( .A(n9358), .Z(n9355) );
  HS65_LH_BFX4 U10158 ( .A(n9353), .Z(n9356) );
  HS65_LH_BFX4 U10160 ( .A(n9361), .Z(n9358) );
  HS65_LH_BFX4 U10161 ( .A(n9356), .Z(n9359) );
  HS65_LH_BFX4 U10163 ( .A(n9364), .Z(n9361) );
  HS65_LH_BFX4 U10164 ( .A(n9359), .Z(n9362) );
  HS65_LH_BFX4 U10166 ( .A(n9367), .Z(n9364) );
  HS65_LH_BFX4 U10167 ( .A(n9362), .Z(n9365) );
  HS65_LH_BFX4 U10169 ( .A(n9370), .Z(n9367) );
  HS65_LH_BFX4 U10170 ( .A(n9365), .Z(n9368) );
  HS65_LH_BFX4 U10172 ( .A(n9375), .Z(n9370) );
  HS65_LH_BFX4 U10173 ( .A(n9368), .Z(n9371) );
  HS65_LH_CNIVX3 U10175 ( .A(n9382), .Z(n9373) );
  HS65_LH_CNIVX3 U10176 ( .A(n9373), .Z(n9374) );
  HS65_LH_BFX4 U10177 ( .A(n9380), .Z(n9375) );
  HS65_LH_BFX4 U10179 ( .A(n9371), .Z(n9377) );
  HS65_LH_BFX4 U10182 ( .A(n9381), .Z(n9380) );
  HS65_LH_BFX4 U10183 ( .A(n9383), .Z(n9381) );
  HS65_LH_BFX4 U10184 ( .A(n9385), .Z(n9382) );
  HS65_LH_BFX4 U10185 ( .A(n9384), .Z(n9383) );
  HS65_LH_BFX4 U10186 ( .A(n9386), .Z(n9384) );
  HS65_LH_BFX4 U10187 ( .A(n9387), .Z(n9385) );
  HS65_LH_BFX4 U10188 ( .A(n9388), .Z(n9386) );
  HS65_LH_BFX4 U10189 ( .A(n9389), .Z(n9387) );
  HS65_LH_BFX4 U10190 ( .A(\u_DataPath/u_execute/psw_status_i [0]), .Z(n9388)
         );
  HS65_LH_BFX4 U10191 ( .A(n9377), .Z(n9389) );
  HS65_LH_BFX4 U10219 ( .A(n9420), .Z(n9417) );
  HS65_LH_BFX4 U10222 ( .A(n9423), .Z(n9420) );
  HS65_LH_BFX4 U10225 ( .A(n9426), .Z(n9423) );
  HS65_LH_BFX4 U10228 ( .A(n9429), .Z(n9426) );
  HS65_LH_BFX4 U10231 ( .A(n9432), .Z(n9429) );
  HS65_LH_BFX4 U10234 ( .A(n9435), .Z(n9432) );
  HS65_LH_BFX4 U10237 ( .A(n9438), .Z(n9435) );
  HS65_LH_BFX4 U10240 ( .A(n9441), .Z(n9438) );
  HS65_LH_BFX4 U10243 ( .A(n9444), .Z(n9441) );
  HS65_LH_BFX4 U10246 ( .A(n9447), .Z(n9444) );
  HS65_LH_BFX4 U10249 ( .A(n9450), .Z(n9447) );
  HS65_LH_BFX4 U10252 ( .A(n9452), .Z(n9450) );
  HS65_LH_BFX4 U10254 ( .A(n9455), .Z(n9452) );
  HS65_LH_BFX4 U10257 ( .A(n9458), .Z(n9455) );
  HS65_LH_BFX4 U10260 ( .A(n9461), .Z(n9458) );
  HS65_LH_BFX4 U10263 ( .A(n9464), .Z(n9461) );
  HS65_LH_BFX4 U10266 ( .A(n9466), .Z(n9464) );
  HS65_LH_BFX4 U10268 ( .A(n9468), .Z(n9466) );
  HS65_LH_BFX4 U10270 ( .A(n9470), .Z(n9468) );
  HS65_LH_BFX4 U10272 ( .A(n9472), .Z(n9470) );
  HS65_LH_BFX4 U10274 ( .A(n9474), .Z(n9472) );
  HS65_LH_BFX4 U10276 ( .A(n9475), .Z(n9474) );
  HS65_LH_BFX4 U10277 ( .A(n9476), .Z(n9475) );
  HS65_LH_BFX4 U10278 ( .A(\u_DataPath/u_idexreg/N40 ), .Z(n9476) );
  HS65_LH_BFX4 U10279 ( .A(n9479), .Z(n9477) );
  HS65_LH_BFX4 U10280 ( .A(\u_DataPath/immediate_ext_dec_i [2]), .Z(n9478) );
  HS65_LH_BFX4 U10281 ( .A(n11675), .Z(n9479) );
  HS65_LH_BFX4 U10282 ( .A(n9481), .Z(n9480) );
  HS65_LH_BFX4 U10283 ( .A(n9482), .Z(n9481) );
  HS65_LH_BFX4 U10284 ( .A(n13642), .Z(n9482) );
  HS65_LH_BFX4 U10285 ( .A(n9484), .Z(n9483) );
  HS65_LH_BFX4 U10286 ( .A(n9485), .Z(n9484) );
  HS65_LH_BFX4 U10287 ( .A(n9486), .Z(n9485) );
  HS65_LH_BFX4 U10288 ( .A(n9487), .Z(n9486) );
  HS65_LH_BFX4 U10289 ( .A(n9488), .Z(n9487) );
  HS65_LH_BFX4 U10290 ( .A(n9489), .Z(n9488) );
  HS65_LH_BFX4 U10291 ( .A(n9490), .Z(n9489) );
  HS65_LH_BFX4 U10292 ( .A(n9491), .Z(n9490) );
  HS65_LH_BFX4 U10293 ( .A(n9492), .Z(n9491) );
  HS65_LH_BFX4 U10294 ( .A(n9493), .Z(n9492) );
  HS65_LH_BFX4 U10295 ( .A(n9494), .Z(n9493) );
  HS65_LH_BFX4 U10296 ( .A(n9495), .Z(n9494) );
  HS65_LH_BFX4 U10297 ( .A(n9496), .Z(n9495) );
  HS65_LH_BFX4 U10298 ( .A(n9497), .Z(n9496) );
  HS65_LH_BFX4 U10299 ( .A(n9498), .Z(n9497) );
  HS65_LH_BFX4 U10300 ( .A(n9499), .Z(n9498) );
  HS65_LH_BFX4 U10301 ( .A(n9500), .Z(n9499) );
  HS65_LH_BFX4 U10302 ( .A(n9501), .Z(n9500) );
  HS65_LH_BFX4 U10303 ( .A(n9502), .Z(n9501) );
  HS65_LH_BFX4 U10304 ( .A(n9503), .Z(n9502) );
  HS65_LH_BFX4 U10305 ( .A(n9504), .Z(n9503) );
  HS65_LH_BFX4 U10306 ( .A(n9505), .Z(n9504) );
  HS65_LH_BFX4 U10307 ( .A(n9506), .Z(n9505) );
  HS65_LH_BFX4 U10308 ( .A(n9507), .Z(n9506) );
  HS65_LH_BFX4 U10309 ( .A(\u_DataPath/u_exmemreg/N12 ), .Z(n9507) );
  HS65_LH_BFX2 U10310 ( .A(n40907), .Z(n9508) );
  HS65_LH_BFX4 U10326 ( .A(n9526), .Z(n9524) );
  HS65_LH_BFX4 U10328 ( .A(n9528), .Z(n9526) );
  HS65_LH_BFX4 U10330 ( .A(n9532), .Z(n9528) );
  HS65_LH_BFX4 U10334 ( .A(n9533), .Z(n9532) );
  HS65_LH_BFX4 U10335 ( .A(n9535), .Z(n9533) );
  HS65_LH_BFX4 U10337 ( .A(n9539), .Z(n9535) );
  HS65_LH_BFX4 U10340 ( .A(n9551), .Z(n9538) );
  HS65_LH_BFX4 U10341 ( .A(n9541), .Z(n9539) );
  HS65_LH_BFX4 U10342 ( .A(\u_DataPath/regfile_addr_out_towb_i [3]), .Z(n9540)
         );
  HS65_LH_BFX4 U10343 ( .A(n9543), .Z(n9541) );
  HS65_LH_BFX4 U10345 ( .A(n9545), .Z(n9543) );
  HS65_LH_CNIVX3 U10346 ( .A(n9548), .Z(n9544) );
  HS65_LH_CNIVX3 U10347 ( .A(n9544), .Z(n9545) );
  HS65_LH_BFX4 U10350 ( .A(n9550), .Z(n9548) );
  HS65_LH_BFX4 U10352 ( .A(n9552), .Z(n9550) );
  HS65_LH_BFX4 U10353 ( .A(\u_DataPath/reg_write_i ), .Z(n9551) );
  HS65_LH_BFX4 U10354 ( .A(n9553), .Z(n9552) );
  HS65_LH_BFX4 U10355 ( .A(n9554), .Z(n9553) );
  HS65_LH_BFX4 U10356 ( .A(n9555), .Z(n9554) );
  HS65_LH_BFX4 U10357 ( .A(n9556), .Z(n9555) );
  HS65_LH_BFX4 U10358 ( .A(n9557), .Z(n9556) );
  HS65_LH_BFX4 U10359 ( .A(n9558), .Z(n9557) );
  HS65_LH_BFX4 U10360 ( .A(n9559), .Z(n9558) );
  HS65_LH_BFX4 U10361 ( .A(n15210), .Z(n9559) );
  HS65_LH_BFX4 U10362 ( .A(n9564), .Z(n9560) );
  HS65_LH_BFX4 U10363 ( .A(\u_DataPath/RFaddr_out_memwb_i [0]), .Z(n9561) );
  HS65_LH_BFX4 U10364 ( .A(n9561), .Z(n9562) );
  HS65_LH_BFX4 U10365 ( .A(n9562), .Z(n9563) );
  HS65_LH_BFX4 U10366 ( .A(n14039), .Z(n9564) );
  HS65_LH_BFX4 U10367 ( .A(n9563), .Z(n9565) );
  HS65_LH_BFX4 U10368 ( .A(n9565), .Z(n9566) );
  HS65_LH_BFX4 U10369 ( .A(n9566), .Z(n9567) );
  HS65_LH_BFX4 U10370 ( .A(n9569), .Z(n9568) );
  HS65_LH_BFX4 U10371 ( .A(n9570), .Z(n9569) );
  HS65_LH_BFX4 U10372 ( .A(n9571), .Z(n9570) );
  HS65_LH_BFX4 U10373 ( .A(n9572), .Z(n9571) );
  HS65_LH_BFX4 U10374 ( .A(n9573), .Z(n9572) );
  HS65_LH_BFX4 U10375 ( .A(n9574), .Z(n9573) );
  HS65_LH_BFX4 U10376 ( .A(n9575), .Z(n9574) );
  HS65_LH_BFX4 U10377 ( .A(n9576), .Z(n9575) );
  HS65_LH_BFX4 U10378 ( .A(n9577), .Z(n9576) );
  HS65_LH_BFX4 U10379 ( .A(n9578), .Z(n9577) );
  HS65_LH_BFX4 U10380 ( .A(n9579), .Z(n9578) );
  HS65_LH_BFX4 U10381 ( .A(n9580), .Z(n9579) );
  HS65_LH_BFX4 U10382 ( .A(n9581), .Z(n9580) );
  HS65_LH_BFX4 U10383 ( .A(n9582), .Z(n9581) );
  HS65_LH_BFX4 U10384 ( .A(n9567), .Z(n9582) );
  HS65_LH_BFX4 U10385 ( .A(n9585), .Z(n9583) );
  HS65_LH_BFX4 U10386 ( .A(n9586), .Z(n9584) );
  HS65_LH_BFX4 U10387 ( .A(n9591), .Z(n9585) );
  HS65_LH_BFX4 U10388 ( .A(n9588), .Z(n9586) );
  HS65_LH_BFX4 U10389 ( .A(n9602), .Z(n9587) );
  HS65_LH_BFX4 U10390 ( .A(n9590), .Z(n9588) );
  HS65_LH_BFX4 U10391 ( .A(n9599), .Z(n9589) );
  HS65_LH_BFX4 U10392 ( .A(n9592), .Z(n9590) );
  HS65_LH_BFX4 U10393 ( .A(n9593), .Z(n9591) );
  HS65_LH_BFX4 U10394 ( .A(n9594), .Z(n9592) );
  HS65_LH_BFX4 U10395 ( .A(n9595), .Z(n9593) );
  HS65_LH_BFX4 U10396 ( .A(n9596), .Z(n9594) );
  HS65_LH_BFX4 U10397 ( .A(n9597), .Z(n9595) );
  HS65_LH_BFX4 U10398 ( .A(n9600), .Z(n9596) );
  HS65_LH_BFX4 U10399 ( .A(n9589), .Z(n9597) );
  HS65_LH_CNIVX3 U10400 ( .A(n9587), .Z(n9598) );
  HS65_LH_CNIVX3 U10401 ( .A(n9598), .Z(n9599) );
  HS65_LH_BFX4 U10402 ( .A(n9601), .Z(n9600) );
  HS65_LH_BFX4 U10403 ( .A(n9605), .Z(n9601) );
  HS65_LH_BFX4 U10404 ( .A(n9604), .Z(n9602) );
  HS65_LH_CNIVX3 U10405 ( .A(n9607), .Z(n9603) );
  HS65_LH_CNIVX3 U10406 ( .A(n9603), .Z(n9604) );
  HS65_LH_BFX4 U10407 ( .A(n9608), .Z(n9605) );
  HS65_LH_CNIVX3 U10408 ( .A(n9610), .Z(n9606) );
  HS65_LH_CNIVX3 U10409 ( .A(n9606), .Z(n9607) );
  HS65_LH_BFX4 U10410 ( .A(n9611), .Z(n9608) );
  HS65_LH_CNIVX3 U10411 ( .A(n9613), .Z(n9609) );
  HS65_LH_CNIVX3 U10412 ( .A(n9609), .Z(n9610) );
  HS65_LH_BFX4 U10413 ( .A(n9614), .Z(n9611) );
  HS65_LH_CNIVX3 U10414 ( .A(n9616), .Z(n9612) );
  HS65_LH_CNIVX3 U10415 ( .A(n9612), .Z(n9613) );
  HS65_LH_BFX4 U10416 ( .A(n9617), .Z(n9614) );
  HS65_LH_CNIVX3 U10417 ( .A(n9619), .Z(n9615) );
  HS65_LH_CNIVX3 U10418 ( .A(n9615), .Z(n9616) );
  HS65_LH_BFX4 U10419 ( .A(n9620), .Z(n9617) );
  HS65_LH_CNIVX3 U10420 ( .A(n9622), .Z(n9618) );
  HS65_LH_CNIVX3 U10421 ( .A(n9618), .Z(n9619) );
  HS65_LH_BFX4 U10422 ( .A(n9623), .Z(n9620) );
  HS65_LH_CNIVX3 U10423 ( .A(n9625), .Z(n9621) );
  HS65_LH_CNIVX3 U10424 ( .A(n9621), .Z(n9622) );
  HS65_LH_BFX4 U10425 ( .A(n9626), .Z(n9623) );
  HS65_LH_CNIVX3 U10426 ( .A(n9628), .Z(n9624) );
  HS65_LH_CNIVX3 U10427 ( .A(n9624), .Z(n9625) );
  HS65_LH_BFX4 U10428 ( .A(n9629), .Z(n9626) );
  HS65_LH_CNIVX3 U10429 ( .A(n9631), .Z(n9627) );
  HS65_LH_CNIVX3 U10430 ( .A(n9627), .Z(n9628) );
  HS65_LH_BFX4 U10431 ( .A(n9632), .Z(n9629) );
  HS65_LH_CNIVX3 U10432 ( .A(n9634), .Z(n9630) );
  HS65_LH_CNIVX3 U10433 ( .A(n9630), .Z(n9631) );
  HS65_LH_BFX4 U10434 ( .A(n9635), .Z(n9632) );
  HS65_LH_CNIVX3 U10435 ( .A(n9637), .Z(n9633) );
  HS65_LH_CNIVX3 U10436 ( .A(n9633), .Z(n9634) );
  HS65_LH_BFX4 U10437 ( .A(n9638), .Z(n9635) );
  HS65_LH_CNIVX3 U10438 ( .A(n9642), .Z(n9636) );
  HS65_LH_CNIVX3 U10439 ( .A(n9636), .Z(n9637) );
  HS65_LH_BFX4 U10440 ( .A(n9639), .Z(n9638) );
  HS65_LH_BFX4 U10441 ( .A(n9640), .Z(n9639) );
  HS65_LH_BFX4 U10442 ( .A(n9643), .Z(n9640) );
  HS65_LH_CNIVX3 U10443 ( .A(n9641), .Z(n9642) );
  HS65_LH_BFX4 U10444 ( .A(n9644), .Z(n9643) );
  HS65_LH_BFX4 U10445 ( .A(\u_DataPath/u_idexreg/N36 ), .Z(n9644) );
  HS65_LH_BFX4 U10446 ( .A(n9649), .Z(n9645) );
  HS65_LH_BFX4 U10447 ( .A(\u_DataPath/RFaddr_out_memwb_i [1]), .Z(n9646) );
  HS65_LH_BFX4 U10448 ( .A(n9646), .Z(n9647) );
  HS65_LH_BFX4 U10449 ( .A(n9647), .Z(n9648) );
  HS65_LH_BFX4 U10450 ( .A(n14040), .Z(n9649) );
  HS65_LH_BFX4 U10451 ( .A(n9648), .Z(n9650) );
  HS65_LH_BFX4 U10452 ( .A(n9650), .Z(n9651) );
  HS65_LH_BFX4 U10453 ( .A(n9653), .Z(n9652) );
  HS65_LH_BFX4 U10454 ( .A(n9654), .Z(n9653) );
  HS65_LH_BFX4 U10455 ( .A(n9655), .Z(n9654) );
  HS65_LH_BFX4 U10456 ( .A(n9656), .Z(n9655) );
  HS65_LH_BFX4 U10457 ( .A(n9657), .Z(n9656) );
  HS65_LH_BFX4 U10458 ( .A(n9658), .Z(n9657) );
  HS65_LH_BFX4 U10459 ( .A(n9659), .Z(n9658) );
  HS65_LH_BFX4 U10460 ( .A(n9660), .Z(n9659) );
  HS65_LH_BFX4 U10461 ( .A(n9661), .Z(n9660) );
  HS65_LH_BFX4 U10462 ( .A(n9662), .Z(n9661) );
  HS65_LH_BFX4 U10463 ( .A(n9663), .Z(n9662) );
  HS65_LH_BFX4 U10464 ( .A(n9664), .Z(n9663) );
  HS65_LH_BFX4 U10465 ( .A(n9665), .Z(n9664) );
  HS65_LH_BFX4 U10466 ( .A(n9666), .Z(n9665) );
  HS65_LH_BFX4 U10467 ( .A(n9667), .Z(n9666) );
  HS65_LH_BFX4 U10468 ( .A(n9651), .Z(n9667) );
  HS65_LH_BFX4 U10469 ( .A(n9670), .Z(n9668) );
  HS65_LH_BFX4 U10470 ( .A(n9671), .Z(n9669) );
  HS65_LH_BFX4 U10471 ( .A(n9672), .Z(n9670) );
  HS65_LH_BFX4 U10472 ( .A(n9673), .Z(n9671) );
  HS65_LH_BFX4 U10473 ( .A(n9674), .Z(n9672) );
  HS65_LH_BFX4 U10474 ( .A(n9675), .Z(n9673) );
  HS65_LH_BFX4 U10475 ( .A(n9676), .Z(n9674) );
  HS65_LH_BFX4 U10476 ( .A(n9677), .Z(n9675) );
  HS65_LH_BFX4 U10477 ( .A(n9678), .Z(n9676) );
  HS65_LH_BFX4 U10478 ( .A(n9679), .Z(n9677) );
  HS65_LH_BFX4 U10479 ( .A(n9680), .Z(n9678) );
  HS65_LH_BFX4 U10480 ( .A(n9681), .Z(n9679) );
  HS65_LH_BFX4 U10481 ( .A(n9682), .Z(n9680) );
  HS65_LH_BFX4 U10482 ( .A(n9683), .Z(n9681) );
  HS65_LH_BFX4 U10483 ( .A(n9684), .Z(n9682) );
  HS65_LH_BFX4 U10484 ( .A(n9685), .Z(n9683) );
  HS65_LH_BFX4 U10485 ( .A(n9686), .Z(n9684) );
  HS65_LH_BFX4 U10486 ( .A(n9687), .Z(n9685) );
  HS65_LH_BFX4 U10487 ( .A(n9688), .Z(n9686) );
  HS65_LH_BFX4 U10488 ( .A(n9689), .Z(n9687) );
  HS65_LH_BFX4 U10489 ( .A(n9690), .Z(n9688) );
  HS65_LH_BFX4 U10490 ( .A(n9691), .Z(n9689) );
  HS65_LH_BFX4 U10491 ( .A(n9692), .Z(n9690) );
  HS65_LH_BFX4 U10492 ( .A(n9693), .Z(n9691) );
  HS65_LH_BFX4 U10493 ( .A(n9694), .Z(n9692) );
  HS65_LH_BFX4 U10494 ( .A(n9695), .Z(n9693) );
  HS65_LH_BFX4 U10495 ( .A(n9696), .Z(n9694) );
  HS65_LH_BFX4 U10496 ( .A(n9697), .Z(n9695) );
  HS65_LH_BFX4 U10497 ( .A(n9698), .Z(n9696) );
  HS65_LH_BFX4 U10498 ( .A(n9699), .Z(n9697) );
  HS65_LH_BFX4 U10499 ( .A(n9700), .Z(n9698) );
  HS65_LH_BFX4 U10500 ( .A(n9701), .Z(n9699) );
  HS65_LH_BFX4 U10501 ( .A(n13537), .Z(n9700) );
  HS65_LH_BFX4 U10502 ( .A(n9703), .Z(n9701) );
  HS65_LH_BFX4 U10503 ( .A(\u_DataPath/u_idexreg/N42 ), .Z(n9702) );
  HS65_LH_BFX4 U10504 ( .A(n9705), .Z(n9703) );
  HS65_LH_BFX4 U10505 ( .A(n9702), .Z(n9704) );
  HS65_LH_BFX4 U10506 ( .A(n9707), .Z(n9705) );
  HS65_LH_BFX4 U10507 ( .A(n9704), .Z(n9706) );
  HS65_LH_BFX4 U10508 ( .A(n9709), .Z(n9707) );
  HS65_LH_BFX4 U10509 ( .A(n9706), .Z(n9708) );
  HS65_LH_BFX4 U10510 ( .A(n9711), .Z(n9709) );
  HS65_LH_BFX4 U10511 ( .A(n9708), .Z(n9710) );
  HS65_LH_BFX4 U10512 ( .A(n9712), .Z(n9711) );
  HS65_LH_BFX4 U10513 ( .A(n9713), .Z(n9712) );
  HS65_LH_BFX4 U10514 ( .A(n9714), .Z(n9713) );
  HS65_LH_BFX4 U10515 ( .A(\u_DataPath/u_idexreg/N37 ), .Z(n9714) );
  HS65_LH_BFX4 U10516 ( .A(n9717), .Z(n9715) );
  HS65_LH_BFX4 U10517 ( .A(\u_DataPath/RFaddr_out_memwb_i [2]), .Z(n9716) );
  HS65_LH_BFX4 U10518 ( .A(n14041), .Z(n9717) );
  HS65_LH_BFX4 U10519 ( .A(n9716), .Z(n9718) );
  HS65_LH_BFX4 U10520 ( .A(n9718), .Z(n9719) );
  HS65_LH_BFX4 U10521 ( .A(n9719), .Z(n9720) );
  HS65_LH_BFX4 U10522 ( .A(n9720), .Z(n9721) );
  HS65_LH_BFX4 U10523 ( .A(n9723), .Z(n9722) );
  HS65_LH_BFX4 U10524 ( .A(n9724), .Z(n9723) );
  HS65_LH_BFX4 U10525 ( .A(n9725), .Z(n9724) );
  HS65_LH_BFX4 U10526 ( .A(n9726), .Z(n9725) );
  HS65_LH_BFX4 U10527 ( .A(n9727), .Z(n9726) );
  HS65_LH_BFX4 U10528 ( .A(n9728), .Z(n9727) );
  HS65_LH_BFX4 U10529 ( .A(n9729), .Z(n9728) );
  HS65_LH_BFX4 U10530 ( .A(n9730), .Z(n9729) );
  HS65_LH_BFX4 U10531 ( .A(n9731), .Z(n9730) );
  HS65_LH_BFX4 U10532 ( .A(n9732), .Z(n9731) );
  HS65_LH_BFX4 U10533 ( .A(n9733), .Z(n9732) );
  HS65_LH_BFX4 U10534 ( .A(n9734), .Z(n9733) );
  HS65_LH_BFX4 U10535 ( .A(n9735), .Z(n9734) );
  HS65_LH_BFX4 U10536 ( .A(n9736), .Z(n9735) );
  HS65_LH_BFX4 U10537 ( .A(n9737), .Z(n9736) );
  HS65_LH_BFX4 U10538 ( .A(n9721), .Z(n9737) );
  HS65_LH_BFX4 U10539 ( .A(n9740), .Z(n9738) );
  HS65_LH_BFX4 U10540 ( .A(n9741), .Z(n9739) );
  HS65_LH_BFX4 U10541 ( .A(n9746), .Z(n9740) );
  HS65_LH_BFX4 U10542 ( .A(n9743), .Z(n9741) );
  HS65_LH_BFX4 U10543 ( .A(n9744), .Z(n9742) );
  HS65_LH_BFX4 U10544 ( .A(n9745), .Z(n9743) );
  HS65_LH_BFX4 U10545 ( .A(n9752), .Z(n9744) );
  HS65_LH_BFX4 U10546 ( .A(n9747), .Z(n9745) );
  HS65_LH_BFX4 U10547 ( .A(n9748), .Z(n9746) );
  HS65_LH_BFX4 U10548 ( .A(n9749), .Z(n9747) );
  HS65_LH_BFX4 U10549 ( .A(n9750), .Z(n9748) );
  HS65_LH_BFX4 U10550 ( .A(n9751), .Z(n9749) );
  HS65_LH_BFX4 U10551 ( .A(n9742), .Z(n9750) );
  HS65_LH_BFX4 U10552 ( .A(n9753), .Z(n9751) );
  HS65_LH_BFX4 U10553 ( .A(n9754), .Z(n9752) );
  HS65_LH_BFX4 U10554 ( .A(n9757), .Z(n9753) );
  HS65_LH_BFX4 U10555 ( .A(n9756), .Z(n9754) );
  HS65_LH_CNIVX3 U10556 ( .A(n9759), .Z(n9755) );
  HS65_LH_CNIVX3 U10557 ( .A(n9755), .Z(n9756) );
  HS65_LH_BFX4 U10558 ( .A(n9758), .Z(n9757) );
  HS65_LH_BFX4 U10559 ( .A(n9762), .Z(n9758) );
  HS65_LH_BFX4 U10560 ( .A(n9761), .Z(n9759) );
  HS65_LH_CNIVX3 U10561 ( .A(n9764), .Z(n9760) );
  HS65_LH_CNIVX3 U10562 ( .A(n9760), .Z(n9761) );
  HS65_LH_BFX4 U10563 ( .A(n9765), .Z(n9762) );
  HS65_LH_CNIVX3 U10564 ( .A(n9767), .Z(n9763) );
  HS65_LH_CNIVX3 U10565 ( .A(n9763), .Z(n9764) );
  HS65_LH_BFX4 U10566 ( .A(n9768), .Z(n9765) );
  HS65_LH_CNIVX3 U10567 ( .A(n9770), .Z(n9766) );
  HS65_LH_CNIVX3 U10568 ( .A(n9766), .Z(n9767) );
  HS65_LH_BFX4 U10569 ( .A(n9769), .Z(n9768) );
  HS65_LH_BFX4 U10570 ( .A(n9773), .Z(n9769) );
  HS65_LH_BFX4 U10571 ( .A(n9772), .Z(n9770) );
  HS65_LH_CNIVX3 U10572 ( .A(n9775), .Z(n9771) );
  HS65_LH_CNIVX3 U10573 ( .A(n9771), .Z(n9772) );
  HS65_LH_BFX4 U10574 ( .A(n9776), .Z(n9773) );
  HS65_LH_CNIVX3 U10575 ( .A(n9778), .Z(n9774) );
  HS65_LH_CNIVX3 U10576 ( .A(n9774), .Z(n9775) );
  HS65_LH_BFX4 U10577 ( .A(n9779), .Z(n9776) );
  HS65_LH_CNIVX3 U10578 ( .A(n9781), .Z(n9777) );
  HS65_LH_CNIVX3 U10579 ( .A(n9777), .Z(n9778) );
  HS65_LH_BFX4 U10580 ( .A(n9782), .Z(n9779) );
  HS65_LH_CNIVX3 U10581 ( .A(n9784), .Z(n9780) );
  HS65_LH_CNIVX3 U10582 ( .A(n9780), .Z(n9781) );
  HS65_LH_BFX4 U10583 ( .A(n9785), .Z(n9782) );
  HS65_LH_CNIVX3 U10584 ( .A(n9787), .Z(n9783) );
  HS65_LH_CNIVX3 U10585 ( .A(n9783), .Z(n9784) );
  HS65_LH_BFX4 U10586 ( .A(n9788), .Z(n9785) );
  HS65_LH_CNIVX3 U10587 ( .A(n9790), .Z(n9786) );
  HS65_LH_CNIVX3 U10588 ( .A(n9786), .Z(n9787) );
  HS65_LH_BFX4 U10589 ( .A(n9791), .Z(n9788) );
  HS65_LH_CNIVX3 U10590 ( .A(n9795), .Z(n9789) );
  HS65_LH_CNIVX3 U10591 ( .A(n9789), .Z(n9790) );
  HS65_LH_BFX4 U10592 ( .A(n9792), .Z(n9791) );
  HS65_LH_BFX4 U10593 ( .A(n9793), .Z(n9792) );
  HS65_LH_BFX4 U10594 ( .A(n9796), .Z(n9793) );
  HS65_LH_CNIVX3 U10595 ( .A(n9794), .Z(n9795) );
  HS65_LH_BFX4 U10596 ( .A(n9797), .Z(n9796) );
  HS65_LH_BFX4 U10597 ( .A(\u_DataPath/u_idexreg/N38 ), .Z(n9797) );
  HS65_LH_BFX4 U10598 ( .A(n9801), .Z(n9798) );
  HS65_LH_BFX4 U10599 ( .A(\u_DataPath/RFaddr_out_memwb_i [3]), .Z(n9799) );
  HS65_LH_BFX4 U10600 ( .A(n9799), .Z(n9800) );
  HS65_LH_BFX4 U10601 ( .A(n14042), .Z(n9801) );
  HS65_LH_BFX4 U10602 ( .A(n9800), .Z(n9802) );
  HS65_LH_BFX4 U10603 ( .A(n9804), .Z(n9803) );
  HS65_LH_BFX4 U10604 ( .A(n9805), .Z(n9804) );
  HS65_LH_BFX4 U10605 ( .A(n9806), .Z(n9805) );
  HS65_LH_BFX4 U10606 ( .A(n9807), .Z(n9806) );
  HS65_LH_BFX4 U10607 ( .A(n9808), .Z(n9807) );
  HS65_LH_BFX4 U10608 ( .A(n9809), .Z(n9808) );
  HS65_LH_BFX4 U10609 ( .A(n9810), .Z(n9809) );
  HS65_LH_BFX4 U10610 ( .A(n9811), .Z(n9810) );
  HS65_LH_BFX4 U10611 ( .A(n9812), .Z(n9811) );
  HS65_LH_BFX4 U10612 ( .A(n9813), .Z(n9812) );
  HS65_LH_BFX4 U10613 ( .A(n9814), .Z(n9813) );
  HS65_LH_BFX4 U10614 ( .A(n9815), .Z(n9814) );
  HS65_LH_BFX4 U10615 ( .A(n9816), .Z(n9815) );
  HS65_LH_BFX4 U10616 ( .A(n9817), .Z(n9816) );
  HS65_LH_BFX4 U10617 ( .A(n9818), .Z(n9817) );
  HS65_LH_BFX4 U10618 ( .A(n9819), .Z(n9818) );
  HS65_LH_BFX4 U10619 ( .A(n9820), .Z(n9819) );
  HS65_LH_BFX4 U10620 ( .A(n9802), .Z(n9820) );
  HS65_LH_BFX4 U10621 ( .A(n9823), .Z(n9821) );
  HS65_LH_BFX4 U10622 ( .A(n9824), .Z(n9822) );
  HS65_LH_BFX4 U10623 ( .A(n9825), .Z(n9823) );
  HS65_LH_BFX4 U10624 ( .A(n9826), .Z(n9824) );
  HS65_LH_BFX4 U10625 ( .A(n9827), .Z(n9825) );
  HS65_LH_BFX4 U10626 ( .A(n9828), .Z(n9826) );
  HS65_LH_BFX4 U10627 ( .A(n9829), .Z(n9827) );
  HS65_LH_BFX4 U10628 ( .A(n9830), .Z(n9828) );
  HS65_LH_BFX4 U10629 ( .A(n9831), .Z(n9829) );
  HS65_LH_BFX4 U10630 ( .A(n9832), .Z(n9830) );
  HS65_LH_BFX4 U10631 ( .A(n9833), .Z(n9831) );
  HS65_LH_BFX4 U10632 ( .A(n9834), .Z(n9832) );
  HS65_LH_BFX4 U10633 ( .A(n9835), .Z(n9833) );
  HS65_LH_BFX4 U10634 ( .A(n9836), .Z(n9834) );
  HS65_LH_BFX4 U10635 ( .A(n9837), .Z(n9835) );
  HS65_LH_BFX4 U10636 ( .A(n9838), .Z(n9836) );
  HS65_LH_BFX4 U10637 ( .A(n9839), .Z(n9837) );
  HS65_LH_BFX4 U10638 ( .A(n9840), .Z(n9838) );
  HS65_LH_BFX4 U10639 ( .A(n9841), .Z(n9839) );
  HS65_LH_BFX4 U10640 ( .A(n9842), .Z(n9840) );
  HS65_LH_BFX4 U10641 ( .A(n9843), .Z(n9841) );
  HS65_LH_BFX4 U10642 ( .A(n9844), .Z(n9842) );
  HS65_LH_BFX4 U10643 ( .A(n9845), .Z(n9843) );
  HS65_LH_BFX4 U10644 ( .A(n9846), .Z(n9844) );
  HS65_LH_BFX4 U10645 ( .A(n9847), .Z(n9845) );
  HS65_LH_BFX4 U10646 ( .A(n9848), .Z(n9846) );
  HS65_LH_BFX4 U10647 ( .A(n9849), .Z(n9847) );
  HS65_LH_BFX4 U10648 ( .A(n9850), .Z(n9848) );
  HS65_LH_BFX4 U10649 ( .A(n9851), .Z(n9849) );
  HS65_LH_BFX4 U10650 ( .A(n9852), .Z(n9850) );
  HS65_LH_BFX4 U10651 ( .A(n9853), .Z(n9851) );
  HS65_LH_BFX4 U10652 ( .A(n9854), .Z(n9852) );
  HS65_LH_BFX4 U10653 ( .A(n9855), .Z(n9853) );
  HS65_LH_BFX4 U10654 ( .A(n9856), .Z(n9854) );
  HS65_LH_BFX4 U10655 ( .A(n9857), .Z(n9855) );
  HS65_LH_BFX4 U10656 ( .A(n9858), .Z(n9856) );
  HS65_LH_BFX4 U10657 ( .A(n9859), .Z(n9857) );
  HS65_LH_BFX4 U10658 ( .A(n9860), .Z(n9858) );
  HS65_LH_BFX4 U10659 ( .A(n9861), .Z(n9859) );
  HS65_LH_BFX4 U10660 ( .A(n13531), .Z(n9860) );
  HS65_LH_BFX4 U10661 ( .A(n9863), .Z(n9861) );
  HS65_LH_BFX4 U10662 ( .A(\u_DataPath/u_idexreg/N44 ), .Z(n9862) );
  HS65_LH_BFX4 U10663 ( .A(n9865), .Z(n9863) );
  HS65_LH_BFX4 U10664 ( .A(n9862), .Z(n9864) );
  HS65_LH_BFX4 U10665 ( .A(n9866), .Z(n9865) );
  HS65_LH_BFX4 U10666 ( .A(n9867), .Z(n9866) );
  HS65_LH_BFX4 U10667 ( .A(\u_DataPath/u_idexreg/N39 ), .Z(n9867) );
  HS65_LH_BFX4 U10668 ( .A(n9871), .Z(n9868) );
  HS65_LH_BFX4 U10669 ( .A(n9872), .Z(n9869) );
  HS65_LH_BFX4 U10670 ( .A(n9873), .Z(n9870) );
  HS65_LH_BFX4 U10671 ( .A(n9874), .Z(n9871) );
  HS65_LH_BFX4 U10672 ( .A(n9875), .Z(n9872) );
  HS65_LH_BFX4 U10673 ( .A(n9876), .Z(n9873) );
  HS65_LH_BFX4 U10674 ( .A(n9880), .Z(n9874) );
  HS65_LH_BFX4 U10675 ( .A(n9878), .Z(n9875) );
  HS65_LH_BFX4 U10676 ( .A(n9879), .Z(n9876) );
  HS65_LH_BFX4 U10677 ( .A(\u_DataPath/u_idexreg/N19 ), .Z(n9877) );
  HS65_LH_BFX4 U10678 ( .A(n9881), .Z(n9878) );
  HS65_LH_BFX4 U10679 ( .A(n9882), .Z(n9879) );
  HS65_LH_BFX4 U10680 ( .A(n9883), .Z(n9880) );
  HS65_LH_BFX4 U10681 ( .A(n9884), .Z(n9881) );
  HS65_LH_BFX4 U10682 ( .A(n9885), .Z(n9882) );
  HS65_LH_BFX4 U10683 ( .A(n9886), .Z(n9883) );
  HS65_LH_BFX4 U10684 ( .A(n9887), .Z(n9884) );
  HS65_LH_BFX4 U10685 ( .A(n9888), .Z(n9885) );
  HS65_LH_BFX4 U10686 ( .A(n9889), .Z(n9886) );
  HS65_LH_BFX4 U10687 ( .A(n9890), .Z(n9887) );
  HS65_LH_BFX4 U10688 ( .A(n9891), .Z(n9888) );
  HS65_LH_BFX4 U10689 ( .A(n9893), .Z(n9889) );
  HS65_LH_BFX4 U10690 ( .A(n9892), .Z(n9890) );
  HS65_LH_BFX4 U10691 ( .A(n9898), .Z(n9891) );
  HS65_LH_BFX4 U10692 ( .A(n9897), .Z(n9892) );
  HS65_LH_BFX4 U10693 ( .A(n9895), .Z(n9893) );
  HS65_LH_CNIVX3 U10694 ( .A(n9900), .Z(n9894) );
  HS65_LH_CNIVX3 U10695 ( .A(n9894), .Z(n9895) );
  HS65_LH_CNIVX3 U10696 ( .A(n9902), .Z(n9896) );
  HS65_LH_CNIVX3 U10697 ( .A(n9896), .Z(n9897) );
  HS65_LH_BFX4 U10698 ( .A(n9903), .Z(n9898) );
  HS65_LH_CNIVX3 U10699 ( .A(n9906), .Z(n9899) );
  HS65_LH_CNIVX3 U10700 ( .A(n9899), .Z(n9900) );
  HS65_LH_CNIVX3 U10701 ( .A(n9910), .Z(n9901) );
  HS65_LH_CNIVX3 U10702 ( .A(n9901), .Z(n9902) );
  HS65_LH_BFX4 U10703 ( .A(n9904), .Z(n9903) );
  HS65_LH_BFX4 U10704 ( .A(n9911), .Z(n9904) );
  HS65_LH_BFX4 U10705 ( .A(\u_DataPath/idex_rt_i [4]), .Z(n9905) );
  HS65_LH_BFX4 U10706 ( .A(n9908), .Z(n9906) );
  HS65_LH_CNIVX3 U10707 ( .A(n9915), .Z(n9907) );
  HS65_LH_CNIVX3 U10708 ( .A(n9907), .Z(n9908) );
  HS65_LH_CNIVX3 U10709 ( .A(n9913), .Z(n9909) );
  HS65_LH_CNIVX3 U10710 ( .A(n9909), .Z(n9910) );
  HS65_LH_BFX4 U10711 ( .A(n9914), .Z(n9911) );
  HS65_LH_CNIVX3 U10712 ( .A(n9917), .Z(n9912) );
  HS65_LH_CNIVX3 U10713 ( .A(n9912), .Z(n9913) );
  HS65_LH_BFX4 U10714 ( .A(n9918), .Z(n9914) );
  HS65_LH_BFX4 U10715 ( .A(n9919), .Z(n9915) );
  HS65_LH_CNIVX3 U10716 ( .A(n9924), .Z(n9916) );
  HS65_LH_CNIVX3 U10717 ( .A(n9916), .Z(n9917) );
  HS65_LH_BFX4 U10718 ( .A(n9920), .Z(n9918) );
  HS65_LH_BFX4 U10719 ( .A(n9922), .Z(n9919) );
  HS65_LH_BFX4 U10720 ( .A(n9925), .Z(n9920) );
  HS65_LH_BFX4 U10721 ( .A(n9905), .Z(n9921) );
  HS65_LH_BFX4 U10722 ( .A(n9926), .Z(n9922) );
  HS65_LH_CNIVX3 U10723 ( .A(n9943), .Z(n9923) );
  HS65_LH_CNIVX3 U10724 ( .A(n9923), .Z(n9924) );
  HS65_LH_BFX4 U10725 ( .A(n9927), .Z(n9925) );
  HS65_LH_BFX4 U10726 ( .A(n9929), .Z(n9926) );
  HS65_LH_BFX4 U10727 ( .A(n9930), .Z(n9927) );
  HS65_LH_BFX4 U10728 ( .A(n9921), .Z(n9928) );
  HS65_LH_BFX4 U10729 ( .A(n9932), .Z(n9929) );
  HS65_LH_BFX4 U10730 ( .A(n9933), .Z(n9930) );
  HS65_LH_BFX4 U10731 ( .A(n9928), .Z(n9931) );
  HS65_LH_BFX4 U10732 ( .A(n9935), .Z(n9932) );
  HS65_LH_BFX4 U10733 ( .A(n9936), .Z(n9933) );
  HS65_LH_BFX4 U10734 ( .A(n9931), .Z(n9934) );
  HS65_LH_BFX4 U10735 ( .A(n9938), .Z(n9935) );
  HS65_LH_BFX4 U10736 ( .A(n9939), .Z(n9936) );
  HS65_LH_BFX4 U10737 ( .A(n9934), .Z(n9937) );
  HS65_LH_BFX4 U10738 ( .A(n9941), .Z(n9938) );
  HS65_LH_BFX4 U10739 ( .A(n9944), .Z(n9939) );
  HS65_LH_BFX4 U10740 ( .A(n9937), .Z(n9940) );
  HS65_LH_BFX4 U10741 ( .A(n9945), .Z(n9941) );
  HS65_LH_CNIVX3 U10742 ( .A(n9940), .Z(n9942) );
  HS65_LH_CNIVX3 U10743 ( .A(n9942), .Z(n9943) );
  HS65_LH_BFX4 U10744 ( .A(n9946), .Z(n9944) );
  HS65_LH_BFX4 U10745 ( .A(n9877), .Z(n9945) );
  HS65_LH_BFX4 U10746 ( .A(n9947), .Z(n9946) );
  HS65_LH_BFX4 U10747 ( .A(n9948), .Z(n9947) );
  HS65_LH_BFX4 U10748 ( .A(\u_DataPath/u_idexreg/N40 ), .Z(n9948) );
  HS65_LH_BFX4 U10749 ( .A(n12505), .Z(n9949) );
  HS65_LH_BFX4 U10750 ( .A(n12552), .Z(n9950) );
  HS65_LH_BFX4 U10751 ( .A(n12599), .Z(n9951) );
  HS65_LH_BFX4 U10752 ( .A(n9953), .Z(n9952) );
  HS65_LH_BFX4 U10753 ( .A(n9954), .Z(n9953) );
  HS65_LH_BFX4 U10754 ( .A(n9955), .Z(n9954) );
  HS65_LH_BFX4 U10755 ( .A(n9956), .Z(n9955) );
  HS65_LH_BFX4 U10756 ( .A(n9957), .Z(n9956) );
  HS65_LH_BFX4 U10757 ( .A(n9958), .Z(n9957) );
  HS65_LH_BFX4 U10758 ( .A(n9959), .Z(n9958) );
  HS65_LH_BFX4 U10759 ( .A(n9960), .Z(n9959) );
  HS65_LH_BFX4 U10760 ( .A(n9961), .Z(n9960) );
  HS65_LH_BFX4 U10761 ( .A(n12644), .Z(n9961) );
  HS65_LH_BFX4 U10762 ( .A(n12673), .Z(n9962) );
  HS65_LH_BFX4 U10763 ( .A(n12718), .Z(n9963) );
  HS65_LH_BFX4 U10764 ( .A(n12763), .Z(n9964) );
  HS65_LH_BFX4 U10765 ( .A(n12807), .Z(n9965) );
  HS65_LH_BFX4 U10766 ( .A(n12852), .Z(n9966) );
  HS65_LH_BFX4 U10767 ( .A(n12897), .Z(n9967) );
  HS65_LH_BFX4 U10768 ( .A(n12942), .Z(n9968) );
  HS65_LH_BFX4 U10769 ( .A(n12987), .Z(n9969) );
  HS65_LH_BFX4 U10770 ( .A(n13032), .Z(n9970) );
  HS65_LH_BFX4 U10771 ( .A(n13077), .Z(n9971) );
  HS65_LH_BFX4 U10772 ( .A(n13122), .Z(n9972) );
  HS65_LH_BFX4 U10773 ( .A(n13167), .Z(n9973) );
  HS65_LH_BFX4 U10774 ( .A(n13212), .Z(n9974) );
  HS65_LH_BFX4 U10775 ( .A(n13257), .Z(n9975) );
  HS65_LH_BFX4 U10776 ( .A(n13302), .Z(n9976) );
  HS65_LH_BFX4 U10777 ( .A(n11921), .Z(n9977) );
  HS65_LH_BFX4 U10778 ( .A(n11966), .Z(n9978) );
  HS65_LH_BFX4 U10779 ( .A(n12011), .Z(n9979) );
  HS65_LH_BFX4 U10780 ( .A(n12056), .Z(n9980) );
  HS65_LH_BFX4 U10781 ( .A(n12101), .Z(n9981) );
  HS65_LH_BFX4 U10782 ( .A(n12146), .Z(n9982) );
  HS65_LH_BFX4 U10783 ( .A(n12191), .Z(n9983) );
  HS65_LH_BFX4 U10784 ( .A(n12236), .Z(n9984) );
  HS65_LH_BFX4 U10785 ( .A(n13347), .Z(n9985) );
  HS65_LH_BFX4 U10786 ( .A(n13392), .Z(n9986) );
  HS65_LH_BFX4 U10787 ( .A(n13437), .Z(n9987) );
  HS65_LH_BFX4 U10788 ( .A(n13482), .Z(n9988) );
  HS65_LH_BFX4 U10789 ( .A(n13540), .Z(n9989) );
  HS65_LH_BFX4 U10790 ( .A(n9991), .Z(n9990) );
  HS65_LH_BFX4 U10791 ( .A(n9992), .Z(n9991) );
  HS65_LH_BFX4 U10792 ( .A(n9993), .Z(n9992) );
  HS65_LH_BFX4 U10793 ( .A(n9994), .Z(n9993) );
  HS65_LH_BFX4 U10794 ( .A(n9995), .Z(n9994) );
  HS65_LH_BFX4 U10795 ( .A(n9996), .Z(n9995) );
  HS65_LH_BFX4 U10796 ( .A(n9997), .Z(n9996) );
  HS65_LH_BFX4 U10797 ( .A(n9998), .Z(n9997) );
  HS65_LH_BFX4 U10798 ( .A(n9999), .Z(n9998) );
  HS65_LH_BFX4 U10799 ( .A(n10000), .Z(n9999) );
  HS65_LH_BFX4 U10800 ( .A(n10001), .Z(n10000) );
  HS65_LH_BFX4 U10801 ( .A(n10002), .Z(n10001) );
  HS65_LH_BFX4 U10802 ( .A(n10003), .Z(n10002) );
  HS65_LH_BFX4 U10803 ( .A(n10004), .Z(n10003) );
  HS65_LH_BFX4 U10804 ( .A(n10005), .Z(n10004) );
  HS65_LH_BFX4 U10805 ( .A(n10006), .Z(n10005) );
  HS65_LH_BFX4 U10806 ( .A(n10007), .Z(n10006) );
  HS65_LH_BFX4 U10807 ( .A(n10008), .Z(n10007) );
  HS65_LH_BFX4 U10808 ( .A(n10009), .Z(n10008) );
  HS65_LH_BFX4 U10809 ( .A(n10010), .Z(n10009) );
  HS65_LH_BFX4 U10810 ( .A(n10011), .Z(n10010) );
  HS65_LH_BFX4 U10811 ( .A(n10012), .Z(n10011) );
  HS65_LH_BFX4 U10812 ( .A(n10013), .Z(n10012) );
  HS65_LH_BFX4 U10813 ( .A(n10014), .Z(n10013) );
  HS65_LH_BFX4 U10814 ( .A(\u_DataPath/cw_memwb_i [2]), .Z(n10014) );
  HS65_LH_BFX4 U10815 ( .A(n10016), .Z(n10015) );
  HS65_LH_BFX4 U10816 ( .A(n10017), .Z(n10016) );
  HS65_LH_BFX4 U10817 ( .A(n10018), .Z(n10017) );
  HS65_LH_BFX4 U10818 ( .A(n10019), .Z(n10018) );
  HS65_LH_BFX4 U10819 ( .A(n10020), .Z(n10019) );
  HS65_LH_BFX4 U10820 ( .A(n10021), .Z(n10020) );
  HS65_LH_BFX4 U10821 ( .A(n10022), .Z(n10021) );
  HS65_LH_BFX4 U10822 ( .A(n10023), .Z(n10022) );
  HS65_LH_BFX4 U10823 ( .A(n10024), .Z(n10023) );
  HS65_LH_BFX4 U10824 ( .A(n10025), .Z(n10024) );
  HS65_LH_BFX4 U10825 ( .A(n10026), .Z(n10025) );
  HS65_LH_BFX4 U10826 ( .A(n10027), .Z(n10026) );
  HS65_LH_BFX4 U10827 ( .A(n10028), .Z(n10027) );
  HS65_LH_BFX4 U10828 ( .A(n10029), .Z(n10028) );
  HS65_LH_BFX4 U10829 ( .A(n10030), .Z(n10029) );
  HS65_LH_BFX4 U10830 ( .A(n10031), .Z(n10030) );
  HS65_LH_BFX4 U10831 ( .A(n10032), .Z(n10031) );
  HS65_LH_BFX4 U10832 ( .A(n10033), .Z(n10032) );
  HS65_LH_BFX4 U10833 ( .A(n10034), .Z(n10033) );
  HS65_LH_BFX4 U10834 ( .A(n10035), .Z(n10034) );
  HS65_LH_BFX4 U10835 ( .A(n10036), .Z(n10035) );
  HS65_LH_BFX4 U10836 ( .A(n10037), .Z(n10036) );
  HS65_LH_BFX4 U10837 ( .A(n10038), .Z(n10037) );
  HS65_LH_BFX4 U10838 ( .A(n10039), .Z(n10038) );
  HS65_LH_BFX4 U10839 ( .A(\u_DataPath/cw_exmem_i [10]), .Z(n10039) );
  HS65_LH_BFX4 U10840 ( .A(n10041), .Z(n10040) );
  HS65_LH_BFX4 U10841 ( .A(n10042), .Z(n10041) );
  HS65_LH_BFX4 U10842 ( .A(n10043), .Z(n10042) );
  HS65_LH_BFX4 U10843 ( .A(n10044), .Z(n10043) );
  HS65_LH_BFX4 U10844 ( .A(n10045), .Z(n10044) );
  HS65_LH_BFX4 U10845 ( .A(n10046), .Z(n10045) );
  HS65_LH_BFX4 U10846 ( .A(n10047), .Z(n10046) );
  HS65_LH_BFX4 U10847 ( .A(n10048), .Z(n10047) );
  HS65_LH_BFX4 U10848 ( .A(n10049), .Z(n10048) );
  HS65_LH_BFX4 U10849 ( .A(n10050), .Z(n10049) );
  HS65_LH_BFX4 U10850 ( .A(n10051), .Z(n10050) );
  HS65_LH_BFX4 U10851 ( .A(n10052), .Z(n10051) );
  HS65_LH_BFX4 U10852 ( .A(n10053), .Z(n10052) );
  HS65_LH_BFX4 U10853 ( .A(n10054), .Z(n10053) );
  HS65_LH_BFX4 U10854 ( .A(n10055), .Z(n10054) );
  HS65_LH_BFX4 U10855 ( .A(n10056), .Z(n10055) );
  HS65_LH_BFX4 U10856 ( .A(n10057), .Z(n10056) );
  HS65_LH_BFX4 U10857 ( .A(n10058), .Z(n10057) );
  HS65_LH_BFX4 U10858 ( .A(n10059), .Z(n10058) );
  HS65_LH_BFX4 U10859 ( .A(n10060), .Z(n10059) );
  HS65_LH_BFX4 U10860 ( .A(n10061), .Z(n10060) );
  HS65_LH_BFX4 U10861 ( .A(n10062), .Z(n10061) );
  HS65_LH_BFX4 U10862 ( .A(n10063), .Z(n10062) );
  HS65_LH_BFX4 U10863 ( .A(n10064), .Z(n10063) );
  HS65_LH_BFX4 U10864 ( .A(\u_DataPath/cw_memwb_i [0]), .Z(n10064) );
  HS65_LH_BFX4 U10865 ( .A(n10066), .Z(n10065) );
  HS65_LH_BFX4 U10866 ( .A(n10067), .Z(n10066) );
  HS65_LH_BFX4 U10867 ( .A(n10068), .Z(n10067) );
  HS65_LH_BFX4 U10868 ( .A(n10069), .Z(n10068) );
  HS65_LH_BFX4 U10869 ( .A(n10070), .Z(n10069) );
  HS65_LH_BFX4 U10870 ( .A(n10071), .Z(n10070) );
  HS65_LH_BFX4 U10871 ( .A(n10072), .Z(n10071) );
  HS65_LH_BFX4 U10872 ( .A(n10073), .Z(n10072) );
  HS65_LH_BFX4 U10873 ( .A(n10074), .Z(n10073) );
  HS65_LH_BFX4 U10874 ( .A(n10075), .Z(n10074) );
  HS65_LH_BFX4 U10875 ( .A(n10076), .Z(n10075) );
  HS65_LH_BFX4 U10876 ( .A(n10077), .Z(n10076) );
  HS65_LH_BFX4 U10877 ( .A(n10078), .Z(n10077) );
  HS65_LH_BFX4 U10878 ( .A(n10079), .Z(n10078) );
  HS65_LH_BFX4 U10879 ( .A(n10080), .Z(n10079) );
  HS65_LH_BFX4 U10880 ( .A(n10081), .Z(n10080) );
  HS65_LH_BFX4 U10881 ( .A(n10082), .Z(n10081) );
  HS65_LH_BFX4 U10882 ( .A(n10083), .Z(n10082) );
  HS65_LH_BFX4 U10883 ( .A(n10084), .Z(n10083) );
  HS65_LH_BFX4 U10884 ( .A(n10085), .Z(n10084) );
  HS65_LH_BFX4 U10885 ( .A(n10086), .Z(n10085) );
  HS65_LH_BFX4 U10886 ( .A(n10087), .Z(n10086) );
  HS65_LH_BFX4 U10887 ( .A(n10088), .Z(n10087) );
  HS65_LH_BFX4 U10888 ( .A(n10089), .Z(n10088) );
  HS65_LH_BFX4 U10889 ( .A(\u_DataPath/u_idexreg/N10 ), .Z(n10089) );
  HS65_LH_BFX4 U10890 ( .A(n10091), .Z(n10090) );
  HS65_LH_BFX4 U10891 ( .A(n10093), .Z(n10091) );
  HS65_LH_BFX4 U10892 ( .A(\u_DataPath/u_idexreg/N11 ), .Z(n10092) );
  HS65_LH_BFX4 U10893 ( .A(n10095), .Z(n10093) );
  HS65_LH_BFX4 U10894 ( .A(n10092), .Z(n10094) );
  HS65_LH_BFX4 U10895 ( .A(n14046), .Z(n10095) );
  HS65_LH_BFX4 U10896 ( .A(n10094), .Z(n10096) );
  HS65_LH_BFX4 U10897 ( .A(n10096), .Z(n10097) );
  HS65_LH_BFX4 U10898 ( .A(n10097), .Z(n10098) );
  HS65_LH_BFX4 U10899 ( .A(n10098), .Z(n10099) );
  HS65_LH_BFX4 U10900 ( .A(n10099), .Z(n10100) );
  HS65_LH_BFX4 U10901 ( .A(n10100), .Z(n10101) );
  HS65_LH_BFX4 U10902 ( .A(n12480), .Z(n10102) );
  HS65_LH_BFX4 U10903 ( .A(n10104), .Z(n10103) );
  HS65_LH_BFX4 U10904 ( .A(n10105), .Z(n10104) );
  HS65_LH_BFX4 U10905 ( .A(n10106), .Z(n10105) );
  HS65_LH_BFX4 U10906 ( .A(n10107), .Z(n10106) );
  HS65_LH_BFX4 U10907 ( .A(n10108), .Z(n10107) );
  HS65_LH_BFX4 U10908 ( .A(n10109), .Z(n10108) );
  HS65_LH_BFX4 U10909 ( .A(n10110), .Z(n10109) );
  HS65_LH_BFX4 U10910 ( .A(n10111), .Z(n10110) );
  HS65_LH_BFX4 U10911 ( .A(n10112), .Z(n10111) );
  HS65_LH_BFX4 U10912 ( .A(n10113), .Z(n10112) );
  HS65_LH_BFX4 U10913 ( .A(n10114), .Z(n10113) );
  HS65_LH_BFX4 U10914 ( .A(n10115), .Z(n10114) );
  HS65_LH_BFX4 U10915 ( .A(n10116), .Z(n10115) );
  HS65_LH_BFX4 U10916 ( .A(n10117), .Z(n10116) );
  HS65_LH_BFX4 U10917 ( .A(n10118), .Z(n10117) );
  HS65_LH_BFX4 U10918 ( .A(n10119), .Z(n10118) );
  HS65_LH_BFX4 U10919 ( .A(n10120), .Z(n10119) );
  HS65_LH_BFX4 U10920 ( .A(n10121), .Z(n10120) );
  HS65_LH_BFX4 U10921 ( .A(n10122), .Z(n10121) );
  HS65_LH_BFX4 U10922 ( .A(n10123), .Z(n10122) );
  HS65_LH_BFX4 U10923 ( .A(n10124), .Z(n10123) );
  HS65_LH_BFX4 U10924 ( .A(n10125), .Z(n10124) );
  HS65_LH_BFX4 U10925 ( .A(n10126), .Z(n10125) );
  HS65_LH_BFX4 U10926 ( .A(n10127), .Z(n10126) );
  HS65_LH_BFX4 U10927 ( .A(\u_DataPath/u_idexreg/N16 ), .Z(n10127) );
  HS65_LH_BFX4 U10928 ( .A(n10129), .Z(n10128) );
  HS65_LH_BFX4 U10929 ( .A(n10130), .Z(n10129) );
  HS65_LH_BFX4 U10930 ( .A(n10131), .Z(n10130) );
  HS65_LH_BFX4 U10931 ( .A(n10132), .Z(n10131) );
  HS65_LH_BFX4 U10932 ( .A(n10133), .Z(n10132) );
  HS65_LH_BFX4 U10933 ( .A(n10134), .Z(n10133) );
  HS65_LH_BFX4 U10934 ( .A(n10135), .Z(n10134) );
  HS65_LH_BFX4 U10935 ( .A(n10136), .Z(n10135) );
  HS65_LH_BFX4 U10936 ( .A(n10137), .Z(n10136) );
  HS65_LH_BFX4 U10937 ( .A(n10138), .Z(n10137) );
  HS65_LH_BFX4 U10938 ( .A(n10139), .Z(n10138) );
  HS65_LH_BFX4 U10939 ( .A(n10140), .Z(n10139) );
  HS65_LH_BFX4 U10940 ( .A(n10141), .Z(n10140) );
  HS65_LH_BFX4 U10941 ( .A(n10142), .Z(n10141) );
  HS65_LH_BFX4 U10942 ( .A(n10147), .Z(n10142) );
  HS65_LH_BFX4 U10943 ( .A(\u_DataPath/u_idexreg/N13 ), .Z(n10143) );
  HS65_LH_BFX4 U10944 ( .A(n10143), .Z(n10144) );
  HS65_LH_BFX4 U10945 ( .A(n10144), .Z(n10145) );
  HS65_LH_BFX4 U10946 ( .A(n10145), .Z(n10146) );
  HS65_LH_BFX4 U10947 ( .A(n10149), .Z(n10147) );
  HS65_LH_BFX4 U10948 ( .A(n10146), .Z(n10148) );
  HS65_LH_BFX4 U10949 ( .A(n10150), .Z(n10149) );
  HS65_LH_BFX4 U10950 ( .A(n10483), .Z(n10150) );
  HS65_LH_BFX4 U10951 ( .A(n13639), .Z(n10151) );
  HS65_LH_BFX4 U10953 ( .A(\u_DataPath/jump_i ), .Z(n10153) );
  HS65_LH_BFX4 U10954 ( .A(n10159), .Z(n10154) );
  HS65_LH_BFX4 U10955 ( .A(n10160), .Z(n10155) );
  HS65_LH_BFX4 U10956 ( .A(n12637), .Z(n10156) );
  HS65_LH_BFX4 U10958 ( .A(n10162), .Z(n10158) );
  HS65_LH_BFX4 U10959 ( .A(n10163), .Z(n10159) );
  HS65_LH_BFX4 U10960 ( .A(n10164), .Z(n10160) );
  HS65_LH_BFX4 U10962 ( .A(n10166), .Z(n10162) );
  HS65_LH_BFX4 U10963 ( .A(n10167), .Z(n10163) );
  HS65_LH_BFX4 U10964 ( .A(n10168), .Z(n10164) );
  HS65_LH_BFX4 U10966 ( .A(n10170), .Z(n10166) );
  HS65_LH_BFX4 U10967 ( .A(n10171), .Z(n10167) );
  HS65_LH_BFX4 U10968 ( .A(n10172), .Z(n10168) );
  HS65_LH_BFX4 U10970 ( .A(n10174), .Z(n10170) );
  HS65_LH_BFX4 U10971 ( .A(n10175), .Z(n10171) );
  HS65_LH_BFX4 U10972 ( .A(n10176), .Z(n10172) );
  HS65_LH_BFX4 U10974 ( .A(n10182), .Z(n10174) );
  HS65_LH_BFX4 U10975 ( .A(n10179), .Z(n10175) );
  HS65_LH_BFX4 U10976 ( .A(n10180), .Z(n10176) );
  HS65_LH_BFX4 U10978 ( .A(n10153), .Z(n10178) );
  HS65_LH_BFX4 U10979 ( .A(n10183), .Z(n10179) );
  HS65_LH_BFX4 U10980 ( .A(n10184), .Z(n10180) );
  HS65_LH_BFX4 U10982 ( .A(n10186), .Z(n10182) );
  HS65_LH_BFX4 U10983 ( .A(n10187), .Z(n10183) );
  HS65_LH_BFX4 U10984 ( .A(n10188), .Z(n10184) );
  HS65_LH_BFX4 U10986 ( .A(n10190), .Z(n10186) );
  HS65_LH_BFX4 U10987 ( .A(n10191), .Z(n10187) );
  HS65_LH_BFX4 U10988 ( .A(n10192), .Z(n10188) );
  HS65_LH_BFX4 U10990 ( .A(n10194), .Z(n10190) );
  HS65_LH_BFX4 U10991 ( .A(n10195), .Z(n10191) );
  HS65_LH_BFX4 U10992 ( .A(n10196), .Z(n10192) );
  HS65_LH_BFX4 U10994 ( .A(n10198), .Z(n10194) );
  HS65_LH_BFX4 U10995 ( .A(n10199), .Z(n10195) );
  HS65_LH_BFX4 U10996 ( .A(n10200), .Z(n10196) );
  HS65_LH_BFX4 U10998 ( .A(n10202), .Z(n10198) );
  HS65_LH_BFX4 U10999 ( .A(n10203), .Z(n10199) );
  HS65_LH_BFX4 U11000 ( .A(n10204), .Z(n10200) );
  HS65_LH_BFX4 U11002 ( .A(n10206), .Z(n10202) );
  HS65_LH_BFX4 U11003 ( .A(n10207), .Z(n10203) );
  HS65_LH_BFX4 U11004 ( .A(n10208), .Z(n10204) );
  HS65_LH_BFX4 U11006 ( .A(n10210), .Z(n10206) );
  HS65_LH_BFX4 U11007 ( .A(n10211), .Z(n10207) );
  HS65_LH_BFX4 U11008 ( .A(n10212), .Z(n10208) );
  HS65_LH_BFX4 U11010 ( .A(n10214), .Z(n10210) );
  HS65_LH_BFX4 U11011 ( .A(n10215), .Z(n10211) );
  HS65_LH_BFX4 U11012 ( .A(n10216), .Z(n10212) );
  HS65_LH_BFX4 U11014 ( .A(n10218), .Z(n10214) );
  HS65_LH_BFX4 U11015 ( .A(n10219), .Z(n10215) );
  HS65_LH_BFX4 U11016 ( .A(n10220), .Z(n10216) );
  HS65_LH_BFX4 U11018 ( .A(n10222), .Z(n10218) );
  HS65_LH_BFX4 U11019 ( .A(n10223), .Z(n10219) );
  HS65_LH_BFX4 U11020 ( .A(n10224), .Z(n10220) );
  HS65_LH_BFX4 U11022 ( .A(n10225), .Z(n10222) );
  HS65_LH_BFX4 U11023 ( .A(n10226), .Z(n10223) );
  HS65_LH_BFX4 U11024 ( .A(n10227), .Z(n10224) );
  HS65_LH_BFX4 U11025 ( .A(n10178), .Z(n10225) );
  HS65_LH_BFX4 U11026 ( .A(n10229), .Z(n10226) );
  HS65_LH_BFX4 U11027 ( .A(n10230), .Z(n10227) );
  HS65_LH_BFX4 U11028 ( .A(n15477), .Z(n10228) );
  HS65_LH_BFX4 U11029 ( .A(n10231), .Z(n10229) );
  HS65_LH_BFX4 U11030 ( .A(n10232), .Z(n10230) );
  HS65_LH_BFX4 U11031 ( .A(n10233), .Z(n10231) );
  HS65_LH_BFX4 U11032 ( .A(n10234), .Z(n10232) );
  HS65_LH_BFX4 U11033 ( .A(n10235), .Z(n10233) );
  HS65_LH_BFX4 U11034 ( .A(n10236), .Z(n10234) );
  HS65_LH_BFX4 U11035 ( .A(n10237), .Z(n10235) );
  HS65_LH_BFX4 U11036 ( .A(n10238), .Z(n10236) );
  HS65_LH_BFX4 U11037 ( .A(n10239), .Z(n10237) );
  HS65_LH_BFX4 U11038 ( .A(n10240), .Z(n10238) );
  HS65_LH_BFX4 U11039 ( .A(\u_DataPath/branch_target_i [2]), .Z(n10239) );
  HS65_LH_BFX4 U11040 ( .A(\u_DataPath/jump_address_i [2]), .Z(n10240) );
  HS65_LH_BFX4 U11041 ( .A(n10242), .Z(n10241) );
  HS65_LH_BFX4 U11042 ( .A(n10243), .Z(n10242) );
  HS65_LH_BFX4 U11043 ( .A(n10244), .Z(n10243) );
  HS65_LH_BFX4 U11044 ( .A(n10753), .Z(n10244) );
  HS65_LH_BFX4 U11045 ( .A(n10246), .Z(n10245) );
  HS65_LH_BFX4 U11046 ( .A(n10247), .Z(n10246) );
  HS65_LH_BFX4 U11047 ( .A(n10248), .Z(n10247) );
  HS65_LH_BFX4 U11048 ( .A(n10249), .Z(n10248) );
  HS65_LH_BFX4 U11049 ( .A(n10250), .Z(n10249) );
  HS65_LH_BFX4 U11050 ( .A(n10251), .Z(n10250) );
  HS65_LH_BFX4 U11051 ( .A(n10252), .Z(n10251) );
  HS65_LH_BFX4 U11052 ( .A(n10253), .Z(n10252) );
  HS65_LH_BFX4 U11053 ( .A(n10254), .Z(n10253) );
  HS65_LH_BFX4 U11054 ( .A(n10255), .Z(n10254) );
  HS65_LH_BFX4 U11055 ( .A(n10256), .Z(n10255) );
  HS65_LH_BFX4 U11056 ( .A(n10257), .Z(n10256) );
  HS65_LH_BFX4 U11057 ( .A(n10258), .Z(n10257) );
  HS65_LH_BFX4 U11058 ( .A(n10259), .Z(n10258) );
  HS65_LH_BFX4 U11059 ( .A(n10260), .Z(n10259) );
  HS65_LH_BFX4 U11060 ( .A(n10261), .Z(n10260) );
  HS65_LH_BFX4 U11061 ( .A(n10262), .Z(n10261) );
  HS65_LH_BFX4 U11062 ( .A(n10263), .Z(n10262) );
  HS65_LH_BFX4 U11063 ( .A(n10264), .Z(n10263) );
  HS65_LH_BFX4 U11064 ( .A(n10265), .Z(n10264) );
  HS65_LH_BFX4 U11065 ( .A(n10266), .Z(n10265) );
  HS65_LH_BFX4 U11066 ( .A(n10267), .Z(n10266) );
  HS65_LH_BFX4 U11067 ( .A(n10268), .Z(n10267) );
  HS65_LH_BFX4 U11068 ( .A(n10269), .Z(n10268) );
  HS65_LH_BFX4 U11069 ( .A(\u_DataPath/u_idexreg/N15 ), .Z(n10269) );
  HS65_LH_BFX4 U11070 ( .A(n10271), .Z(n10270) );
  HS65_LH_BFX4 U11071 ( .A(n10272), .Z(n10271) );
  HS65_LH_BFX4 U11072 ( .A(n10273), .Z(n10272) );
  HS65_LH_BFX4 U11073 ( .A(n10274), .Z(n10273) );
  HS65_LH_BFX4 U11074 ( .A(n10275), .Z(n10274) );
  HS65_LH_BFX4 U11075 ( .A(n10276), .Z(n10275) );
  HS65_LH_BFX4 U11076 ( .A(n10277), .Z(n10276) );
  HS65_LH_BFX4 U11077 ( .A(n10278), .Z(n10277) );
  HS65_LH_BFX4 U11078 ( .A(n10279), .Z(n10278) );
  HS65_LH_BFX4 U11079 ( .A(n10280), .Z(n10279) );
  HS65_LH_BFX4 U11080 ( .A(n10281), .Z(n10280) );
  HS65_LH_BFX4 U11081 ( .A(n10282), .Z(n10281) );
  HS65_LH_BFX4 U11082 ( .A(n10283), .Z(n10282) );
  HS65_LH_BFX4 U11083 ( .A(n10284), .Z(n10283) );
  HS65_LH_BFX4 U11084 ( .A(n10285), .Z(n10284) );
  HS65_LH_BFX4 U11085 ( .A(n10286), .Z(n10285) );
  HS65_LH_BFX4 U11086 ( .A(n10287), .Z(n10286) );
  HS65_LH_BFX4 U11087 ( .A(n10288), .Z(n10287) );
  HS65_LH_BFX4 U11088 ( .A(n10290), .Z(n10288) );
  HS65_LH_BFX4 U11089 ( .A(\u_DataPath/cw_exmem_i [4]), .Z(n10289) );
  HS65_LH_BFX4 U11090 ( .A(n10291), .Z(n10290) );
  HS65_LH_BFX4 U11091 ( .A(n10292), .Z(n10291) );
  HS65_LH_BFX4 U11092 ( .A(n11636), .Z(n10292) );
  HS65_LH_BFX4 U11093 ( .A(n10294), .Z(n10293) );
  HS65_LH_BFX4 U11094 ( .A(n10295), .Z(n10294) );
  HS65_LH_BFX4 U11095 ( .A(n10296), .Z(n10295) );
  HS65_LH_BFX4 U11096 ( .A(n10297), .Z(n10296) );
  HS65_LH_BFX4 U11097 ( .A(n10298), .Z(n10297) );
  HS65_LH_BFX4 U11098 ( .A(n10299), .Z(n10298) );
  HS65_LH_BFX4 U11099 ( .A(n10300), .Z(n10299) );
  HS65_LH_BFX4 U11100 ( .A(n10301), .Z(n10300) );
  HS65_LH_BFX4 U11101 ( .A(n10302), .Z(n10301) );
  HS65_LH_BFX4 U11102 ( .A(n10303), .Z(n10302) );
  HS65_LH_BFX4 U11103 ( .A(n10304), .Z(n10303) );
  HS65_LH_BFX4 U11104 ( .A(n10305), .Z(n10304) );
  HS65_LH_BFX4 U11105 ( .A(n10306), .Z(n10305) );
  HS65_LH_BFX4 U11106 ( .A(n10307), .Z(n10306) );
  HS65_LH_BFX4 U11107 ( .A(n10308), .Z(n10307) );
  HS65_LH_BFX4 U11108 ( .A(n10313), .Z(n10308) );
  HS65_LH_BFX4 U11109 ( .A(\u_DataPath/cw_exmem_i [6]), .Z(n10309) );
  HS65_LH_BFX4 U11110 ( .A(n10309), .Z(n10310) );
  HS65_LH_BFX4 U11111 ( .A(n10310), .Z(n10311) );
  HS65_LH_BFX4 U11112 ( .A(n10311), .Z(n10312) );
  HS65_LH_BFX4 U11113 ( .A(n10314), .Z(n10313) );
  HS65_LH_BFX4 U11114 ( .A(n10315), .Z(n10314) );
  HS65_LH_BFX4 U11115 ( .A(n10482), .Z(n10315) );
  HS65_LH_BFX4 U11116 ( .A(n10317), .Z(n10316) );
  HS65_LH_BFX4 U11117 ( .A(n10318), .Z(n10317) );
  HS65_LH_BFX4 U11118 ( .A(n13646), .Z(n10318) );
  HS65_LH_BFX4 U11119 ( .A(opcode_i[0]), .Z(n10319) );
  HS65_LH_BFX4 U11120 ( .A(n10319), .Z(n10320) );
  HS65_LH_BFX4 U11121 ( .A(n10322), .Z(n10321) );
  HS65_LH_BFX4 U11122 ( .A(n10323), .Z(n10322) );
  HS65_LH_BFX4 U11123 ( .A(n10324), .Z(n10323) );
  HS65_LH_BFX4 U11124 ( .A(n10325), .Z(n10324) );
  HS65_LH_BFX4 U11125 ( .A(n10326), .Z(n10325) );
  HS65_LH_BFX4 U11126 ( .A(n10327), .Z(n10326) );
  HS65_LH_BFX4 U11127 ( .A(n10328), .Z(n10327) );
  HS65_LH_BFX4 U11128 ( .A(n10329), .Z(n10328) );
  HS65_LH_BFX4 U11129 ( .A(n10330), .Z(n10329) );
  HS65_LH_BFX4 U11130 ( .A(n10331), .Z(n10330) );
  HS65_LH_BFX4 U11131 ( .A(n10332), .Z(n10331) );
  HS65_LH_BFX4 U11132 ( .A(n10333), .Z(n10332) );
  HS65_LH_BFX4 U11133 ( .A(n10334), .Z(n10333) );
  HS65_LH_BFX4 U11134 ( .A(n10335), .Z(n10334) );
  HS65_LH_BFX4 U11135 ( .A(n10336), .Z(n10335) );
  HS65_LH_BFX4 U11136 ( .A(n10337), .Z(n10336) );
  HS65_LH_BFX4 U11137 ( .A(n10338), .Z(n10337) );
  HS65_LH_BFX4 U11138 ( .A(n10339), .Z(n10338) );
  HS65_LH_BFX4 U11139 ( .A(n10340), .Z(n10339) );
  HS65_LH_BFX4 U11140 ( .A(n10341), .Z(n10340) );
  HS65_LH_BFX4 U11141 ( .A(n10342), .Z(n10341) );
  HS65_LH_BFX4 U11142 ( .A(n10343), .Z(n10342) );
  HS65_LH_BFX4 U11143 ( .A(n10344), .Z(n10343) );
  HS65_LH_BFX4 U11144 ( .A(n10345), .Z(n10344) );
  HS65_LH_BFX4 U11145 ( .A(\u_DataPath/u_idexreg/N8 ), .Z(n10345) );
  HS65_LH_BFX4 U11146 ( .A(n10347), .Z(n10346) );
  HS65_LH_BFX4 U11147 ( .A(n10348), .Z(n10347) );
  HS65_LH_BFX4 U11148 ( .A(n10349), .Z(n10348) );
  HS65_LH_BFX4 U11149 ( .A(n10350), .Z(n10349) );
  HS65_LH_BFX4 U11150 ( .A(n10351), .Z(n10350) );
  HS65_LH_BFX4 U11151 ( .A(n10352), .Z(n10351) );
  HS65_LH_BFX4 U11152 ( .A(n10353), .Z(n10352) );
  HS65_LH_BFX4 U11153 ( .A(n10354), .Z(n10353) );
  HS65_LH_BFX4 U11154 ( .A(n10355), .Z(n10354) );
  HS65_LH_BFX4 U11155 ( .A(n10356), .Z(n10355) );
  HS65_LH_BFX4 U11156 ( .A(n10357), .Z(n10356) );
  HS65_LH_BFX4 U11157 ( .A(n10358), .Z(n10357) );
  HS65_LH_BFX4 U11158 ( .A(n10359), .Z(n10358) );
  HS65_LH_BFX4 U11159 ( .A(n10360), .Z(n10359) );
  HS65_LH_BFX4 U11160 ( .A(n10361), .Z(n10360) );
  HS65_LH_BFX4 U11161 ( .A(n10362), .Z(n10361) );
  HS65_LH_BFX4 U11162 ( .A(n10363), .Z(n10362) );
  HS65_LH_BFX4 U11163 ( .A(n10364), .Z(n10363) );
  HS65_LH_BFX4 U11164 ( .A(n10365), .Z(n10364) );
  HS65_LH_BFX4 U11165 ( .A(n10366), .Z(n10365) );
  HS65_LH_BFX4 U11166 ( .A(n10367), .Z(n10366) );
  HS65_LH_BFX4 U11167 ( .A(n10368), .Z(n10367) );
  HS65_LH_BFX4 U11168 ( .A(n10369), .Z(n10368) );
  HS65_LH_BFX4 U11169 ( .A(n10370), .Z(n10369) );
  HS65_LH_BFX4 U11170 ( .A(\u_DataPath/cw_exmem_i [1]), .Z(n10370) );
  HS65_LH_BFX4 U11171 ( .A(opcode_i[5]), .Z(n10371) );
  HS65_LH_BFX4 U11173 ( .A(n10382), .Z(n10373) );
  HS65_LH_BFX4 U11176 ( .A(\u_DataPath/cw_to_ex_i [20]), .Z(n10376) );
  HS65_LH_BFX4 U11179 ( .A(n10376), .Z(n10379) );
  HS65_LH_BFX4 U11182 ( .A(n10385), .Z(n10382) );
  HS65_LH_BFX4 U11185 ( .A(n10387), .Z(n10385) );
  HS65_LH_BFX4 U11187 ( .A(n10390), .Z(n10387) );
  HS65_LH_BFX4 U11190 ( .A(n10393), .Z(n10390) );
  HS65_LH_BFX4 U11193 ( .A(n10396), .Z(n10393) );
  HS65_LH_BFX4 U11196 ( .A(n10400), .Z(n10396) );
  HS65_LH_BFX4 U11200 ( .A(n10404), .Z(n10400) );
  HS65_LH_BFX4 U11204 ( .A(n10408), .Z(n10404) );
  HS65_LH_BFX4 U11208 ( .A(n10412), .Z(n10408) );
  HS65_LH_BFX4 U11212 ( .A(n10416), .Z(n10412) );
  HS65_LH_BFX4 U11216 ( .A(n10420), .Z(n10416) );
  HS65_LH_BFX4 U11220 ( .A(n10424), .Z(n10420) );
  HS65_LH_BFX4 U11224 ( .A(n10428), .Z(n10424) );
  HS65_LH_BFX4 U11228 ( .A(n10432), .Z(n10428) );
  HS65_LH_BFX4 U11232 ( .A(n10438), .Z(n10432) );
  HS65_LH_BFX4 U11238 ( .A(n14045), .Z(n10438) );
  HS65_LH_BFX4 U11243 ( .A(opcode_i[1]), .Z(n10443) );
  HS65_LH_BFX4 U11244 ( .A(n10443), .Z(n10444) );
  HS65_LH_BFX4 U11245 ( .A(n10444), .Z(n10445) );
  HS65_LH_BFX4 U11246 ( .A(n10445), .Z(n10446) );
  HS65_LH_BFX4 U11247 ( .A(opcode_i[2]), .Z(n10447) );
  HS65_LH_BFX4 U11248 ( .A(n10447), .Z(n10448) );
  HS65_LH_BFX4 U11249 ( .A(n10448), .Z(n10449) );
  HS65_LH_BFX4 U11250 ( .A(n10449), .Z(n10450) );
  HS65_LH_BFX4 U11251 ( .A(n10454), .Z(n10451) );
  HS65_LH_BFX2 U11252 ( .A(n12485), .Z(n10452) );
  HS65_LH_BFX4 U11253 ( .A(n10451), .Z(n10453) );
  HS65_LH_BFX4 U11254 ( .A(n13652), .Z(n10454) );
  HS65_LH_BFX4 U11256 ( .A(n10459), .Z(n10456) );
  HS65_LH_BFX4 U11257 ( .A(n10460), .Z(n10457) );
  HS65_LH_BFX4 U11259 ( .A(n10462), .Z(n10459) );
  HS65_LH_BFX4 U11260 ( .A(n10463), .Z(n10460) );
  HS65_LH_BFX4 U11262 ( .A(n10465), .Z(n10462) );
  HS65_LH_BFX4 U11263 ( .A(n10466), .Z(n10463) );
  HS65_LH_BFX4 U11265 ( .A(n10468), .Z(n10465) );
  HS65_LH_BFX4 U11266 ( .A(n10469), .Z(n10466) );
  HS65_LH_BFX4 U11268 ( .A(n10472), .Z(n10468) );
  HS65_LH_BFX4 U11269 ( .A(n10471), .Z(n10469) );
  HS65_LH_BFX4 U11271 ( .A(n10474), .Z(n10471) );
  HS65_LH_BFX4 U11272 ( .A(n13613), .Z(n10472) );
  HS65_LH_BFX4 U11274 ( .A(n10476), .Z(n10474) );
  HS65_LH_BFX4 U11276 ( .A(n10478), .Z(n10476) );
  HS65_LH_BFX4 U11278 ( .A(n11622), .Z(n10478) );
  HS65_LH_BFX4 U11280 ( .A(n13591), .Z(n10480) );
  HS65_LH_BFX4 U11281 ( .A(n10101), .Z(n10481) );
  HS65_LH_BFX4 U11282 ( .A(n13528), .Z(n10482) );
  HS65_LH_BFX4 U11283 ( .A(n13527), .Z(n10483) );
  HS65_LH_BFX4 U11285 ( .A(n10486), .Z(n10485) );
  HS65_LH_BFX4 U11286 ( .A(n10488), .Z(n10486) );
  HS65_LH_BFX4 U11288 ( .A(n10490), .Z(n10488) );
  HS65_LH_BFX4 U11290 ( .A(n10492), .Z(n10490) );
  HS65_LH_BFX4 U11292 ( .A(n10494), .Z(n10492) );
  HS65_LH_BFX4 U11294 ( .A(n10496), .Z(n10494) );
  HS65_LH_BFX4 U11296 ( .A(n10498), .Z(n10496) );
  HS65_LH_BFX4 U11298 ( .A(n10500), .Z(n10498) );
  HS65_LH_BFX4 U11300 ( .A(n10502), .Z(n10500) );
  HS65_LH_BFX4 U11302 ( .A(n10504), .Z(n10502) );
  HS65_LH_BFX4 U11304 ( .A(n10506), .Z(n10504) );
  HS65_LH_BFX4 U11306 ( .A(n10508), .Z(n10506) );
  HS65_LH_BFX4 U11308 ( .A(n10510), .Z(n10508) );
  HS65_LH_BFX4 U11310 ( .A(n10512), .Z(n10510) );
  HS65_LH_BFX4 U11312 ( .A(n10514), .Z(n10512) );
  HS65_LH_BFX4 U11314 ( .A(n10516), .Z(n10514) );
  HS65_LH_BFX4 U11316 ( .A(n10518), .Z(n10516) );
  HS65_LH_BFX4 U11318 ( .A(n10519), .Z(n10518) );
  HS65_LH_BFX4 U11319 ( .A(n10520), .Z(n10519) );
  HS65_LH_BFX4 U11320 ( .A(n10521), .Z(n10520) );
  HS65_LH_BFX4 U11321 ( .A(n10522), .Z(n10521) );
  HS65_LH_BFX4 U11322 ( .A(n10523), .Z(n10522) );
  HS65_LH_BFX4 U11323 ( .A(n10524), .Z(n10523) );
  HS65_LH_BFX4 U11324 ( .A(n10525), .Z(n10524) );
  HS65_LH_BFX4 U11325 ( .A(n10526), .Z(n10525) );
  HS65_LH_BFX4 U11326 ( .A(\u_DataPath/cw_to_ex_i [19]), .Z(n10526) );
  HS65_LH_BFX4 U11351 ( .A(n9318), .Z(n10551) );
  HS65_LH_BFX4 U11353 ( .A(\u_DataPath/cw_tomem_i [3]), .Z(n10553) );
  HS65_LH_BFX4 U11354 ( .A(n14073), .Z(n10554) );
  HS65_LH_BFX4 U11355 ( .A(\u_DataPath/cw_tomem_i [7]), .Z(n10555) );
  HS65_LH_BFX4 U11356 ( .A(n14064), .Z(n10556) );
  HS65_LH_BFX4 U11357 ( .A(\u_DataPath/cw_tomem_i [8]), .Z(n10557) );
  HS65_LH_BFX4 U11358 ( .A(n14075), .Z(n10558) );
  HS65_LH_BFX4 U11359 ( .A(n10551), .Z(n10559) );
  HS65_LH_BFX4 U11360 ( .A(n10567), .Z(n10560) );
  HS65_LH_BFX4 U11361 ( .A(n10553), .Z(n10561) );
  HS65_LH_BFX4 U11362 ( .A(n10555), .Z(n10562) );
  HS65_LH_BFX4 U11363 ( .A(n10556), .Z(n10563) );
  HS65_LH_BFX4 U11364 ( .A(n10557), .Z(n10564) );
  HS65_LH_BFX4 U11365 ( .A(n10576), .Z(n10565) );
  HS65_LH_BFX4 U11366 ( .A(n10559), .Z(n10566) );
  HS65_LH_BFX4 U11367 ( .A(n10578), .Z(n10567) );
  HS65_LH_BFX4 U11368 ( .A(n10561), .Z(n10568) );
  HS65_LH_BFX4 U11369 ( .A(n10562), .Z(n10569) );
  HS65_LH_BFX4 U11370 ( .A(n10564), .Z(n10570) );
  HS65_LH_BFX4 U11371 ( .A(n10563), .Z(n10571) );
  HS65_LH_CNIVX3 U11372 ( .A(n10583), .Z(n10572) );
  HS65_LH_CNIVX3 U11373 ( .A(n10572), .Z(n10573) );
  HS65_LH_CNIVX3 U11374 ( .A(n10596), .Z(n10574) );
  HS65_LH_CNIVX3 U11375 ( .A(n10574), .Z(n10575) );
  HS65_LH_BFX4 U11376 ( .A(n10586), .Z(n10576) );
  HS65_LH_BFX4 U11377 ( .A(n10566), .Z(n10577) );
  HS65_LH_BFX4 U11378 ( .A(n10590), .Z(n10578) );
  HS65_LH_BFX4 U11379 ( .A(n10568), .Z(n10579) );
  HS65_LH_BFX4 U11380 ( .A(n10571), .Z(n10580) );
  HS65_LH_BFX4 U11381 ( .A(\u_DataPath/cw_tomem_i [5]), .Z(n10581) );
  HS65_LH_CNIVX3 U11382 ( .A(n10603), .Z(n10582) );
  HS65_LH_CNIVX3 U11383 ( .A(n10582), .Z(n10583) );
  HS65_LH_CNIVX3 U11384 ( .A(n10608), .Z(n10584) );
  HS65_LH_CNIVX3 U11385 ( .A(n10584), .Z(n10585) );
  HS65_LH_BFX4 U11386 ( .A(n10681), .Z(n10586) );
  HS65_LH_BFX4 U11387 ( .A(n10577), .Z(n10587) );
  HS65_LH_CNIVX3 U11388 ( .A(n10599), .Z(n10588) );
  HS65_LH_CNIVX3 U11389 ( .A(n10588), .Z(n10589) );
  HS65_LH_BFX4 U11390 ( .A(n10600), .Z(n10590) );
  HS65_LH_BFX4 U11391 ( .A(n10558), .Z(n10591) );
  HS65_LH_BFX4 U11392 ( .A(n10601), .Z(n10592) );
  HS65_LH_BFX4 U11393 ( .A(n10579), .Z(n10593) );
  HS65_LH_BFX4 U11394 ( .A(n10569), .Z(n10594) );
  HS65_LH_CNIVX3 U11395 ( .A(n10607), .Z(n10595) );
  HS65_LH_CNIVX3 U11396 ( .A(n10595), .Z(n10596) );
  HS65_LH_BFX4 U11397 ( .A(n10587), .Z(n10597) );
  HS65_LH_CNIVX3 U11398 ( .A(n10611), .Z(n10598) );
  HS65_LH_CNIVX3 U11399 ( .A(n10598), .Z(n10599) );
  HS65_LH_BFX4 U11400 ( .A(n10623), .Z(n10600) );
  HS65_LH_BFX4 U11401 ( .A(n10613), .Z(n10601) );
  HS65_LH_BFX4 U11402 ( .A(n10593), .Z(n10602) );
  HS65_LH_BFX4 U11403 ( .A(n10605), .Z(n10603) );
  HS65_LH_CNIVX3 U11404 ( .A(n10616), .Z(n10604) );
  HS65_LH_CNIVX3 U11405 ( .A(n10604), .Z(n10605) );
  HS65_LH_CNIVX3 U11406 ( .A(n10618), .Z(n10606) );
  HS65_LH_CNIVX3 U11407 ( .A(n10606), .Z(n10607) );
  HS65_LH_BFX4 U11408 ( .A(n10619), .Z(n10608) );
  HS65_LH_BFX4 U11409 ( .A(n10597), .Z(n10609) );
  HS65_LH_CNIVX3 U11410 ( .A(n10622), .Z(n10610) );
  HS65_LH_CNIVX3 U11411 ( .A(n10610), .Z(n10611) );
  HS65_LH_BFX4 U11412 ( .A(\u_DataPath/dataOut_exe_i [1]), .Z(n10612) );
  HS65_LH_BFX4 U11413 ( .A(n10624), .Z(n10613) );
  HS65_LH_BFX4 U11414 ( .A(n10602), .Z(n10614) );
  HS65_LH_CNIVX3 U11415 ( .A(n10626), .Z(n10615) );
  HS65_LH_CNIVX3 U11416 ( .A(n10615), .Z(n10616) );
  HS65_LH_CNIVX3 U11417 ( .A(n10628), .Z(n10617) );
  HS65_LH_CNIVX3 U11418 ( .A(n10617), .Z(n10618) );
  HS65_LH_BFX4 U11419 ( .A(n10630), .Z(n10619) );
  HS65_LH_BFX4 U11420 ( .A(n10609), .Z(n10620) );
  HS65_LH_CNIVX3 U11421 ( .A(n10633), .Z(n10621) );
  HS65_LH_CNIVX3 U11422 ( .A(n10621), .Z(n10622) );
  HS65_LH_BFX4 U11423 ( .A(n10645), .Z(n10623) );
  HS65_LH_BFX4 U11424 ( .A(n10635), .Z(n10624) );
  HS65_LH_CNIVX3 U11425 ( .A(n10637), .Z(n10625) );
  HS65_LH_CNIVX3 U11426 ( .A(n10625), .Z(n10626) );
  HS65_LH_CNIVX3 U11427 ( .A(n10639), .Z(n10627) );
  HS65_LH_CNIVX3 U11428 ( .A(n10627), .Z(n10628) );
  HS65_LH_BFX4 U11429 ( .A(n10614), .Z(n10629) );
  HS65_LH_BFX4 U11430 ( .A(n10641), .Z(n10630) );
  HS65_LH_BFX4 U11431 ( .A(n10620), .Z(n10631) );
  HS65_LH_CNIVX3 U11432 ( .A(n10643), .Z(n10632) );
  HS65_LH_CNIVX3 U11433 ( .A(n10632), .Z(n10633) );
  HS65_LH_BFX4 U11434 ( .A(n10612), .Z(n10634) );
  HS65_LH_BFX4 U11435 ( .A(n10646), .Z(n10635) );
  HS65_LH_CNIVX3 U11436 ( .A(n10648), .Z(n10636) );
  HS65_LH_CNIVX3 U11437 ( .A(n10636), .Z(n10637) );
  HS65_LH_CNIVX3 U11438 ( .A(n10650), .Z(n10638) );
  HS65_LH_CNIVX3 U11439 ( .A(n10638), .Z(n10639) );
  HS65_LH_BFX4 U11440 ( .A(n10629), .Z(n10640) );
  HS65_LH_BFX4 U11441 ( .A(n10651), .Z(n10641) );
  HS65_LH_CNIVX3 U11442 ( .A(n10656), .Z(n10642) );
  HS65_LH_CNIVX3 U11443 ( .A(n10642), .Z(n10643) );
  HS65_LH_BFX4 U11444 ( .A(n10631), .Z(n10644) );
  HS65_LH_BFX4 U11445 ( .A(n10668), .Z(n10645) );
  HS65_LH_BFX4 U11446 ( .A(n10659), .Z(n10646) );
  HS65_LH_CNIVX3 U11447 ( .A(n10661), .Z(n10647) );
  HS65_LH_CNIVX3 U11448 ( .A(n10647), .Z(n10648) );
  HS65_LH_CNIVX3 U11449 ( .A(n10663), .Z(n10649) );
  HS65_LH_CNIVX3 U11450 ( .A(n10649), .Z(n10650) );
  HS65_LH_BFX4 U11451 ( .A(n10654), .Z(n10651) );
  HS65_LH_BFX4 U11452 ( .A(n10640), .Z(n10652) );
  HS65_LH_CNIVX3 U11453 ( .A(n10674), .Z(n10653) );
  HS65_LH_CNIVX3 U11454 ( .A(n10653), .Z(n10654) );
  HS65_LH_CNIVX3 U11455 ( .A(n10666), .Z(n10655) );
  HS65_LH_CNIVX3 U11456 ( .A(n10655), .Z(n10656) );
  HS65_LH_BFX4 U11457 ( .A(n10644), .Z(n10657) );
  HS65_LH_BFX4 U11458 ( .A(n10634), .Z(n10658) );
  HS65_LH_BFX4 U11459 ( .A(n10669), .Z(n10659) );
  HS65_LH_CNIVX3 U11460 ( .A(n10671), .Z(n10660) );
  HS65_LH_CNIVX3 U11461 ( .A(n10660), .Z(n10661) );
  HS65_LH_CNIVX3 U11462 ( .A(n10673), .Z(n10662) );
  HS65_LH_CNIVX3 U11463 ( .A(n10662), .Z(n10663) );
  HS65_LH_BFX4 U11464 ( .A(n10652), .Z(n10664) );
  HS65_LH_CNIVX3 U11465 ( .A(n10689), .Z(n10665) );
  HS65_LH_CNIVX3 U11466 ( .A(n10665), .Z(n10666) );
  HS65_LH_BFX4 U11467 ( .A(n10657), .Z(n10667) );
  HS65_LH_BFX4 U11468 ( .A(n10692), .Z(n10668) );
  HS65_LH_BFX4 U11469 ( .A(n10693), .Z(n10669) );
  HS65_LH_CNIVX3 U11470 ( .A(n10685), .Z(n10670) );
  HS65_LH_CNIVX3 U11471 ( .A(n10670), .Z(n10671) );
  HS65_LH_CNIVX3 U11472 ( .A(n10687), .Z(n10672) );
  HS65_LH_CNIVX3 U11473 ( .A(n10672), .Z(n10673) );
  HS65_LH_BFX4 U11474 ( .A(n10698), .Z(n10674) );
  HS65_LH_CNIVX3 U11475 ( .A(n10591), .Z(n10675) );
  HS65_LH_CNIVX3 U11476 ( .A(n10675), .Z(n10676) );
  HS65_LH_CNIVX3 U11477 ( .A(n10700), .Z(n10677) );
  HS65_LH_CNIVX3 U11478 ( .A(n10677), .Z(n10678) );
  HS65_LH_BFX4 U11479 ( .A(n10664), .Z(n10679) );
  HS65_LH_CNIVX3 U11480 ( .A(n15704), .Z(n10680) );
  HS65_LH_CNIVX3 U11481 ( .A(n10680), .Z(n10681) );
  HS65_LH_BFX4 U11482 ( .A(n10667), .Z(n10682) );
  HS65_LH_BFX4 U11483 ( .A(n10658), .Z(n10683) );
  HS65_LH_CNIVX3 U11484 ( .A(n10695), .Z(n10684) );
  HS65_LH_CNIVX3 U11485 ( .A(n10684), .Z(n10685) );
  HS65_LH_CNIVX3 U11486 ( .A(n10697), .Z(n10686) );
  HS65_LH_CNIVX3 U11487 ( .A(n10686), .Z(n10687) );
  HS65_LH_CNIVX3 U11488 ( .A(n9306), .Z(n10688) );
  HS65_LH_CNIVX3 U11489 ( .A(n10688), .Z(n10689) );
  HS65_LH_BFX4 U11490 ( .A(n10679), .Z(n10690) );
  HS65_LH_BFX4 U11491 ( .A(n10682), .Z(n10691) );
  HS65_LH_BFX4 U11492 ( .A(n10683), .Z(n10692) );
  HS65_LH_BFX4 U11493 ( .A(n10711), .Z(n10693) );
  HS65_LH_CNIVX3 U11494 ( .A(n10706), .Z(n10694) );
  HS65_LH_CNIVX3 U11495 ( .A(n10694), .Z(n10695) );
  HS65_LH_CNIVX3 U11496 ( .A(n10708), .Z(n10696) );
  HS65_LH_CNIVX3 U11497 ( .A(n10696), .Z(n10697) );
  HS65_LH_BFX4 U11498 ( .A(n10581), .Z(n10698) );
  HS65_LH_CNIVX3 U11499 ( .A(n10580), .Z(n10699) );
  HS65_LH_CNIVX3 U11500 ( .A(n10699), .Z(n10700) );
  HS65_LH_BFX4 U11501 ( .A(n10691), .Z(n10701) );
  HS65_LH_BFX4 U11502 ( .A(n10690), .Z(n10702) );
  HS65_LH_CNIVX3 U11503 ( .A(n10718), .Z(n10703) );
  HS65_LH_CNIVX3 U11504 ( .A(n10703), .Z(n10704) );
  HS65_LH_CNIVX3 U11505 ( .A(n10714), .Z(n10705) );
  HS65_LH_CNIVX3 U11506 ( .A(n10705), .Z(n10706) );
  HS65_LH_CNIVX3 U11507 ( .A(n10716), .Z(n10707) );
  HS65_LH_CNIVX3 U11508 ( .A(n10707), .Z(n10708) );
  HS65_LH_CNIVX3 U11509 ( .A(n9293), .Z(n10709) );
  HS65_LH_CNIVX3 U11510 ( .A(n10709), .Z(n10710) );
  HS65_LH_BFX4 U11511 ( .A(n10717), .Z(n10711) );
  HS65_LH_BFX4 U11512 ( .A(n10702), .Z(n10712) );
  HS65_LH_CNIVX3 U11513 ( .A(n10723), .Z(n10713) );
  HS65_LH_CNIVX3 U11514 ( .A(n10713), .Z(n10714) );
  HS65_LH_CNIVX3 U11515 ( .A(n10725), .Z(n10715) );
  HS65_LH_CNIVX3 U11516 ( .A(n10715), .Z(n10716) );
  HS65_LH_BFX4 U11517 ( .A(\u_DataPath/cw_tomem_i [6]), .Z(n10717) );
  HS65_LH_BFX4 U11518 ( .A(n10701), .Z(n10718) );
  HS65_LH_BFX4 U11519 ( .A(n10712), .Z(n10719) );
  HS65_LH_CNIVX3 U11520 ( .A(n14047), .Z(n10720) );
  HS65_LH_CNIVX3 U11521 ( .A(n10720), .Z(n10721) );
  HS65_LH_CNIVX3 U11522 ( .A(n10570), .Z(n10722) );
  HS65_LH_CNIVX3 U11523 ( .A(n10722), .Z(n10723) );
  HS65_LH_CNIVX3 U11524 ( .A(n10594), .Z(n10724) );
  HS65_LH_CNIVX3 U11525 ( .A(n10724), .Z(n10725) );
  HS65_LH_BFX4 U11526 ( .A(n10727), .Z(n10726) );
  HS65_LH_BFX4 U11527 ( .A(n10728), .Z(n10727) );
  HS65_LH_BFX4 U11528 ( .A(n10729), .Z(n10728) );
  HS65_LH_BFX4 U11529 ( .A(n10730), .Z(n10729) );
  HS65_LH_BFX4 U11530 ( .A(n10731), .Z(n10730) );
  HS65_LH_BFX4 U11531 ( .A(n10732), .Z(n10731) );
  HS65_LH_BFX4 U11532 ( .A(n10733), .Z(n10732) );
  HS65_LH_BFX4 U11533 ( .A(n10734), .Z(n10733) );
  HS65_LH_BFX4 U11534 ( .A(n10735), .Z(n10734) );
  HS65_LH_BFX4 U11535 ( .A(n10736), .Z(n10735) );
  HS65_LH_BFX4 U11536 ( .A(n10737), .Z(n10736) );
  HS65_LH_BFX4 U11537 ( .A(n10738), .Z(n10737) );
  HS65_LH_BFX4 U11538 ( .A(n10739), .Z(n10738) );
  HS65_LH_BFX4 U11539 ( .A(n10740), .Z(n10739) );
  HS65_LH_BFX4 U11540 ( .A(n10741), .Z(n10740) );
  HS65_LH_BFX4 U11541 ( .A(n10742), .Z(n10741) );
  HS65_LH_BFX4 U11542 ( .A(n10743), .Z(n10742) );
  HS65_LH_BFX4 U11543 ( .A(n10744), .Z(n10743) );
  HS65_LH_BFX4 U11544 ( .A(n10745), .Z(n10744) );
  HS65_LH_BFX4 U11545 ( .A(n10746), .Z(n10745) );
  HS65_LH_BFX4 U11546 ( .A(n10747), .Z(n10746) );
  HS65_LH_BFX4 U11547 ( .A(n10748), .Z(n10747) );
  HS65_LH_BFX4 U11548 ( .A(n14048), .Z(n10748) );
  HS65_LH_BFX4 U11549 ( .A(\u_DataPath/u_idexreg/N20 ), .Z(n10749) );
  HS65_LH_BFX4 U11550 ( .A(n10756), .Z(n10750) );
  HS65_LH_BFX4 U11551 ( .A(n10757), .Z(n10751) );
  HS65_LH_BFX4 U11553 ( .A(n10759), .Z(n10753) );
  HS65_LH_BFX4 U11554 ( .A(n10760), .Z(n10754) );
  HS65_LH_BFX4 U11555 ( .A(n10761), .Z(n10755) );
  HS65_LH_BFX4 U11556 ( .A(n10762), .Z(n10756) );
  HS65_LH_BFX4 U11557 ( .A(n10763), .Z(n10757) );
  HS65_LH_BFX4 U11559 ( .A(n10765), .Z(n10759) );
  HS65_LH_BFX4 U11560 ( .A(n10766), .Z(n10760) );
  HS65_LH_BFX4 U11561 ( .A(n10767), .Z(n10761) );
  HS65_LH_BFX4 U11562 ( .A(n10768), .Z(n10762) );
  HS65_LH_BFX4 U11563 ( .A(n10769), .Z(n10763) );
  HS65_LH_BFX4 U11565 ( .A(n10773), .Z(n10765) );
  HS65_LH_BFX4 U11566 ( .A(n10774), .Z(n10766) );
  HS65_LH_BFX4 U11567 ( .A(n10775), .Z(n10767) );
  HS65_LH_BFX4 U11568 ( .A(n10776), .Z(n10768) );
  HS65_LH_BFX4 U11569 ( .A(n10771), .Z(n10769) );
  HS65_LH_CNIVX3 U11570 ( .A(n10782), .Z(n10770) );
  HS65_LH_CNIVX3 U11571 ( .A(n10770), .Z(n10771) );
  HS65_LH_BFX4 U11573 ( .A(n10778), .Z(n10773) );
  HS65_LH_BFX4 U11574 ( .A(n10779), .Z(n10774) );
  HS65_LH_BFX4 U11575 ( .A(n10780), .Z(n10775) );
  HS65_LH_BFX4 U11576 ( .A(n10781), .Z(n10776) );
  HS65_LH_BFX4 U11578 ( .A(n10786), .Z(n10778) );
  HS65_LH_BFX4 U11579 ( .A(n10787), .Z(n10779) );
  HS65_LH_BFX4 U11580 ( .A(n10788), .Z(n10780) );
  HS65_LH_BFX4 U11581 ( .A(n10789), .Z(n10781) );
  HS65_LH_BFX4 U11582 ( .A(n10784), .Z(n10782) );
  HS65_LH_CNIVX3 U11583 ( .A(n10791), .Z(n10783) );
  HS65_LH_CNIVX3 U11584 ( .A(n10783), .Z(n10784) );
  HS65_LH_BFX4 U11586 ( .A(n10793), .Z(n10786) );
  HS65_LH_BFX4 U11587 ( .A(n10794), .Z(n10787) );
  HS65_LH_BFX4 U11588 ( .A(n10795), .Z(n10788) );
  HS65_LH_BFX4 U11589 ( .A(n10796), .Z(n10789) );
  HS65_LH_CNIVX3 U11590 ( .A(n10798), .Z(n10790) );
  HS65_LH_CNIVX3 U11591 ( .A(n10790), .Z(n10791) );
  HS65_LH_BFX4 U11593 ( .A(n10800), .Z(n10793) );
  HS65_LH_BFX4 U11594 ( .A(n10801), .Z(n10794) );
  HS65_LH_BFX4 U11595 ( .A(n10802), .Z(n10795) );
  HS65_LH_BFX4 U11596 ( .A(n10803), .Z(n10796) );
  HS65_LH_CNIVX3 U11597 ( .A(n10809), .Z(n10797) );
  HS65_LH_CNIVX3 U11598 ( .A(n10797), .Z(n10798) );
  HS65_LH_BFX4 U11600 ( .A(n10805), .Z(n10800) );
  HS65_LH_BFX4 U11601 ( .A(n10806), .Z(n10801) );
  HS65_LH_BFX4 U11602 ( .A(n10807), .Z(n10802) );
  HS65_LH_BFX4 U11603 ( .A(n10808), .Z(n10803) );
  HS65_LH_BFX4 U11605 ( .A(n10813), .Z(n10805) );
  HS65_LH_BFX4 U11606 ( .A(n10814), .Z(n10806) );
  HS65_LH_BFX4 U11607 ( .A(n10815), .Z(n10807) );
  HS65_LH_BFX4 U11608 ( .A(n10816), .Z(n10808) );
  HS65_LH_BFX4 U11609 ( .A(n10811), .Z(n10809) );
  HS65_LH_CNIVX3 U11610 ( .A(n10818), .Z(n10810) );
  HS65_LH_CNIVX3 U11611 ( .A(n10810), .Z(n10811) );
  HS65_LH_BFX4 U11613 ( .A(n10820), .Z(n10813) );
  HS65_LH_BFX4 U11614 ( .A(n10821), .Z(n10814) );
  HS65_LH_BFX4 U11615 ( .A(n10822), .Z(n10815) );
  HS65_LH_BFX4 U11616 ( .A(n10823), .Z(n10816) );
  HS65_LH_CNIVX3 U11617 ( .A(n10825), .Z(n10817) );
  HS65_LH_CNIVX3 U11618 ( .A(n10817), .Z(n10818) );
  HS65_LH_BFX4 U11620 ( .A(n10827), .Z(n10820) );
  HS65_LH_BFX4 U11621 ( .A(n10828), .Z(n10821) );
  HS65_LH_BFX4 U11622 ( .A(n10829), .Z(n10822) );
  HS65_LH_BFX4 U11623 ( .A(n10830), .Z(n10823) );
  HS65_LH_CNIVX3 U11624 ( .A(n10836), .Z(n10824) );
  HS65_LH_CNIVX3 U11625 ( .A(n10824), .Z(n10825) );
  HS65_LH_BFX4 U11627 ( .A(n10832), .Z(n10827) );
  HS65_LH_BFX4 U11628 ( .A(n10833), .Z(n10828) );
  HS65_LH_BFX4 U11629 ( .A(n10834), .Z(n10829) );
  HS65_LH_BFX4 U11630 ( .A(n10835), .Z(n10830) );
  HS65_LH_BFX4 U11632 ( .A(n10840), .Z(n10832) );
  HS65_LH_BFX4 U11633 ( .A(n10841), .Z(n10833) );
  HS65_LH_BFX4 U11634 ( .A(n10842), .Z(n10834) );
  HS65_LH_BFX4 U11635 ( .A(n10843), .Z(n10835) );
  HS65_LH_BFX4 U11636 ( .A(n10838), .Z(n10836) );
  HS65_LH_CNIVX3 U11637 ( .A(n10845), .Z(n10837) );
  HS65_LH_CNIVX3 U11638 ( .A(n10837), .Z(n10838) );
  HS65_LH_BFX4 U11640 ( .A(n10847), .Z(n10840) );
  HS65_LH_BFX4 U11641 ( .A(n10848), .Z(n10841) );
  HS65_LH_BFX4 U11642 ( .A(n10849), .Z(n10842) );
  HS65_LH_BFX4 U11643 ( .A(n10850), .Z(n10843) );
  HS65_LH_CNIVX3 U11644 ( .A(n10856), .Z(n10844) );
  HS65_LH_CNIVX3 U11645 ( .A(n10844), .Z(n10845) );
  HS65_LH_BFX4 U11647 ( .A(n10852), .Z(n10847) );
  HS65_LH_BFX4 U11648 ( .A(n10853), .Z(n10848) );
  HS65_LH_BFX4 U11649 ( .A(n10854), .Z(n10849) );
  HS65_LH_BFX4 U11650 ( .A(n10855), .Z(n10850) );
  HS65_LH_BFX4 U11652 ( .A(n10860), .Z(n10852) );
  HS65_LH_BFX4 U11653 ( .A(n10861), .Z(n10853) );
  HS65_LH_BFX4 U11654 ( .A(n10862), .Z(n10854) );
  HS65_LH_BFX4 U11655 ( .A(n10863), .Z(n10855) );
  HS65_LH_BFX4 U11656 ( .A(n10858), .Z(n10856) );
  HS65_LH_CNIVX3 U11657 ( .A(n10865), .Z(n10857) );
  HS65_LH_CNIVX3 U11658 ( .A(n10857), .Z(n10858) );
  HS65_LH_BFX4 U11660 ( .A(n10867), .Z(n10860) );
  HS65_LH_BFX4 U11661 ( .A(n10868), .Z(n10861) );
  HS65_LH_BFX4 U11662 ( .A(n10869), .Z(n10862) );
  HS65_LH_BFX4 U11663 ( .A(n10870), .Z(n10863) );
  HS65_LH_CNIVX3 U11664 ( .A(n10872), .Z(n10864) );
  HS65_LH_CNIVX3 U11665 ( .A(n10864), .Z(n10865) );
  HS65_LH_BFX4 U11667 ( .A(n10874), .Z(n10867) );
  HS65_LH_BFX4 U11668 ( .A(n10875), .Z(n10868) );
  HS65_LH_BFX4 U11669 ( .A(n14038), .Z(n10869) );
  HS65_LH_BFX4 U11670 ( .A(n10876), .Z(n10870) );
  HS65_LH_CNIVX3 U11671 ( .A(n10879), .Z(n10871) );
  HS65_LH_CNIVX3 U11672 ( .A(n10871), .Z(n10872) );
  HS65_LH_BFX4 U11674 ( .A(n14043), .Z(n10874) );
  HS65_LH_BFX4 U11675 ( .A(n10877), .Z(n10875) );
  HS65_LH_BFX4 U11676 ( .A(n10878), .Z(n10876) );
  HS65_LH_BFX4 U11677 ( .A(n10880), .Z(n10877) );
  HS65_LH_BFX4 U11678 ( .A(n10881), .Z(n10878) );
  HS65_LH_BFX4 U11679 ( .A(n10882), .Z(n10879) );
  HS65_LH_BFX4 U11680 ( .A(n10883), .Z(n10880) );
  HS65_LH_BFX4 U11681 ( .A(n10886), .Z(n10881) );
  HS65_LH_BFX4 U11682 ( .A(n14049), .Z(n10882) );
  HS65_LH_BFX4 U11683 ( .A(n10885), .Z(n10883) );
  HS65_LH_CNIVX3 U11684 ( .A(\u_DataPath/u_execute/link_value_i [1]), .Z(
        n10884) );
  HS65_LH_CNIVX3 U11685 ( .A(n10884), .Z(n10885) );
  HS65_LH_BFX4 U11686 ( .A(n10887), .Z(n10886) );
  HS65_LH_BFX4 U11687 ( .A(n10888), .Z(n10887) );
  HS65_LH_BFX4 U11688 ( .A(\u_DataPath/u_execute/psw_status_i [1]), .Z(n10888)
         );
  HS65_LH_BFX4 U11689 ( .A(n10890), .Z(n10889) );
  HS65_LH_BFX4 U11690 ( .A(n10894), .Z(n10890) );
  HS65_LH_BFX4 U11691 ( .A(\u_DataPath/RFaddr_out_memwb_i [4]), .Z(n10891) );
  HS65_LH_BFX4 U11692 ( .A(n10891), .Z(n10892) );
  HS65_LH_BFX4 U11693 ( .A(n10892), .Z(n10893) );
  HS65_LH_BFX4 U11694 ( .A(n14050), .Z(n10894) );
  HS65_LH_BFX4 U11695 ( .A(n10893), .Z(n10895) );
  HS65_LH_BFX4 U11696 ( .A(n10895), .Z(n10896) );
  HS65_LH_BFX4 U11697 ( .A(n10896), .Z(n10897) );
  HS65_LH_BFX4 U11698 ( .A(n10897), .Z(n10898) );
  HS65_LH_BFX4 U11699 ( .A(n10898), .Z(n10899) );
  HS65_LH_BFX4 U11700 ( .A(n10899), .Z(n10900) );
  HS65_LH_BFX4 U11701 ( .A(n10900), .Z(n10901) );
  HS65_LH_BFX4 U11702 ( .A(n10901), .Z(n10902) );
  HS65_LH_BFX4 U11703 ( .A(n10902), .Z(n10903) );
  HS65_LH_BFX4 U11704 ( .A(n10903), .Z(n10904) );
  HS65_LH_BFX4 U11705 ( .A(n10904), .Z(n10905) );
  HS65_LH_BFX4 U11706 ( .A(n10905), .Z(n10906) );
  HS65_LH_BFX4 U11707 ( .A(n10906), .Z(n10907) );
  HS65_LH_BFX4 U11708 ( .A(n10907), .Z(n10908) );
  HS65_LH_BFX4 U11709 ( .A(n10908), .Z(n10909) );
  HS65_LH_BFX4 U11710 ( .A(n10909), .Z(n10910) );
  HS65_LH_BFX4 U11711 ( .A(n10910), .Z(n10911) );
  HS65_LH_BFX4 U12217 ( .A(n11418), .Z(n11417) );
  HS65_LH_BFX4 U12218 ( .A(n15624), .Z(n11418) );
  HS65_LH_BFX4 U12236 ( .A(n11437), .Z(n11436) );
  HS65_LH_BFX4 U12237 ( .A(n11438), .Z(n11437) );
  HS65_LH_BFX4 U12238 ( .A(n11439), .Z(n11438) );
  HS65_LH_BFX4 U12239 ( .A(n11440), .Z(n11439) );
  HS65_LH_BFX4 U12240 ( .A(n15626), .Z(n11440) );
  HS65_LH_BFX4 U12256 ( .A(n11457), .Z(n11456) );
  HS65_LH_BFX4 U12257 ( .A(n11458), .Z(n11457) );
  HS65_LH_BFX4 U12258 ( .A(n11459), .Z(n11458) );
  HS65_LH_BFX4 U12259 ( .A(n11460), .Z(n11459) );
  HS65_LH_BFX4 U12260 ( .A(n11461), .Z(n11460) );
  HS65_LH_BFX4 U12261 ( .A(n11462), .Z(n11461) );
  HS65_LH_BFX4 U12262 ( .A(n15628), .Z(n11462) );
  HS65_LH_BFX4 U12275 ( .A(n11476), .Z(n11475) );
  HS65_LH_BFX4 U12276 ( .A(n11477), .Z(n11476) );
  HS65_LH_BFX4 U12277 ( .A(n11478), .Z(n11477) );
  HS65_LH_BFX4 U12278 ( .A(n11479), .Z(n11478) );
  HS65_LH_BFX4 U12279 ( .A(n11480), .Z(n11479) );
  HS65_LH_BFX4 U12280 ( .A(n11481), .Z(n11480) );
  HS65_LH_BFX4 U12281 ( .A(n11482), .Z(n11481) );
  HS65_LH_BFX4 U12282 ( .A(n11483), .Z(n11482) );
  HS65_LH_BFX4 U12283 ( .A(n11484), .Z(n11483) );
  HS65_LH_BFX4 U12284 ( .A(n15630), .Z(n11484) );
  HS65_LH_BFX4 U12295 ( .A(n11496), .Z(n11495) );
  HS65_LH_BFX4 U12296 ( .A(n11497), .Z(n11496) );
  HS65_LH_BFX4 U12297 ( .A(n11498), .Z(n11497) );
  HS65_LH_BFX4 U12298 ( .A(n11499), .Z(n11498) );
  HS65_LH_BFX4 U12299 ( .A(n11500), .Z(n11499) );
  HS65_LH_BFX4 U12300 ( .A(n11501), .Z(n11500) );
  HS65_LH_BFX4 U12301 ( .A(n11502), .Z(n11501) );
  HS65_LH_BFX4 U12302 ( .A(n11503), .Z(n11502) );
  HS65_LH_BFX4 U12303 ( .A(n11504), .Z(n11503) );
  HS65_LH_BFX4 U12304 ( .A(n11505), .Z(n11504) );
  HS65_LH_BFX4 U12305 ( .A(n11506), .Z(n11505) );
  HS65_LH_BFX4 U12306 ( .A(n15632), .Z(n11506) );
  HS65_LH_BFX4 U12314 ( .A(n11515), .Z(n11514) );
  HS65_LH_BFX4 U12315 ( .A(n11516), .Z(n11515) );
  HS65_LH_BFX4 U12316 ( .A(n11517), .Z(n11516) );
  HS65_LH_BFX4 U12317 ( .A(n11518), .Z(n11517) );
  HS65_LH_BFX4 U12318 ( .A(n11519), .Z(n11518) );
  HS65_LH_BFX4 U12319 ( .A(n11520), .Z(n11519) );
  HS65_LH_BFX4 U12320 ( .A(n11521), .Z(n11520) );
  HS65_LH_BFX4 U12321 ( .A(n11522), .Z(n11521) );
  HS65_LH_BFX4 U12322 ( .A(n11523), .Z(n11522) );
  HS65_LH_BFX4 U12323 ( .A(n11524), .Z(n11523) );
  HS65_LH_BFX4 U12324 ( .A(n11525), .Z(n11524) );
  HS65_LH_BFX4 U12325 ( .A(n11526), .Z(n11525) );
  HS65_LH_BFX4 U12326 ( .A(n11527), .Z(n11526) );
  HS65_LH_BFX4 U12327 ( .A(n11528), .Z(n11527) );
  HS65_LH_BFX4 U12328 ( .A(n15634), .Z(n11528) );
  HS65_LH_BFX4 U12334 ( .A(n11535), .Z(n11534) );
  HS65_LH_BFX4 U12335 ( .A(n11536), .Z(n11535) );
  HS65_LH_BFX4 U12336 ( .A(n11537), .Z(n11536) );
  HS65_LH_BFX4 U12337 ( .A(n11538), .Z(n11537) );
  HS65_LH_BFX4 U12338 ( .A(n11539), .Z(n11538) );
  HS65_LH_BFX4 U12339 ( .A(n11540), .Z(n11539) );
  HS65_LH_BFX4 U12340 ( .A(n11541), .Z(n11540) );
  HS65_LH_BFX4 U12341 ( .A(n11542), .Z(n11541) );
  HS65_LH_BFX4 U12342 ( .A(n11543), .Z(n11542) );
  HS65_LH_BFX4 U12343 ( .A(n11544), .Z(n11543) );
  HS65_LH_BFX4 U12344 ( .A(n11545), .Z(n11544) );
  HS65_LH_BFX4 U12345 ( .A(n11546), .Z(n11545) );
  HS65_LH_BFX4 U12346 ( .A(n11547), .Z(n11546) );
  HS65_LH_BFX4 U12347 ( .A(n11548), .Z(n11547) );
  HS65_LH_BFX4 U12348 ( .A(n11549), .Z(n11548) );
  HS65_LH_BFX4 U12349 ( .A(n11550), .Z(n11549) );
  HS65_LH_BFX4 U12350 ( .A(n15636), .Z(n11550) );
  HS65_LH_BFX4 U12353 ( .A(n11554), .Z(n11553) );
  HS65_LH_BFX4 U12354 ( .A(n11555), .Z(n11554) );
  HS65_LH_BFX4 U12355 ( .A(n11556), .Z(n11555) );
  HS65_LH_BFX4 U12356 ( .A(n11557), .Z(n11556) );
  HS65_LH_BFX4 U12357 ( .A(n11558), .Z(n11557) );
  HS65_LH_BFX4 U12358 ( .A(n11559), .Z(n11558) );
  HS65_LH_BFX4 U12359 ( .A(n11560), .Z(n11559) );
  HS65_LH_BFX4 U12360 ( .A(n11561), .Z(n11560) );
  HS65_LH_BFX4 U12361 ( .A(n11562), .Z(n11561) );
  HS65_LH_BFX4 U12362 ( .A(n11563), .Z(n11562) );
  HS65_LH_BFX4 U12363 ( .A(n11564), .Z(n11563) );
  HS65_LH_BFX4 U12364 ( .A(n11565), .Z(n11564) );
  HS65_LH_BFX4 U12365 ( .A(n11566), .Z(n11565) );
  HS65_LH_BFX4 U12366 ( .A(n11567), .Z(n11566) );
  HS65_LH_BFX4 U12367 ( .A(n11568), .Z(n11567) );
  HS65_LH_BFX4 U12368 ( .A(n11569), .Z(n11568) );
  HS65_LH_BFX4 U12369 ( .A(n11570), .Z(n11569) );
  HS65_LH_BFX4 U12370 ( .A(n11571), .Z(n11570) );
  HS65_LH_BFX4 U12371 ( .A(n11572), .Z(n11571) );
  HS65_LH_BFX4 U12372 ( .A(n15638), .Z(n11572) );
  HS65_LH_BFX4 U12373 ( .A(n11574), .Z(n11573) );
  HS65_LH_BFX4 U12374 ( .A(n11575), .Z(n11574) );
  HS65_LH_BFX4 U12375 ( .A(n11576), .Z(n11575) );
  HS65_LH_BFX4 U12376 ( .A(n11577), .Z(n11576) );
  HS65_LH_BFX4 U12377 ( .A(n11578), .Z(n11577) );
  HS65_LH_BFX4 U12378 ( .A(n11579), .Z(n11578) );
  HS65_LH_BFX4 U12379 ( .A(n11580), .Z(n11579) );
  HS65_LH_BFX4 U12380 ( .A(n11581), .Z(n11580) );
  HS65_LH_BFX4 U12381 ( .A(n11582), .Z(n11581) );
  HS65_LH_BFX4 U12382 ( .A(n11583), .Z(n11582) );
  HS65_LH_BFX4 U12383 ( .A(n11584), .Z(n11583) );
  HS65_LH_BFX4 U12384 ( .A(n11585), .Z(n11584) );
  HS65_LH_BFX4 U12385 ( .A(n11586), .Z(n11585) );
  HS65_LH_BFX4 U12386 ( .A(n11587), .Z(n11586) );
  HS65_LH_BFX4 U12387 ( .A(n11588), .Z(n11587) );
  HS65_LH_BFX4 U12388 ( .A(n11589), .Z(n11588) );
  HS65_LH_BFX4 U12389 ( .A(n11590), .Z(n11589) );
  HS65_LH_BFX4 U12390 ( .A(n11591), .Z(n11590) );
  HS65_LH_BFX4 U12391 ( .A(n11592), .Z(n11591) );
  HS65_LH_BFX4 U12392 ( .A(n11593), .Z(n11592) );
  HS65_LH_BFX4 U12393 ( .A(n11594), .Z(n11593) );
  HS65_LH_BFX4 U12394 ( .A(n15639), .Z(n11594) );
  HS65_LH_BFX4 U12395 ( .A(n11596), .Z(n11595) );
  HS65_LH_BFX4 U12396 ( .A(n11597), .Z(n11596) );
  HS65_LH_BFX4 U12397 ( .A(n11598), .Z(n11597) );
  HS65_LH_BFX4 U12398 ( .A(n11599), .Z(n11598) );
  HS65_LH_BFX4 U12399 ( .A(n11600), .Z(n11599) );
  HS65_LH_BFX4 U12400 ( .A(n11601), .Z(n11600) );
  HS65_LH_BFX4 U12401 ( .A(n11602), .Z(n11601) );
  HS65_LH_BFX4 U12402 ( .A(n11603), .Z(n11602) );
  HS65_LH_BFX4 U12403 ( .A(n11604), .Z(n11603) );
  HS65_LH_BFX4 U12404 ( .A(n11605), .Z(n11604) );
  HS65_LH_BFX4 U12405 ( .A(n11606), .Z(n11605) );
  HS65_LH_BFX4 U12406 ( .A(n11607), .Z(n11606) );
  HS65_LH_BFX4 U12407 ( .A(n11608), .Z(n11607) );
  HS65_LH_BFX4 U12408 ( .A(n11609), .Z(n11608) );
  HS65_LH_BFX4 U12409 ( .A(n11610), .Z(n11609) );
  HS65_LH_BFX4 U12410 ( .A(n11611), .Z(n11610) );
  HS65_LH_BFX4 U12411 ( .A(n11612), .Z(n11611) );
  HS65_LH_BFX4 U12412 ( .A(n11613), .Z(n11612) );
  HS65_LH_BFX4 U12413 ( .A(n11614), .Z(n11613) );
  HS65_LH_BFX4 U12414 ( .A(n11615), .Z(n11614) );
  HS65_LH_BFX4 U12415 ( .A(n11616), .Z(n11615) );
  HS65_LH_BFX4 U12416 ( .A(n15642), .Z(n11616) );
  HS65_LH_BFX4 U12418 ( .A(\u_DataPath/u_decode_unit/hdu_0/current_state [0]), 
        .Z(n11618) );
  HS65_LH_BFX4 U12419 ( .A(n10481), .Z(n11619) );
  HS65_LH_BFX4 U12420 ( .A(n11626), .Z(n11620) );
  HS65_LH_BFX4 U12422 ( .A(n11630), .Z(n11622) );
  HS65_LH_BFX4 U12424 ( .A(n11618), .Z(n11624) );
  HS65_LH_BFX4 U12425 ( .A(n11619), .Z(n11625) );
  HS65_LH_BFX4 U12426 ( .A(n11634), .Z(n11626) );
  HS65_LH_BFX4 U12428 ( .A(\u_DataPath/u_decode_unit/hdu_0/current_state [1]), 
        .Z(n11628) );
  HS65_LH_CNIVX3 U12429 ( .A(n11638), .Z(n11629) );
  HS65_LH_CNIVX3 U12430 ( .A(n11629), .Z(n11630) );
  HS65_LH_BFX4 U12432 ( .A(n11624), .Z(n11632) );
  HS65_LH_BFX4 U12433 ( .A(n11625), .Z(n11633) );
  HS65_LH_BFX4 U12434 ( .A(n13541), .Z(n11634) );
  HS65_LH_BFX4 U12436 ( .A(n13585), .Z(n11636) );
  HS65_LH_CNIVX3 U12437 ( .A(n13533), .Z(n11637) );
  HS65_LH_CNIVX3 U12438 ( .A(n11637), .Z(n11638) );
  HS65_LH_BFX4 U12440 ( .A(n11632), .Z(n11640) );
  HS65_LH_BFX4 U12441 ( .A(\u_DataPath/immediate_ext_dec_i [4]), .Z(n11641) );
  HS65_LH_BFX4 U12442 ( .A(n11641), .Z(n11642) );
  HS65_LH_BFX4 U12443 ( .A(n11642), .Z(n11643) );
  HS65_LH_BFX4 U12444 ( .A(n13649), .Z(n11644) );
  HS65_LH_BFX4 U12445 ( .A(n11649), .Z(n11645) );
  HS65_LH_BFX4 U12446 ( .A(\u_DataPath/immediate_ext_dec_i [5]), .Z(n11646) );
  HS65_LH_BFX4 U12447 ( .A(n11646), .Z(n11647) );
  HS65_LH_BFX4 U12448 ( .A(n11647), .Z(n11648) );
  HS65_LH_BFX4 U12449 ( .A(n11650), .Z(n11649) );
  HS65_LH_BFX4 U12450 ( .A(n13641), .Z(n11650) );
  HS65_LH_BFX4 U12451 ( .A(n11652), .Z(n11651) );
  HS65_LH_BFX4 U12452 ( .A(n11653), .Z(n11652) );
  HS65_LH_BFX4 U12453 ( .A(n11654), .Z(n11653) );
  HS65_LH_BFX4 U12454 ( .A(n11655), .Z(n11654) );
  HS65_LH_BFX4 U12455 ( .A(n11656), .Z(n11655) );
  HS65_LH_BFX4 U12456 ( .A(n11657), .Z(n11656) );
  HS65_LH_BFX4 U12457 ( .A(n11658), .Z(n11657) );
  HS65_LH_BFX4 U12458 ( .A(n11659), .Z(n11658) );
  HS65_LH_BFX4 U12459 ( .A(n11660), .Z(n11659) );
  HS65_LH_BFX4 U12460 ( .A(n11661), .Z(n11660) );
  HS65_LH_BFX4 U12461 ( .A(n11662), .Z(n11661) );
  HS65_LH_BFX4 U12462 ( .A(n11663), .Z(n11662) );
  HS65_LH_BFX4 U12463 ( .A(n11664), .Z(n11663) );
  HS65_LH_BFX4 U12464 ( .A(n11665), .Z(n11664) );
  HS65_LH_BFX4 U12465 ( .A(n11666), .Z(n11665) );
  HS65_LH_BFX4 U12466 ( .A(n11667), .Z(n11666) );
  HS65_LH_BFX4 U12467 ( .A(n11668), .Z(n11667) );
  HS65_LH_BFX4 U12468 ( .A(n11669), .Z(n11668) );
  HS65_LH_BFX4 U12469 ( .A(n11670), .Z(n11669) );
  HS65_LH_BFX4 U12470 ( .A(n11671), .Z(n11670) );
  HS65_LH_BFX4 U12471 ( .A(n11672), .Z(n11671) );
  HS65_LH_BFX4 U12472 ( .A(n11673), .Z(n11672) );
  HS65_LH_BFX4 U12473 ( .A(n11674), .Z(n11673) );
  HS65_LH_BFX4 U12474 ( .A(\u_DataPath/immediate_ext_dec_i [6]), .Z(n11674) );
  HS65_LH_BFX4 U12475 ( .A(n11676), .Z(n11675) );
  HS65_LH_BFX4 U12476 ( .A(n11677), .Z(n11676) );
  HS65_LH_BFX4 U12477 ( .A(n11678), .Z(n11677) );
  HS65_LH_BFX4 U12478 ( .A(n11679), .Z(n11678) );
  HS65_LH_BFX4 U12479 ( .A(n11680), .Z(n11679) );
  HS65_LH_BFX4 U12480 ( .A(n11681), .Z(n11680) );
  HS65_LH_BFX4 U12481 ( .A(n11682), .Z(n11681) );
  HS65_LH_BFX4 U12482 ( .A(n11683), .Z(n11682) );
  HS65_LH_BFX4 U12483 ( .A(n11684), .Z(n11683) );
  HS65_LH_BFX4 U12484 ( .A(n11685), .Z(n11684) );
  HS65_LH_BFX4 U12485 ( .A(n11686), .Z(n11685) );
  HS65_LH_BFX4 U12486 ( .A(n11687), .Z(n11686) );
  HS65_LH_BFX4 U12487 ( .A(n11688), .Z(n11687) );
  HS65_LH_BFX4 U12488 ( .A(n11689), .Z(n11688) );
  HS65_LH_BFX4 U12489 ( .A(n11690), .Z(n11689) );
  HS65_LH_BFX4 U12490 ( .A(n11691), .Z(n11690) );
  HS65_LH_BFX4 U12491 ( .A(n11692), .Z(n11691) );
  HS65_LH_BFX4 U12492 ( .A(n11693), .Z(n11692) );
  HS65_LH_BFX4 U12493 ( .A(n11694), .Z(n11693) );
  HS65_LH_BFX4 U12494 ( .A(n11695), .Z(n11694) );
  HS65_LH_BFX4 U12495 ( .A(n11696), .Z(n11695) );
  HS65_LH_BFX4 U12496 ( .A(n11697), .Z(n11696) );
  HS65_LH_BFX4 U12497 ( .A(n11698), .Z(n11697) );
  HS65_LH_BFX4 U12498 ( .A(\u_DataPath/immediate_ext_dec_i [7]), .Z(n11698) );
  HS65_LH_BFX4 U12499 ( .A(n11700), .Z(n11699) );
  HS65_LH_BFX4 U12500 ( .A(n11701), .Z(n11700) );
  HS65_LH_BFX4 U12501 ( .A(n11702), .Z(n11701) );
  HS65_LH_BFX4 U12502 ( .A(n11703), .Z(n11702) );
  HS65_LH_BFX4 U12503 ( .A(n11704), .Z(n11703) );
  HS65_LH_BFX4 U12504 ( .A(n11705), .Z(n11704) );
  HS65_LH_BFX4 U12505 ( .A(n11706), .Z(n11705) );
  HS65_LH_BFX4 U12506 ( .A(n11707), .Z(n11706) );
  HS65_LH_BFX4 U12507 ( .A(n11708), .Z(n11707) );
  HS65_LH_BFX4 U12508 ( .A(n11709), .Z(n11708) );
  HS65_LH_BFX4 U12509 ( .A(n11710), .Z(n11709) );
  HS65_LH_BFX4 U12510 ( .A(n11711), .Z(n11710) );
  HS65_LH_BFX4 U12511 ( .A(n11712), .Z(n11711) );
  HS65_LH_BFX4 U12512 ( .A(n11713), .Z(n11712) );
  HS65_LH_BFX4 U12513 ( .A(n11714), .Z(n11713) );
  HS65_LH_BFX4 U12514 ( .A(n11715), .Z(n11714) );
  HS65_LH_BFX4 U12515 ( .A(n11716), .Z(n11715) );
  HS65_LH_BFX4 U12516 ( .A(n11717), .Z(n11716) );
  HS65_LH_BFX4 U12517 ( .A(n11718), .Z(n11717) );
  HS65_LH_BFX4 U12518 ( .A(n11719), .Z(n11718) );
  HS65_LH_BFX4 U12519 ( .A(n11720), .Z(n11719) );
  HS65_LH_BFX4 U12520 ( .A(n11721), .Z(n11720) );
  HS65_LH_BFX4 U12521 ( .A(n11722), .Z(n11721) );
  HS65_LH_BFX4 U12522 ( .A(\u_DataPath/immediate_ext_dec_i [8]), .Z(n11722) );
  HS65_LH_BFX4 U12523 ( .A(n11724), .Z(n11723) );
  HS65_LH_BFX4 U12524 ( .A(n11725), .Z(n11724) );
  HS65_LH_BFX4 U12525 ( .A(n11726), .Z(n11725) );
  HS65_LH_BFX4 U12526 ( .A(n11727), .Z(n11726) );
  HS65_LH_BFX4 U12527 ( .A(n11728), .Z(n11727) );
  HS65_LH_BFX4 U12528 ( .A(n11729), .Z(n11728) );
  HS65_LH_BFX4 U12529 ( .A(n11730), .Z(n11729) );
  HS65_LH_BFX4 U12530 ( .A(n11731), .Z(n11730) );
  HS65_LH_BFX4 U12531 ( .A(n11732), .Z(n11731) );
  HS65_LH_BFX4 U12532 ( .A(n11733), .Z(n11732) );
  HS65_LH_BFX4 U12533 ( .A(n11734), .Z(n11733) );
  HS65_LH_BFX4 U12534 ( .A(n11735), .Z(n11734) );
  HS65_LH_BFX4 U12535 ( .A(n11736), .Z(n11735) );
  HS65_LH_BFX4 U12536 ( .A(n11737), .Z(n11736) );
  HS65_LH_BFX4 U12537 ( .A(n11738), .Z(n11737) );
  HS65_LH_BFX4 U12538 ( .A(n11739), .Z(n11738) );
  HS65_LH_BFX4 U12539 ( .A(n11740), .Z(n11739) );
  HS65_LH_BFX4 U12540 ( .A(n11741), .Z(n11740) );
  HS65_LH_BFX4 U12541 ( .A(n11742), .Z(n11741) );
  HS65_LH_BFX4 U12542 ( .A(n11743), .Z(n11742) );
  HS65_LH_BFX4 U12543 ( .A(n11744), .Z(n11743) );
  HS65_LH_BFX4 U12544 ( .A(n11745), .Z(n11744) );
  HS65_LH_BFX4 U12545 ( .A(n11746), .Z(n11745) );
  HS65_LH_BFX4 U12546 ( .A(\u_DataPath/immediate_ext_dec_i [9]), .Z(n11746) );
  HS65_LH_BFX4 U12547 ( .A(n11748), .Z(n11747) );
  HS65_LH_BFX4 U12548 ( .A(n11749), .Z(n11748) );
  HS65_LH_BFX4 U12549 ( .A(n11750), .Z(n11749) );
  HS65_LH_BFX4 U12550 ( .A(n11751), .Z(n11750) );
  HS65_LH_BFX4 U12551 ( .A(n11752), .Z(n11751) );
  HS65_LH_BFX4 U12552 ( .A(n11753), .Z(n11752) );
  HS65_LH_BFX4 U12553 ( .A(n11754), .Z(n11753) );
  HS65_LH_BFX4 U12554 ( .A(n11755), .Z(n11754) );
  HS65_LH_BFX4 U12555 ( .A(n11756), .Z(n11755) );
  HS65_LH_BFX4 U12556 ( .A(n11757), .Z(n11756) );
  HS65_LH_BFX4 U12557 ( .A(n11758), .Z(n11757) );
  HS65_LH_BFX4 U12558 ( .A(n11759), .Z(n11758) );
  HS65_LH_BFX4 U12559 ( .A(n11760), .Z(n11759) );
  HS65_LH_BFX4 U12560 ( .A(n11761), .Z(n11760) );
  HS65_LH_BFX4 U12561 ( .A(n11762), .Z(n11761) );
  HS65_LH_BFX4 U12562 ( .A(n11763), .Z(n11762) );
  HS65_LH_BFX4 U12563 ( .A(n11764), .Z(n11763) );
  HS65_LH_BFX4 U12564 ( .A(n11765), .Z(n11764) );
  HS65_LH_BFX4 U12565 ( .A(n11766), .Z(n11765) );
  HS65_LH_BFX4 U12566 ( .A(n11767), .Z(n11766) );
  HS65_LH_BFX4 U12567 ( .A(n11768), .Z(n11767) );
  HS65_LH_BFX4 U12568 ( .A(n11769), .Z(n11768) );
  HS65_LH_BFX4 U12569 ( .A(n11770), .Z(n11769) );
  HS65_LH_BFX4 U12570 ( .A(\u_DataPath/immediate_ext_dec_i [10]), .Z(n11770)
         );
  HS65_LH_BFX4 U12571 ( .A(n11772), .Z(n11771) );
  HS65_LH_BFX4 U12572 ( .A(n11773), .Z(n11772) );
  HS65_LH_BFX4 U12573 ( .A(n11774), .Z(n11773) );
  HS65_LH_BFX4 U12574 ( .A(n11775), .Z(n11774) );
  HS65_LH_BFX4 U12575 ( .A(n11776), .Z(n11775) );
  HS65_LH_BFX4 U12576 ( .A(n11777), .Z(n11776) );
  HS65_LH_BFX4 U12577 ( .A(n11778), .Z(n11777) );
  HS65_LH_BFX4 U12578 ( .A(n11779), .Z(n11778) );
  HS65_LH_BFX4 U12579 ( .A(n11780), .Z(n11779) );
  HS65_LH_BFX4 U12580 ( .A(n11781), .Z(n11780) );
  HS65_LH_BFX4 U12581 ( .A(n11782), .Z(n11781) );
  HS65_LH_BFX4 U12582 ( .A(n11783), .Z(n11782) );
  HS65_LH_BFX4 U12583 ( .A(n11784), .Z(n11783) );
  HS65_LH_BFX4 U12584 ( .A(n11785), .Z(n11784) );
  HS65_LH_BFX4 U12585 ( .A(n11786), .Z(n11785) );
  HS65_LH_BFX4 U12586 ( .A(n11787), .Z(n11786) );
  HS65_LH_BFX4 U12587 ( .A(n11788), .Z(n11787) );
  HS65_LH_BFX4 U12588 ( .A(n11789), .Z(n11788) );
  HS65_LH_BFX4 U12589 ( .A(n11790), .Z(n11789) );
  HS65_LH_BFX4 U12590 ( .A(n11791), .Z(n11790) );
  HS65_LH_BFX4 U12591 ( .A(n11792), .Z(n11791) );
  HS65_LH_BFX4 U12592 ( .A(n11793), .Z(n11792) );
  HS65_LH_BFX4 U12593 ( .A(n11794), .Z(n11793) );
  HS65_LH_BFX4 U12594 ( .A(\u_DataPath/immediate_ext_dec_i [11]), .Z(n11794)
         );
  HS65_LH_BFX4 U12595 ( .A(n11796), .Z(n11795) );
  HS65_LH_BFX4 U12596 ( .A(n11797), .Z(n11796) );
  HS65_LH_BFX4 U12597 ( .A(n11798), .Z(n11797) );
  HS65_LH_BFX4 U12598 ( .A(n11799), .Z(n11798) );
  HS65_LH_BFX4 U12599 ( .A(n11800), .Z(n11799) );
  HS65_LH_BFX4 U12600 ( .A(n11801), .Z(n11800) );
  HS65_LH_BFX4 U12601 ( .A(n11802), .Z(n11801) );
  HS65_LH_BFX4 U12602 ( .A(n11803), .Z(n11802) );
  HS65_LH_BFX4 U12603 ( .A(n11804), .Z(n11803) );
  HS65_LH_BFX4 U12604 ( .A(n11805), .Z(n11804) );
  HS65_LH_BFX4 U12605 ( .A(n11806), .Z(n11805) );
  HS65_LH_BFX4 U12606 ( .A(n11807), .Z(n11806) );
  HS65_LH_BFX4 U12607 ( .A(n11808), .Z(n11807) );
  HS65_LH_BFX4 U12608 ( .A(n11809), .Z(n11808) );
  HS65_LH_BFX4 U12609 ( .A(n11810), .Z(n11809) );
  HS65_LH_BFX4 U12610 ( .A(n11811), .Z(n11810) );
  HS65_LH_BFX4 U12611 ( .A(n11812), .Z(n11811) );
  HS65_LH_BFX4 U12612 ( .A(n11813), .Z(n11812) );
  HS65_LH_BFX4 U12613 ( .A(n11814), .Z(n11813) );
  HS65_LH_BFX4 U12614 ( .A(n11815), .Z(n11814) );
  HS65_LH_BFX4 U12615 ( .A(n11816), .Z(n11815) );
  HS65_LH_BFX4 U12616 ( .A(n11817), .Z(n11816) );
  HS65_LH_BFX4 U12617 ( .A(n11818), .Z(n11817) );
  HS65_LH_BFX4 U12618 ( .A(\u_DataPath/immediate_ext_dec_i [12]), .Z(n11818)
         );
  HS65_LH_BFX4 U12619 ( .A(n11820), .Z(n11819) );
  HS65_LH_BFX4 U12620 ( .A(n11821), .Z(n11820) );
  HS65_LH_BFX4 U12621 ( .A(n11822), .Z(n11821) );
  HS65_LH_BFX4 U12622 ( .A(n11823), .Z(n11822) );
  HS65_LH_BFX4 U12623 ( .A(n11824), .Z(n11823) );
  HS65_LH_BFX4 U12624 ( .A(n11825), .Z(n11824) );
  HS65_LH_BFX4 U12625 ( .A(n11826), .Z(n11825) );
  HS65_LH_BFX4 U12626 ( .A(n11827), .Z(n11826) );
  HS65_LH_BFX4 U12627 ( .A(n11828), .Z(n11827) );
  HS65_LH_BFX4 U12628 ( .A(n11829), .Z(n11828) );
  HS65_LH_BFX4 U12629 ( .A(n11830), .Z(n11829) );
  HS65_LH_BFX4 U12630 ( .A(n11831), .Z(n11830) );
  HS65_LH_BFX4 U12631 ( .A(n11832), .Z(n11831) );
  HS65_LH_BFX4 U12632 ( .A(n11833), .Z(n11832) );
  HS65_LH_BFX4 U12633 ( .A(n11834), .Z(n11833) );
  HS65_LH_BFX4 U12634 ( .A(n11835), .Z(n11834) );
  HS65_LH_BFX4 U12635 ( .A(n11836), .Z(n11835) );
  HS65_LH_BFX4 U12636 ( .A(n11837), .Z(n11836) );
  HS65_LH_BFX4 U12637 ( .A(n11838), .Z(n11837) );
  HS65_LH_BFX4 U12638 ( .A(n11839), .Z(n11838) );
  HS65_LH_BFX4 U12639 ( .A(n11840), .Z(n11839) );
  HS65_LH_BFX4 U12640 ( .A(n11841), .Z(n11840) );
  HS65_LH_BFX4 U12641 ( .A(n11842), .Z(n11841) );
  HS65_LH_BFX4 U12642 ( .A(\u_DataPath/immediate_ext_dec_i [14]), .Z(n11842)
         );
  HS65_LH_BFX4 U12643 ( .A(n11844), .Z(n11843) );
  HS65_LH_BFX4 U12644 ( .A(n11845), .Z(n11844) );
  HS65_LH_BFX4 U12645 ( .A(n11846), .Z(n11845) );
  HS65_LH_BFX4 U12646 ( .A(n11847), .Z(n11846) );
  HS65_LH_BFX4 U12647 ( .A(n11848), .Z(n11847) );
  HS65_LH_BFX4 U12648 ( .A(n11849), .Z(n11848) );
  HS65_LH_BFX4 U12649 ( .A(n11850), .Z(n11849) );
  HS65_LH_BFX4 U12650 ( .A(n11851), .Z(n11850) );
  HS65_LH_BFX4 U12651 ( .A(n11852), .Z(n11851) );
  HS65_LH_BFX4 U12652 ( .A(n11853), .Z(n11852) );
  HS65_LH_BFX4 U12653 ( .A(n11854), .Z(n11853) );
  HS65_LH_BFX4 U12654 ( .A(n11855), .Z(n11854) );
  HS65_LH_BFX4 U12655 ( .A(n11856), .Z(n11855) );
  HS65_LH_BFX4 U12656 ( .A(n11857), .Z(n11856) );
  HS65_LH_BFX4 U12657 ( .A(n11858), .Z(n11857) );
  HS65_LH_BFX4 U12658 ( .A(n11859), .Z(n11858) );
  HS65_LH_BFX4 U12659 ( .A(n11860), .Z(n11859) );
  HS65_LH_BFX4 U12660 ( .A(n11861), .Z(n11860) );
  HS65_LH_BFX4 U12661 ( .A(n11862), .Z(n11861) );
  HS65_LH_BFX4 U12662 ( .A(n11863), .Z(n11862) );
  HS65_LH_BFX4 U12663 ( .A(n11864), .Z(n11863) );
  HS65_LH_BFX4 U12664 ( .A(n11865), .Z(n11864) );
  HS65_LH_BFX4 U12665 ( .A(n11866), .Z(n11865) );
  HS65_LH_BFX4 U12666 ( .A(\u_DataPath/immediate_ext_dec_i [13]), .Z(n11866)
         );
  HS65_LH_BFX4 U12667 ( .A(n11868), .Z(n11867) );
  HS65_LH_BFX4 U12668 ( .A(n11878), .Z(n11868) );
  HS65_LH_BFX4 U12669 ( .A(\u_DataPath/jaddr_i [16]), .Z(n11869) );
  HS65_LH_BFX4 U12670 ( .A(n11869), .Z(n11870) );
  HS65_LH_BFX4 U12671 ( .A(n11870), .Z(n11871) );
  HS65_LH_BFX4 U12672 ( .A(n11871), .Z(n11872) );
  HS65_LH_BFX4 U12673 ( .A(n11872), .Z(n11873) );
  HS65_LH_BFX4 U12674 ( .A(n11873), .Z(n11874) );
  HS65_LH_BFX4 U12675 ( .A(n11874), .Z(n11875) );
  HS65_LH_BFX4 U12676 ( .A(n11875), .Z(n11876) );
  HS65_LH_BFX4 U12677 ( .A(n11876), .Z(n11877) );
  HS65_LH_BFX4 U12678 ( .A(n11879), .Z(n11878) );
  HS65_LH_BFX4 U12679 ( .A(n11880), .Z(n11879) );
  HS65_LH_BFX4 U12680 ( .A(n11881), .Z(n11880) );
  HS65_LH_BFX4 U12681 ( .A(n11882), .Z(n11881) );
  HS65_LH_BFX4 U12682 ( .A(n11883), .Z(n11882) );
  HS65_LH_BFX4 U12683 ( .A(n11884), .Z(n11883) );
  HS65_LH_BFX4 U12684 ( .A(n11885), .Z(n11884) );
  HS65_LH_BFX4 U12685 ( .A(n11886), .Z(n11885) );
  HS65_LH_BFX4 U12686 ( .A(n11887), .Z(n11886) );
  HS65_LH_BFX4 U12687 ( .A(n11888), .Z(n11887) );
  HS65_LH_BFX4 U12688 ( .A(n14051), .Z(n11888) );
  HS65_LH_BFX4 U12689 ( .A(n11890), .Z(n11889) );
  HS65_LH_BFX4 U12690 ( .A(n11891), .Z(n11890) );
  HS65_LH_BFX4 U12691 ( .A(n11892), .Z(n11891) );
  HS65_LH_BFX4 U12692 ( .A(n11893), .Z(n11892) );
  HS65_LH_BFX4 U12693 ( .A(n11894), .Z(n11893) );
  HS65_LH_BFX4 U12694 ( .A(n11895), .Z(n11894) );
  HS65_LH_BFX4 U12695 ( .A(n11896), .Z(n11895) );
  HS65_LH_BFX4 U12696 ( .A(n11897), .Z(n11896) );
  HS65_LH_BFX4 U12697 ( .A(n11898), .Z(n11897) );
  HS65_LH_BFX4 U12698 ( .A(n11899), .Z(n11898) );
  HS65_LH_BFX4 U12699 ( .A(n11900), .Z(n11899) );
  HS65_LH_BFX4 U12700 ( .A(n11901), .Z(n11900) );
  HS65_LH_BFX4 U12701 ( .A(n11902), .Z(n11901) );
  HS65_LH_BFX4 U12702 ( .A(n11903), .Z(n11902) );
  HS65_LH_BFX4 U12703 ( .A(n11904), .Z(n11903) );
  HS65_LH_BFX4 U12704 ( .A(n11905), .Z(n11904) );
  HS65_LH_BFX4 U12705 ( .A(n11906), .Z(n11905) );
  HS65_LH_BFX4 U12706 ( .A(n11907), .Z(n11906) );
  HS65_LH_BFX4 U12707 ( .A(n11908), .Z(n11907) );
  HS65_LH_BFX4 U12708 ( .A(n11909), .Z(n11908) );
  HS65_LH_BFX4 U12709 ( .A(n11910), .Z(n11909) );
  HS65_LH_BFX4 U12710 ( .A(n11911), .Z(n11910) );
  HS65_LH_BFX4 U12711 ( .A(n11912), .Z(n11911) );
  HS65_LH_BFX4 U12712 ( .A(\u_DataPath/immediate_ext_dec_i [15]), .Z(n11912)
         );
  HS65_LH_BFX4 U12713 ( .A(n13885), .Z(n11913) );
  HS65_LH_BFX4 U12714 ( .A(\u_DataPath/immediate_ext_dec_i [1]), .Z(n11914) );
  HS65_LH_BFX4 U12715 ( .A(n11914), .Z(n11915) );
  HS65_LH_BFX4 U12716 ( .A(n13887), .Z(n11916) );
  HS65_LH_BFX4 U12717 ( .A(\u_DataPath/immediate_ext_dec_i [0]), .Z(n11917) );
  HS65_LH_BFX4 U12718 ( .A(n11917), .Z(n11918) );
  HS65_LH_BFX4 U12719 ( .A(n11918), .Z(n11919) );
  HS65_LH_BFX4 U12720 ( .A(n17227), .Z(n11920) );
  HS65_LH_BFX4 U12721 ( .A(n11923), .Z(n11921) );
  HS65_LH_BFX4 U12723 ( .A(n11925), .Z(n11923) );
  HS65_LH_BFX4 U12725 ( .A(n11927), .Z(n11925) );
  HS65_LH_BFX4 U12727 ( .A(n11929), .Z(n11927) );
  HS65_LH_BFX4 U12729 ( .A(n11931), .Z(n11929) );
  HS65_LH_BFX4 U12731 ( .A(n11933), .Z(n11931) );
  HS65_LH_BFX4 U12733 ( .A(n11935), .Z(n11933) );
  HS65_LH_BFX4 U12734 ( .A(n11936), .Z(n11934) );
  HS65_LH_BFX4 U12735 ( .A(n11937), .Z(n11935) );
  HS65_LH_BFX4 U12736 ( .A(n11938), .Z(n11936) );
  HS65_LH_BFX4 U12737 ( .A(n11939), .Z(n11937) );
  HS65_LH_BFX4 U12738 ( .A(n11940), .Z(n11938) );
  HS65_LH_BFX4 U12739 ( .A(n11941), .Z(n11939) );
  HS65_LH_BFX4 U12740 ( .A(n11942), .Z(n11940) );
  HS65_LH_BFX4 U12741 ( .A(n11943), .Z(n11941) );
  HS65_LH_BFX4 U12742 ( .A(n11944), .Z(n11942) );
  HS65_LH_BFX4 U12743 ( .A(n11945), .Z(n11943) );
  HS65_LH_BFX4 U12744 ( .A(n11946), .Z(n11944) );
  HS65_LH_BFX4 U12745 ( .A(n11947), .Z(n11945) );
  HS65_LH_BFX4 U12746 ( .A(n11948), .Z(n11946) );
  HS65_LH_BFX4 U12747 ( .A(n11949), .Z(n11947) );
  HS65_LH_BFX4 U12748 ( .A(n11950), .Z(n11948) );
  HS65_LH_BFX4 U12749 ( .A(n11951), .Z(n11949) );
  HS65_LH_BFX4 U12750 ( .A(n11952), .Z(n11950) );
  HS65_LH_BFX4 U12751 ( .A(n11953), .Z(n11951) );
  HS65_LH_BFX4 U12752 ( .A(n11954), .Z(n11952) );
  HS65_LH_BFX4 U12753 ( .A(n11955), .Z(n11953) );
  HS65_LH_BFX4 U12754 ( .A(n11956), .Z(n11954) );
  HS65_LH_BFX4 U12755 ( .A(n11957), .Z(n11955) );
  HS65_LH_BFX4 U12756 ( .A(n11958), .Z(n11956) );
  HS65_LH_BFX4 U12757 ( .A(n11959), .Z(n11957) );
  HS65_LH_BFX4 U12758 ( .A(n11960), .Z(n11958) );
  HS65_LH_BFX4 U12759 ( .A(n11961), .Z(n11959) );
  HS65_LH_BFX4 U12760 ( .A(n15454), .Z(n11960) );
  HS65_LH_BFX4 U12761 ( .A(n11962), .Z(n11961) );
  HS65_LH_BFX4 U12762 ( .A(n11963), .Z(n11962) );
  HS65_LH_BFX4 U12763 ( .A(n11964), .Z(n11963) );
  HS65_LH_BFX4 U12764 ( .A(\u_DataPath/pc4_to_idexreg_i [19]), .Z(n11964) );
  HS65_LH_BFX4 U12766 ( .A(n11968), .Z(n11966) );
  HS65_LH_BFX4 U12768 ( .A(n11970), .Z(n11968) );
  HS65_LH_BFX4 U12770 ( .A(n11972), .Z(n11970) );
  HS65_LH_BFX4 U12772 ( .A(n11974), .Z(n11972) );
  HS65_LH_BFX4 U12774 ( .A(n11976), .Z(n11974) );
  HS65_LH_BFX4 U12776 ( .A(n11978), .Z(n11976) );
  HS65_LH_BFX4 U12778 ( .A(n11980), .Z(n11978) );
  HS65_LH_BFX4 U12780 ( .A(n11982), .Z(n11980) );
  HS65_LH_BFX4 U12782 ( .A(n11984), .Z(n11982) );
  HS65_LH_BFX4 U12784 ( .A(n11986), .Z(n11984) );
  HS65_LH_BFX4 U12786 ( .A(n11988), .Z(n11986) );
  HS65_LH_BFX4 U12787 ( .A(n11989), .Z(n11987) );
  HS65_LH_BFX4 U12788 ( .A(n11990), .Z(n11988) );
  HS65_LH_BFX4 U12789 ( .A(n11991), .Z(n11989) );
  HS65_LH_BFX4 U12790 ( .A(n11992), .Z(n11990) );
  HS65_LH_BFX4 U12791 ( .A(n11993), .Z(n11991) );
  HS65_LH_BFX4 U12792 ( .A(n11994), .Z(n11992) );
  HS65_LH_BFX4 U12793 ( .A(n11995), .Z(n11993) );
  HS65_LH_BFX4 U12794 ( .A(n11996), .Z(n11994) );
  HS65_LH_BFX4 U12795 ( .A(n11997), .Z(n11995) );
  HS65_LH_BFX4 U12796 ( .A(n11998), .Z(n11996) );
  HS65_LH_BFX4 U12797 ( .A(n11999), .Z(n11997) );
  HS65_LH_BFX4 U12798 ( .A(n12000), .Z(n11998) );
  HS65_LH_BFX4 U12799 ( .A(n12001), .Z(n11999) );
  HS65_LH_BFX4 U12800 ( .A(n12002), .Z(n12000) );
  HS65_LH_BFX4 U12801 ( .A(n12003), .Z(n12001) );
  HS65_LH_BFX4 U12802 ( .A(n12004), .Z(n12002) );
  HS65_LH_BFX4 U12803 ( .A(n12005), .Z(n12003) );
  HS65_LH_BFX4 U12804 ( .A(n12006), .Z(n12004) );
  HS65_LH_BFX4 U12805 ( .A(n14095), .Z(n12005) );
  HS65_LH_BFX4 U12806 ( .A(n12007), .Z(n12006) );
  HS65_LH_BFX4 U12807 ( .A(n12008), .Z(n12007) );
  HS65_LH_BFX4 U12808 ( .A(n12009), .Z(n12008) );
  HS65_LH_BFX4 U12809 ( .A(\u_DataPath/pc4_to_idexreg_i [20]), .Z(n12009) );
  HS65_LH_BFX4 U12810 ( .A(n17225), .Z(n12010) );
  HS65_LH_BFX4 U12811 ( .A(n12013), .Z(n12011) );
  HS65_LH_BFX4 U12813 ( .A(n12015), .Z(n12013) );
  HS65_LH_BFX4 U12815 ( .A(n12017), .Z(n12015) );
  HS65_LH_BFX4 U12817 ( .A(n12019), .Z(n12017) );
  HS65_LH_BFX4 U12819 ( .A(n12021), .Z(n12019) );
  HS65_LH_BFX4 U12821 ( .A(n12023), .Z(n12021) );
  HS65_LH_BFX4 U12823 ( .A(n12025), .Z(n12023) );
  HS65_LH_BFX4 U12825 ( .A(n12027), .Z(n12025) );
  HS65_LH_BFX4 U12827 ( .A(n12029), .Z(n12027) );
  HS65_LH_BFX4 U12829 ( .A(n12031), .Z(n12029) );
  HS65_LH_BFX4 U12831 ( .A(n12033), .Z(n12031) );
  HS65_LH_BFX4 U12833 ( .A(n12035), .Z(n12033) );
  HS65_LH_BFX4 U12835 ( .A(n12037), .Z(n12035) );
  HS65_LH_BFX4 U12836 ( .A(n12038), .Z(n12036) );
  HS65_LH_BFX4 U12837 ( .A(n12039), .Z(n12037) );
  HS65_LH_BFX4 U12838 ( .A(n12040), .Z(n12038) );
  HS65_LH_BFX4 U12839 ( .A(n12041), .Z(n12039) );
  HS65_LH_BFX4 U12840 ( .A(n12042), .Z(n12040) );
  HS65_LH_BFX4 U12841 ( .A(n12043), .Z(n12041) );
  HS65_LH_BFX4 U12842 ( .A(n12044), .Z(n12042) );
  HS65_LH_BFX4 U12843 ( .A(n12045), .Z(n12043) );
  HS65_LH_BFX4 U12844 ( .A(n12046), .Z(n12044) );
  HS65_LH_BFX4 U12845 ( .A(n12047), .Z(n12045) );
  HS65_LH_BFX4 U12846 ( .A(n12048), .Z(n12046) );
  HS65_LH_BFX4 U12847 ( .A(n12049), .Z(n12047) );
  HS65_LH_BFX4 U12848 ( .A(n12050), .Z(n12048) );
  HS65_LH_BFX4 U12849 ( .A(n12051), .Z(n12049) );
  HS65_LH_BFX4 U12850 ( .A(n15457), .Z(n12050) );
  HS65_LH_BFX4 U12851 ( .A(n12052), .Z(n12051) );
  HS65_LH_BFX4 U12852 ( .A(n12053), .Z(n12052) );
  HS65_LH_BFX4 U12853 ( .A(n12054), .Z(n12053) );
  HS65_LH_BFX4 U12854 ( .A(\u_DataPath/pc4_to_idexreg_i [21]), .Z(n12054) );
  HS65_LH_BFX4 U12856 ( .A(n12058), .Z(n12056) );
  HS65_LH_BFX4 U12858 ( .A(n12060), .Z(n12058) );
  HS65_LH_BFX4 U12860 ( .A(n12062), .Z(n12060) );
  HS65_LH_BFX4 U12862 ( .A(n12064), .Z(n12062) );
  HS65_LH_BFX4 U12864 ( .A(n12066), .Z(n12064) );
  HS65_LH_BFX4 U12866 ( .A(n12068), .Z(n12066) );
  HS65_LH_BFX4 U12868 ( .A(n12070), .Z(n12068) );
  HS65_LH_BFX4 U12870 ( .A(n12072), .Z(n12070) );
  HS65_LH_BFX4 U12872 ( .A(n12074), .Z(n12072) );
  HS65_LH_BFX4 U12874 ( .A(n12076), .Z(n12074) );
  HS65_LH_BFX4 U12876 ( .A(n12078), .Z(n12076) );
  HS65_LH_BFX4 U12878 ( .A(n12080), .Z(n12078) );
  HS65_LH_BFX4 U12880 ( .A(n12082), .Z(n12080) );
  HS65_LH_BFX4 U12882 ( .A(n12084), .Z(n12082) );
  HS65_LH_BFX4 U12884 ( .A(n12086), .Z(n12084) );
  HS65_LH_BFX4 U12886 ( .A(n12088), .Z(n12086) );
  HS65_LH_BFX4 U12887 ( .A(n12089), .Z(n12087) );
  HS65_LH_BFX4 U12888 ( .A(n12090), .Z(n12088) );
  HS65_LH_BFX4 U12889 ( .A(n12091), .Z(n12089) );
  HS65_LH_BFX4 U12890 ( .A(n12092), .Z(n12090) );
  HS65_LH_BFX4 U12891 ( .A(n12093), .Z(n12091) );
  HS65_LH_BFX4 U12892 ( .A(n12094), .Z(n12092) );
  HS65_LH_BFX4 U12893 ( .A(n12095), .Z(n12093) );
  HS65_LH_BFX4 U12894 ( .A(n12096), .Z(n12094) );
  HS65_LH_BFX4 U12895 ( .A(n14097), .Z(n12095) );
  HS65_LH_BFX4 U12896 ( .A(n12097), .Z(n12096) );
  HS65_LH_BFX4 U12897 ( .A(n12098), .Z(n12097) );
  HS65_LH_BFX4 U12898 ( .A(n12099), .Z(n12098) );
  HS65_LH_BFX4 U12899 ( .A(\u_DataPath/pc4_to_idexreg_i [22]), .Z(n12099) );
  HS65_LH_BFX4 U12900 ( .A(n17223), .Z(n12100) );
  HS65_LH_BFX4 U12901 ( .A(n12103), .Z(n12101) );
  HS65_LH_BFX4 U12903 ( .A(n12105), .Z(n12103) );
  HS65_LH_BFX4 U12905 ( .A(n12107), .Z(n12105) );
  HS65_LH_BFX4 U12907 ( .A(n12109), .Z(n12107) );
  HS65_LH_BFX4 U12909 ( .A(n12111), .Z(n12109) );
  HS65_LH_BFX4 U12911 ( .A(n12113), .Z(n12111) );
  HS65_LH_BFX4 U12913 ( .A(n12115), .Z(n12113) );
  HS65_LH_BFX4 U12915 ( .A(n12117), .Z(n12115) );
  HS65_LH_BFX4 U12917 ( .A(n12119), .Z(n12117) );
  HS65_LH_BFX4 U12919 ( .A(n12121), .Z(n12119) );
  HS65_LH_BFX4 U12921 ( .A(n12123), .Z(n12121) );
  HS65_LH_BFX4 U12923 ( .A(n12125), .Z(n12123) );
  HS65_LH_BFX4 U12925 ( .A(n12127), .Z(n12125) );
  HS65_LH_BFX4 U12927 ( .A(n12129), .Z(n12127) );
  HS65_LH_BFX4 U12929 ( .A(n12131), .Z(n12129) );
  HS65_LH_BFX4 U12931 ( .A(n12133), .Z(n12131) );
  HS65_LH_BFX4 U12933 ( .A(n12135), .Z(n12133) );
  HS65_LH_BFX4 U12935 ( .A(n12137), .Z(n12135) );
  HS65_LH_BFX4 U12937 ( .A(n12139), .Z(n12137) );
  HS65_LH_BFX4 U12938 ( .A(n12140), .Z(n12138) );
  HS65_LH_BFX4 U12939 ( .A(n12141), .Z(n12139) );
  HS65_LH_BFX4 U12940 ( .A(n15460), .Z(n12140) );
  HS65_LH_BFX4 U12941 ( .A(n12142), .Z(n12141) );
  HS65_LH_BFX4 U12942 ( .A(n12143), .Z(n12142) );
  HS65_LH_BFX4 U12943 ( .A(n12144), .Z(n12143) );
  HS65_LH_BFX4 U12944 ( .A(\u_DataPath/pc4_to_idexreg_i [23]), .Z(n12144) );
  HS65_LH_BFX4 U12946 ( .A(n12148), .Z(n12146) );
  HS65_LH_BFX4 U12948 ( .A(n12150), .Z(n12148) );
  HS65_LH_BFX4 U12950 ( .A(n12152), .Z(n12150) );
  HS65_LH_BFX4 U12952 ( .A(n12154), .Z(n12152) );
  HS65_LH_BFX4 U12954 ( .A(n12156), .Z(n12154) );
  HS65_LH_BFX4 U12956 ( .A(n12158), .Z(n12156) );
  HS65_LH_BFX4 U12958 ( .A(n12160), .Z(n12158) );
  HS65_LH_BFX4 U12960 ( .A(n12162), .Z(n12160) );
  HS65_LH_BFX4 U12962 ( .A(n12164), .Z(n12162) );
  HS65_LH_BFX4 U12964 ( .A(n12166), .Z(n12164) );
  HS65_LH_BFX4 U12966 ( .A(n12168), .Z(n12166) );
  HS65_LH_BFX4 U12968 ( .A(n12170), .Z(n12168) );
  HS65_LH_BFX4 U12970 ( .A(n12172), .Z(n12170) );
  HS65_LH_BFX4 U12972 ( .A(n12174), .Z(n12172) );
  HS65_LH_BFX4 U12974 ( .A(n12176), .Z(n12174) );
  HS65_LH_BFX4 U12976 ( .A(n12178), .Z(n12176) );
  HS65_LH_BFX4 U12978 ( .A(n12180), .Z(n12178) );
  HS65_LH_BFX4 U12980 ( .A(n12182), .Z(n12180) );
  HS65_LH_BFX4 U12982 ( .A(n12184), .Z(n12182) );
  HS65_LH_BFX4 U12984 ( .A(n12186), .Z(n12184) );
  HS65_LH_BFX4 U12986 ( .A(n12187), .Z(n12186) );
  HS65_LH_BFX4 U12987 ( .A(n12188), .Z(n12187) );
  HS65_LH_BFX4 U12988 ( .A(n12189), .Z(n12188) );
  HS65_LH_BFX4 U12989 ( .A(\u_DataPath/pc4_to_idexreg_i [24]), .Z(n12189) );
  HS65_LH_BFX4 U12990 ( .A(n17221), .Z(n12190) );
  HS65_LH_BFX4 U12991 ( .A(n12193), .Z(n12191) );
  HS65_LH_BFX4 U12993 ( .A(n12195), .Z(n12193) );
  HS65_LH_BFX4 U12995 ( .A(n12197), .Z(n12195) );
  HS65_LH_BFX4 U12997 ( .A(n12199), .Z(n12197) );
  HS65_LH_BFX4 U12999 ( .A(n12201), .Z(n12199) );
  HS65_LH_BFX4 U13001 ( .A(n12203), .Z(n12201) );
  HS65_LH_BFX4 U13003 ( .A(n12205), .Z(n12203) );
  HS65_LH_BFX4 U13005 ( .A(n12207), .Z(n12205) );
  HS65_LH_BFX4 U13007 ( .A(n12209), .Z(n12207) );
  HS65_LH_BFX4 U13009 ( .A(n12211), .Z(n12209) );
  HS65_LH_BFX4 U13011 ( .A(n12213), .Z(n12211) );
  HS65_LH_BFX4 U13013 ( .A(n12215), .Z(n12213) );
  HS65_LH_BFX4 U13015 ( .A(n12217), .Z(n12215) );
  HS65_LH_BFX4 U13017 ( .A(n12219), .Z(n12217) );
  HS65_LH_BFX4 U13019 ( .A(n12221), .Z(n12219) );
  HS65_LH_BFX4 U13021 ( .A(n12223), .Z(n12221) );
  HS65_LH_BFX4 U13023 ( .A(n12225), .Z(n12223) );
  HS65_LH_BFX4 U13025 ( .A(n12227), .Z(n12225) );
  HS65_LH_BFX4 U13027 ( .A(n12229), .Z(n12227) );
  HS65_LH_BFX4 U13029 ( .A(n12231), .Z(n12229) );
  HS65_LH_BFX4 U13031 ( .A(n12232), .Z(n12231) );
  HS65_LH_BFX4 U13032 ( .A(n12233), .Z(n12232) );
  HS65_LH_BFX4 U13033 ( .A(n12234), .Z(n12233) );
  HS65_LH_BFX4 U13034 ( .A(\u_DataPath/pc4_to_idexreg_i [25]), .Z(n12234) );
  HS65_LH_BFX4 U13036 ( .A(n12238), .Z(n12236) );
  HS65_LH_BFX4 U13038 ( .A(n12240), .Z(n12238) );
  HS65_LH_BFX4 U13040 ( .A(n12242), .Z(n12240) );
  HS65_LH_BFX4 U13042 ( .A(n12244), .Z(n12242) );
  HS65_LH_BFX4 U13044 ( .A(n12246), .Z(n12244) );
  HS65_LH_BFX4 U13046 ( .A(n12248), .Z(n12246) );
  HS65_LH_BFX4 U13048 ( .A(n12250), .Z(n12248) );
  HS65_LH_BFX4 U13050 ( .A(n12252), .Z(n12250) );
  HS65_LH_BFX4 U13052 ( .A(n12254), .Z(n12252) );
  HS65_LH_BFX4 U13054 ( .A(n12256), .Z(n12254) );
  HS65_LH_BFX4 U13056 ( .A(n12258), .Z(n12256) );
  HS65_LH_BFX4 U13058 ( .A(n12260), .Z(n12258) );
  HS65_LH_BFX4 U13060 ( .A(n12262), .Z(n12260) );
  HS65_LH_BFX4 U13062 ( .A(n12264), .Z(n12262) );
  HS65_LH_BFX4 U13064 ( .A(n12266), .Z(n12264) );
  HS65_LH_BFX4 U13066 ( .A(n12268), .Z(n12266) );
  HS65_LH_BFX4 U13068 ( .A(n12270), .Z(n12268) );
  HS65_LH_BFX4 U13070 ( .A(n12272), .Z(n12270) );
  HS65_LH_BFX4 U13072 ( .A(n12274), .Z(n12272) );
  HS65_LH_BFX4 U13074 ( .A(n12276), .Z(n12274) );
  HS65_LH_BFX4 U13076 ( .A(n12277), .Z(n12276) );
  HS65_LH_BFX4 U13077 ( .A(n12278), .Z(n12277) );
  HS65_LH_BFX4 U13078 ( .A(n12279), .Z(n12278) );
  HS65_LH_BFX4 U13079 ( .A(\u_DataPath/pc4_to_idexreg_i [26]), .Z(n12279) );
  HS65_LH_BFX4 U13080 ( .A(n12281), .Z(n12280) );
  HS65_LH_BFX4 U13081 ( .A(n12291), .Z(n12281) );
  HS65_LH_BFX4 U13082 ( .A(\u_DataPath/jaddr_i [17]), .Z(n12282) );
  HS65_LH_BFX4 U13083 ( .A(n12282), .Z(n12283) );
  HS65_LH_BFX4 U13084 ( .A(n12283), .Z(n12284) );
  HS65_LH_BFX4 U13085 ( .A(n12284), .Z(n12285) );
  HS65_LH_BFX4 U13086 ( .A(n12285), .Z(n12286) );
  HS65_LH_BFX4 U13087 ( .A(n12286), .Z(n12287) );
  HS65_LH_BFX4 U13088 ( .A(n12287), .Z(n12288) );
  HS65_LH_BFX4 U13089 ( .A(n12288), .Z(n12289) );
  HS65_LH_BFX4 U13090 ( .A(n12289), .Z(n12290) );
  HS65_LH_BFX4 U13091 ( .A(n12292), .Z(n12291) );
  HS65_LH_BFX4 U13092 ( .A(n12293), .Z(n12292) );
  HS65_LH_BFX4 U13093 ( .A(n12294), .Z(n12293) );
  HS65_LH_BFX4 U13094 ( .A(n12295), .Z(n12294) );
  HS65_LH_BFX4 U13095 ( .A(n12296), .Z(n12295) );
  HS65_LH_BFX4 U13096 ( .A(n12297), .Z(n12296) );
  HS65_LH_BFX4 U13097 ( .A(n12298), .Z(n12297) );
  HS65_LH_BFX4 U13098 ( .A(n12299), .Z(n12298) );
  HS65_LH_BFX4 U13099 ( .A(n12300), .Z(n12299) );
  HS65_LH_BFX4 U13100 ( .A(n12301), .Z(n12300) );
  HS65_LH_BFX4 U13101 ( .A(n14052), .Z(n12301) );
  HS65_LH_BFX4 U13102 ( .A(n12324), .Z(n12302) );
  HS65_LH_BFX4 U13103 ( .A(\u_DataPath/jaddr_i [18]), .Z(n12303) );
  HS65_LH_BFX4 U13104 ( .A(n12303), .Z(n12304) );
  HS65_LH_BFX4 U13105 ( .A(n12304), .Z(n12305) );
  HS65_LH_BFX4 U13106 ( .A(n12305), .Z(n12306) );
  HS65_LH_BFX4 U13107 ( .A(n12306), .Z(n12307) );
  HS65_LH_BFX4 U13108 ( .A(n12307), .Z(n12308) );
  HS65_LH_BFX4 U13109 ( .A(n12308), .Z(n12309) );
  HS65_LH_BFX4 U13110 ( .A(n12309), .Z(n12310) );
  HS65_LH_BFX4 U13111 ( .A(n12310), .Z(n12311) );
  HS65_LH_BFX4 U13112 ( .A(n12311), .Z(n12312) );
  HS65_LH_BFX4 U13113 ( .A(n12312), .Z(n12313) );
  HS65_LH_BFX4 U13114 ( .A(n12313), .Z(n12314) );
  HS65_LH_BFX4 U13115 ( .A(n12314), .Z(n12315) );
  HS65_LH_BFX4 U13116 ( .A(n12315), .Z(n12316) );
  HS65_LH_BFX4 U13117 ( .A(n12316), .Z(n12317) );
  HS65_LH_BFX4 U13118 ( .A(n12317), .Z(n12318) );
  HS65_LH_BFX4 U13119 ( .A(n12318), .Z(n12319) );
  HS65_LH_BFX4 U13120 ( .A(n12319), .Z(n12320) );
  HS65_LH_BFX4 U13121 ( .A(n12320), .Z(n12321) );
  HS65_LH_BFX4 U13122 ( .A(n12321), .Z(n12322) );
  HS65_LH_CNIVX3 U13123 ( .A(n12322), .Z(n12323) );
  HS65_LH_CNIVX3 U13124 ( .A(n12323), .Z(n12324) );
  HS65_LH_BFX4 U13125 ( .A(n12327), .Z(n12325) );
  HS65_LH_BFX4 U13126 ( .A(n12338), .Z(n12326) );
  HS65_LH_BFX4 U13127 ( .A(n12326), .Z(n12327) );
  HS65_LH_BFX4 U13128 ( .A(n12336), .Z(n12328) );
  HS65_LH_BFX4 U13129 ( .A(n12328), .Z(n12329) );
  HS65_LH_BFX4 U13130 ( .A(n12329), .Z(n12330) );
  HS65_LH_BFX4 U13131 ( .A(n12330), .Z(n12331) );
  HS65_LH_BFX4 U13132 ( .A(n12331), .Z(n12332) );
  HS65_LH_BFX4 U13133 ( .A(n12332), .Z(n12333) );
  HS65_LH_BFX4 U13134 ( .A(n12333), .Z(n12334) );
  HS65_LH_BFX4 U13135 ( .A(n12334), .Z(n12335) );
  HS65_LH_BFX4 U13136 ( .A(n12337), .Z(n12336) );
  HS65_LH_BFX4 U13137 ( .A(n12340), .Z(n12337) );
  HS65_LH_BFX4 U13138 ( .A(n12339), .Z(n12338) );
  HS65_LH_BFX4 U13139 ( .A(n12335), .Z(n12339) );
  HS65_LH_BFX4 U13140 ( .A(n12341), .Z(n12340) );
  HS65_LH_BFX4 U13141 ( .A(n12342), .Z(n12341) );
  HS65_LH_BFX4 U13142 ( .A(n12343), .Z(n12342) );
  HS65_LH_BFX4 U13143 ( .A(n12344), .Z(n12343) );
  HS65_LH_BFX4 U13144 ( .A(n12345), .Z(n12344) );
  HS65_LH_BFX4 U13145 ( .A(n12346), .Z(n12345) );
  HS65_LH_BFX4 U13146 ( .A(n14054), .Z(n12346) );
  HS65_LH_BFX4 U13147 ( .A(n12370), .Z(n12347) );
  HS65_LH_BFX4 U13148 ( .A(\u_DataPath/jaddr_i [20]), .Z(n12348) );
  HS65_LH_BFX4 U13149 ( .A(n12348), .Z(n12349) );
  HS65_LH_BFX4 U13150 ( .A(n12349), .Z(n12350) );
  HS65_LH_BFX4 U13151 ( .A(n12350), .Z(n12351) );
  HS65_LH_BFX4 U13152 ( .A(n12351), .Z(n12352) );
  HS65_LH_BFX4 U13153 ( .A(n12352), .Z(n12353) );
  HS65_LH_BFX4 U13154 ( .A(n12353), .Z(n12354) );
  HS65_LH_BFX4 U13155 ( .A(n12354), .Z(n12355) );
  HS65_LH_BFX4 U13156 ( .A(n12355), .Z(n12356) );
  HS65_LH_BFX4 U13157 ( .A(n12356), .Z(n12357) );
  HS65_LH_BFX4 U13158 ( .A(n12357), .Z(n12358) );
  HS65_LH_BFX4 U13159 ( .A(n12358), .Z(n12359) );
  HS65_LH_BFX4 U13160 ( .A(n12359), .Z(n12360) );
  HS65_LH_BFX4 U13161 ( .A(n12360), .Z(n12361) );
  HS65_LH_BFX4 U13162 ( .A(n12361), .Z(n12362) );
  HS65_LH_BFX4 U13163 ( .A(n12362), .Z(n12363) );
  HS65_LH_BFX4 U13164 ( .A(n12363), .Z(n12364) );
  HS65_LH_BFX4 U13165 ( .A(n12364), .Z(n12365) );
  HS65_LH_BFX4 U13166 ( .A(n12365), .Z(n12366) );
  HS65_LH_BFX4 U13167 ( .A(n12366), .Z(n12367) );
  HS65_LH_BFX4 U13168 ( .A(n12367), .Z(n12368) );
  HS65_LH_CNIVX3 U13169 ( .A(n12368), .Z(n12369) );
  HS65_LH_CNIVX3 U13170 ( .A(n12369), .Z(n12370) );
  HS65_LH_BFX4 U13171 ( .A(\u_DataPath/jaddr_i [21]), .Z(n12371) );
  HS65_LH_BFX4 U13172 ( .A(n12371), .Z(n12372) );
  HS65_LH_BFX4 U13173 ( .A(n12372), .Z(n12373) );
  HS65_LH_BFX4 U13174 ( .A(n12373), .Z(n12374) );
  HS65_LH_BFX4 U13175 ( .A(n12374), .Z(n12375) );
  HS65_LH_BFX4 U13176 ( .A(n12375), .Z(n12376) );
  HS65_LH_BFX4 U13177 ( .A(n12376), .Z(n12377) );
  HS65_LH_BFX4 U13178 ( .A(n12377), .Z(n12378) );
  HS65_LH_BFX4 U13179 ( .A(n12378), .Z(n12379) );
  HS65_LH_BFX4 U13180 ( .A(n12379), .Z(n12380) );
  HS65_LH_BFX4 U13181 ( .A(n12380), .Z(n12381) );
  HS65_LH_BFX4 U13182 ( .A(n12383), .Z(n12382) );
  HS65_LH_BFX4 U13183 ( .A(n12384), .Z(n12383) );
  HS65_LH_BFX4 U13184 ( .A(n12385), .Z(n12384) );
  HS65_LH_BFX4 U13185 ( .A(n12386), .Z(n12385) );
  HS65_LH_BFX4 U13186 ( .A(n12387), .Z(n12386) );
  HS65_LH_BFX4 U13187 ( .A(n12388), .Z(n12387) );
  HS65_LH_BFX4 U13188 ( .A(n12389), .Z(n12388) );
  HS65_LH_BFX4 U13189 ( .A(n12390), .Z(n12389) );
  HS65_LH_BFX4 U13190 ( .A(n12391), .Z(n12390) );
  HS65_LH_BFX4 U13191 ( .A(n12392), .Z(n12391) );
  HS65_LH_BFX4 U13192 ( .A(n14055), .Z(n12392) );
  HS65_LH_BFX4 U13193 ( .A(n12395), .Z(n12393) );
  HS65_LH_BFX4 U13194 ( .A(n13578), .Z(n12394) );
  HS65_LH_BFX4 U13195 ( .A(n12394), .Z(n12395) );
  HS65_LH_BFX4 U13196 ( .A(\u_DataPath/jaddr_i [22]), .Z(n12396) );
  HS65_LH_BFX4 U13197 ( .A(n12396), .Z(n12397) );
  HS65_LH_BFX4 U13198 ( .A(n12397), .Z(n12398) );
  HS65_LH_BFX4 U13199 ( .A(n12398), .Z(n12399) );
  HS65_LH_BFX4 U13200 ( .A(n12399), .Z(n12400) );
  HS65_LH_BFX4 U13201 ( .A(n12400), .Z(n12401) );
  HS65_LH_BFX4 U13202 ( .A(n12401), .Z(n12402) );
  HS65_LH_BFX4 U13203 ( .A(n12402), .Z(n12403) );
  HS65_LH_BFX4 U13204 ( .A(n12403), .Z(n12404) );
  HS65_LH_BFX4 U13205 ( .A(n12404), .Z(n12405) );
  HS65_LH_BFX4 U13206 ( .A(n12405), .Z(n12406) );
  HS65_LH_BFX4 U13207 ( .A(n12406), .Z(n12407) );
  HS65_LH_BFX4 U13208 ( .A(n12407), .Z(n12408) );
  HS65_LH_BFX4 U13209 ( .A(n12408), .Z(n12409) );
  HS65_LH_BFX4 U13210 ( .A(n12409), .Z(n12410) );
  HS65_LH_BFX4 U13211 ( .A(n12410), .Z(n12411) );
  HS65_LH_BFX4 U13212 ( .A(n12411), .Z(n12412) );
  HS65_LH_BFX4 U13213 ( .A(n12412), .Z(n12413) );
  HS65_LH_BFX4 U13214 ( .A(n12416), .Z(n12414) );
  HS65_LH_BFX4 U13215 ( .A(n12426), .Z(n12415) );
  HS65_LH_BFX4 U13216 ( .A(n12415), .Z(n12416) );
  HS65_LH_BFX4 U13217 ( .A(\u_DataPath/jaddr_i [23]), .Z(n12417) );
  HS65_LH_BFX4 U13218 ( .A(n12417), .Z(n12418) );
  HS65_LH_BFX4 U13219 ( .A(n12418), .Z(n12419) );
  HS65_LH_BFX4 U13220 ( .A(n12419), .Z(n12420) );
  HS65_LH_BFX4 U13221 ( .A(n12420), .Z(n12421) );
  HS65_LH_BFX4 U13222 ( .A(n12421), .Z(n12422) );
  HS65_LH_BFX4 U13223 ( .A(n12422), .Z(n12423) );
  HS65_LH_BFX4 U13224 ( .A(n12423), .Z(n12424) );
  HS65_LH_BFX4 U13225 ( .A(n12424), .Z(n12425) );
  HS65_LH_BFX4 U13226 ( .A(n12427), .Z(n12426) );
  HS65_LH_BFX4 U13227 ( .A(n12428), .Z(n12427) );
  HS65_LH_BFX4 U13228 ( .A(n12429), .Z(n12428) );
  HS65_LH_BFX4 U13229 ( .A(n12430), .Z(n12429) );
  HS65_LH_BFX4 U13230 ( .A(n12431), .Z(n12430) );
  HS65_LH_BFX4 U13231 ( .A(n12432), .Z(n12431) );
  HS65_LH_BFX4 U13232 ( .A(n12433), .Z(n12432) );
  HS65_LH_BFX4 U13233 ( .A(n12434), .Z(n12433) );
  HS65_LH_BFX4 U13234 ( .A(n12435), .Z(n12434) );
  HS65_LH_BFX4 U13235 ( .A(n14056), .Z(n12435) );
  HS65_LH_BFX4 U13236 ( .A(n12438), .Z(n12436) );
  HS65_LH_BFX4 U13237 ( .A(n12446), .Z(n12437) );
  HS65_LH_BFX4 U13238 ( .A(n12437), .Z(n12438) );
  HS65_LH_BFX4 U13239 ( .A(\u_DataPath/jaddr_i [24]), .Z(n12439) );
  HS65_LH_BFX4 U13240 ( .A(n12439), .Z(n12440) );
  HS65_LH_BFX4 U13241 ( .A(n12440), .Z(n12441) );
  HS65_LH_BFX4 U13242 ( .A(n12441), .Z(n12442) );
  HS65_LH_BFX4 U13243 ( .A(n12442), .Z(n12443) );
  HS65_LH_BFX4 U13244 ( .A(n12443), .Z(n12444) );
  HS65_LH_BFX4 U13245 ( .A(n12444), .Z(n12445) );
  HS65_LH_BFX4 U13246 ( .A(n12447), .Z(n12446) );
  HS65_LH_BFX4 U13247 ( .A(n12448), .Z(n12447) );
  HS65_LH_BFX4 U13248 ( .A(n12449), .Z(n12448) );
  HS65_LH_BFX4 U13249 ( .A(n12450), .Z(n12449) );
  HS65_LH_BFX4 U13250 ( .A(n12451), .Z(n12450) );
  HS65_LH_BFX4 U13251 ( .A(n12453), .Z(n12451) );
  HS65_LH_BFX4 U13252 ( .A(n12445), .Z(n12452) );
  HS65_LH_BFX4 U13253 ( .A(n12454), .Z(n12453) );
  HS65_LH_BFX4 U13254 ( .A(n12455), .Z(n12454) );
  HS65_LH_BFX4 U13255 ( .A(n12456), .Z(n12455) );
  HS65_LH_BFX4 U13256 ( .A(n12457), .Z(n12456) );
  HS65_LH_BFX4 U13257 ( .A(n14057), .Z(n12457) );
  HS65_LH_BFX4 U13258 ( .A(n12471), .Z(n12458) );
  HS65_LH_BFX4 U13259 ( .A(\u_DataPath/jaddr_i [25]), .Z(n12459) );
  HS65_LH_BFX4 U13260 ( .A(n12459), .Z(n12460) );
  HS65_LH_BFX4 U13261 ( .A(n12460), .Z(n12461) );
  HS65_LH_BFX4 U13262 ( .A(n12461), .Z(n12462) );
  HS65_LH_BFX4 U13263 ( .A(n12462), .Z(n12463) );
  HS65_LH_BFX4 U13264 ( .A(n12463), .Z(n12464) );
  HS65_LH_BFX4 U13265 ( .A(n12464), .Z(n12465) );
  HS65_LH_BFX4 U13266 ( .A(n12465), .Z(n12466) );
  HS65_LH_BFX4 U13267 ( .A(n12466), .Z(n12467) );
  HS65_LH_BFX4 U13268 ( .A(n12467), .Z(n12468) );
  HS65_LH_BFX4 U13269 ( .A(n12468), .Z(n12469) );
  HS65_LH_BFX4 U13270 ( .A(n12469), .Z(n12470) );
  HS65_LH_BFX4 U13271 ( .A(n12472), .Z(n12471) );
  HS65_LH_BFX4 U13272 ( .A(n12473), .Z(n12472) );
  HS65_LH_BFX4 U13273 ( .A(n12474), .Z(n12473) );
  HS65_LH_BFX4 U13274 ( .A(n12475), .Z(n12474) );
  HS65_LH_BFX4 U13275 ( .A(n12476), .Z(n12475) );
  HS65_LH_BFX4 U13276 ( .A(n12477), .Z(n12476) );
  HS65_LH_BFX4 U13277 ( .A(n12478), .Z(n12477) );
  HS65_LH_BFX4 U13278 ( .A(n14058), .Z(n12478) );
  HS65_LH_BFX4 U13279 ( .A(n12470), .Z(n12479) );
  HS65_LH_BFX4 U13280 ( .A(n12482), .Z(n12480) );
  HS65_LH_BFX4 U13281 ( .A(n13654), .Z(n12481) );
  HS65_LH_BFX4 U13282 ( .A(n12481), .Z(n12482) );
  HS65_LH_BFX4 U13283 ( .A(opcode_i[3]), .Z(n12483) );
  HS65_LH_BFX4 U13284 ( .A(n10371), .Z(n12484) );
  HS65_LH_BFX2 U13285 ( .A(n12493), .Z(n12485) );
  HS65_LH_BFX4 U13286 ( .A(n12484), .Z(n12486) );
  HS65_LH_BFX4 U13288 ( .A(n12486), .Z(n12488) );
  HS65_LH_BFX2 U13289 ( .A(n15707), .Z(n12489) );
  HS65_LH_BFX4 U13290 ( .A(n12492), .Z(n12490) );
  HS65_LH_BFX2 U13291 ( .A(n12489), .Z(n12491) );
  HS65_LH_BFX4 U13292 ( .A(n12494), .Z(n12492) );
  HS65_LH_BFX2 U13293 ( .A(n12498), .Z(n12493) );
  HS65_LH_BFX4 U13294 ( .A(n13640), .Z(n12494) );
  HS65_LH_BFX2 U13295 ( .A(n12491), .Z(n12495) );
  HS65_LH_BFX2 U13296 ( .A(n12495), .Z(n12496) );
  HS65_LH_BFX2 U13297 ( .A(n12496), .Z(n12497) );
  HS65_LH_BFX2 U13298 ( .A(n12499), .Z(n12498) );
  HS65_LH_BFX2 U13299 ( .A(n12500), .Z(n12499) );
  HS65_LH_BFX2 U13300 ( .A(n12501), .Z(n12500) );
  HS65_LH_BFX2 U13301 ( .A(n12502), .Z(n12501) );
  HS65_LH_BFX2 U13302 ( .A(n12503), .Z(n12502) );
  HS65_LH_BFX2 U13303 ( .A(n12497), .Z(n12503) );
  HS65_LH_BFX4 U13304 ( .A(n12506), .Z(n12504) );
  HS65_LH_BFX4 U13305 ( .A(n12507), .Z(n12505) );
  HS65_LH_BFX4 U13306 ( .A(n12508), .Z(n12506) );
  HS65_LH_BFX4 U13307 ( .A(n12509), .Z(n12507) );
  HS65_LH_BFX4 U13308 ( .A(n12510), .Z(n12508) );
  HS65_LH_BFX4 U13309 ( .A(n12511), .Z(n12509) );
  HS65_LH_BFX4 U13310 ( .A(n12512), .Z(n12510) );
  HS65_LH_BFX4 U13311 ( .A(n12513), .Z(n12511) );
  HS65_LH_BFX4 U13312 ( .A(n12514), .Z(n12512) );
  HS65_LH_BFX4 U13313 ( .A(n12515), .Z(n12513) );
  HS65_LH_BFX4 U13314 ( .A(n12516), .Z(n12514) );
  HS65_LH_BFX4 U13315 ( .A(n12517), .Z(n12515) );
  HS65_LH_BFX4 U13316 ( .A(n12518), .Z(n12516) );
  HS65_LH_BFX4 U13317 ( .A(n12519), .Z(n12517) );
  HS65_LH_BFX4 U13318 ( .A(n12520), .Z(n12518) );
  HS65_LH_BFX4 U13319 ( .A(n12521), .Z(n12519) );
  HS65_LH_BFX4 U13320 ( .A(n12522), .Z(n12520) );
  HS65_LH_BFX4 U13321 ( .A(n12523), .Z(n12521) );
  HS65_LH_BFX4 U13322 ( .A(n12524), .Z(n12522) );
  HS65_LH_BFX4 U13323 ( .A(n12525), .Z(n12523) );
  HS65_LH_BFX4 U13324 ( .A(n12526), .Z(n12524) );
  HS65_LH_BFX4 U13325 ( .A(n12527), .Z(n12525) );
  HS65_LH_BFX4 U13326 ( .A(n12528), .Z(n12526) );
  HS65_LH_BFX4 U13327 ( .A(n12529), .Z(n12527) );
  HS65_LH_BFX4 U13328 ( .A(n12530), .Z(n12528) );
  HS65_LH_BFX4 U13329 ( .A(n12531), .Z(n12529) );
  HS65_LH_BFX4 U13330 ( .A(n12532), .Z(n12530) );
  HS65_LH_BFX4 U13331 ( .A(n12533), .Z(n12531) );
  HS65_LH_BFX4 U13332 ( .A(n12534), .Z(n12532) );
  HS65_LH_BFX4 U13333 ( .A(n12535), .Z(n12533) );
  HS65_LH_BFX4 U13334 ( .A(n12536), .Z(n12534) );
  HS65_LH_BFX4 U13335 ( .A(n12537), .Z(n12535) );
  HS65_LH_BFX4 U13336 ( .A(n12538), .Z(n12536) );
  HS65_LH_BFX4 U13337 ( .A(n12539), .Z(n12537) );
  HS65_LH_BFX4 U13338 ( .A(n12540), .Z(n12538) );
  HS65_LH_BFX4 U13339 ( .A(n12541), .Z(n12539) );
  HS65_LH_BFX4 U13340 ( .A(n12542), .Z(n12540) );
  HS65_LH_BFX4 U13341 ( .A(n12543), .Z(n12541) );
  HS65_LH_BFX4 U13342 ( .A(n12544), .Z(n12542) );
  HS65_LH_BFX4 U13343 ( .A(n12545), .Z(n12543) );
  HS65_LH_BFX4 U13344 ( .A(n12546), .Z(n12544) );
  HS65_LH_BFX4 U13345 ( .A(n12547), .Z(n12545) );
  HS65_LH_BFX4 U13346 ( .A(n12548), .Z(n12546) );
  HS65_LH_BFX4 U13347 ( .A(n12549), .Z(n12547) );
  HS65_LH_BFX4 U13348 ( .A(\u_DataPath/pc_4_i [0]), .Z(n12548) );
  HS65_LH_BFX4 U13349 ( .A(n12550), .Z(n12549) );
  HS65_LH_BFX4 U13350 ( .A(\u_DataPath/pc4_to_idexreg_i [0]), .Z(n12550) );
  HS65_LH_BFX4 U13351 ( .A(n12553), .Z(n12551) );
  HS65_LH_BFX4 U13352 ( .A(n12554), .Z(n12552) );
  HS65_LH_BFX4 U13353 ( .A(n12555), .Z(n12553) );
  HS65_LH_BFX4 U13354 ( .A(n12556), .Z(n12554) );
  HS65_LH_BFX4 U13355 ( .A(n12557), .Z(n12555) );
  HS65_LH_BFX4 U13356 ( .A(n12558), .Z(n12556) );
  HS65_LH_BFX4 U13357 ( .A(n12559), .Z(n12557) );
  HS65_LH_BFX4 U13358 ( .A(n12560), .Z(n12558) );
  HS65_LH_BFX4 U13359 ( .A(n12561), .Z(n12559) );
  HS65_LH_BFX4 U13360 ( .A(n12562), .Z(n12560) );
  HS65_LH_BFX4 U13361 ( .A(n12563), .Z(n12561) );
  HS65_LH_BFX4 U13362 ( .A(n12564), .Z(n12562) );
  HS65_LH_BFX4 U13363 ( .A(n12565), .Z(n12563) );
  HS65_LH_BFX4 U13364 ( .A(n12566), .Z(n12564) );
  HS65_LH_BFX4 U13365 ( .A(n12567), .Z(n12565) );
  HS65_LH_BFX4 U13366 ( .A(n12568), .Z(n12566) );
  HS65_LH_BFX4 U13367 ( .A(n12569), .Z(n12567) );
  HS65_LH_BFX4 U13368 ( .A(n12570), .Z(n12568) );
  HS65_LH_BFX4 U13369 ( .A(n12571), .Z(n12569) );
  HS65_LH_BFX4 U13370 ( .A(n12572), .Z(n12570) );
  HS65_LH_BFX4 U13371 ( .A(n12573), .Z(n12571) );
  HS65_LH_BFX4 U13372 ( .A(n12574), .Z(n12572) );
  HS65_LH_BFX4 U13373 ( .A(n12575), .Z(n12573) );
  HS65_LH_BFX4 U13374 ( .A(n12576), .Z(n12574) );
  HS65_LH_BFX4 U13375 ( .A(n12577), .Z(n12575) );
  HS65_LH_BFX4 U13376 ( .A(n12578), .Z(n12576) );
  HS65_LH_BFX4 U13377 ( .A(n12579), .Z(n12577) );
  HS65_LH_BFX4 U13378 ( .A(n12580), .Z(n12578) );
  HS65_LH_BFX4 U13379 ( .A(n12581), .Z(n12579) );
  HS65_LH_BFX4 U13380 ( .A(n12582), .Z(n12580) );
  HS65_LH_BFX4 U13381 ( .A(n12583), .Z(n12581) );
  HS65_LH_BFX4 U13382 ( .A(n12584), .Z(n12582) );
  HS65_LH_BFX4 U13383 ( .A(n12585), .Z(n12583) );
  HS65_LH_BFX4 U13384 ( .A(n12586), .Z(n12584) );
  HS65_LH_BFX4 U13385 ( .A(n12587), .Z(n12585) );
  HS65_LH_BFX4 U13386 ( .A(n12588), .Z(n12586) );
  HS65_LH_BFX4 U13387 ( .A(n12589), .Z(n12587) );
  HS65_LH_BFX4 U13388 ( .A(n12590), .Z(n12588) );
  HS65_LH_BFX4 U13389 ( .A(n12591), .Z(n12589) );
  HS65_LH_BFX4 U13390 ( .A(n12592), .Z(n12590) );
  HS65_LH_BFX4 U13391 ( .A(n12593), .Z(n12591) );
  HS65_LH_BFX4 U13392 ( .A(n12594), .Z(n12592) );
  HS65_LH_BFX4 U13393 ( .A(n12595), .Z(n12593) );
  HS65_LH_BFX4 U13394 ( .A(n12596), .Z(n12594) );
  HS65_LH_BFX4 U13395 ( .A(\u_DataPath/pc_4_i [1]), .Z(n12595) );
  HS65_LH_BFX4 U13396 ( .A(n12597), .Z(n12596) );
  HS65_LH_BFX4 U13397 ( .A(\u_DataPath/pc4_to_idexreg_i [1]), .Z(n12597) );
  HS65_LH_BFX4 U13398 ( .A(n12600), .Z(n12598) );
  HS65_LH_BFX4 U13399 ( .A(n12601), .Z(n12599) );
  HS65_LH_BFX4 U13400 ( .A(n12602), .Z(n12600) );
  HS65_LH_BFX4 U13401 ( .A(n12603), .Z(n12601) );
  HS65_LH_BFX4 U13402 ( .A(n12604), .Z(n12602) );
  HS65_LH_BFX4 U13403 ( .A(n12605), .Z(n12603) );
  HS65_LH_BFX4 U13404 ( .A(n12606), .Z(n12604) );
  HS65_LH_BFX4 U13405 ( .A(n12607), .Z(n12605) );
  HS65_LH_BFX4 U13406 ( .A(n12608), .Z(n12606) );
  HS65_LH_BFX4 U13407 ( .A(n12609), .Z(n12607) );
  HS65_LH_BFX4 U13408 ( .A(n12610), .Z(n12608) );
  HS65_LH_BFX4 U13409 ( .A(n12611), .Z(n12609) );
  HS65_LH_BFX4 U13410 ( .A(n12612), .Z(n12610) );
  HS65_LH_BFX4 U13411 ( .A(n12613), .Z(n12611) );
  HS65_LH_BFX4 U13412 ( .A(n12614), .Z(n12612) );
  HS65_LH_BFX4 U13413 ( .A(n12615), .Z(n12613) );
  HS65_LH_BFX4 U13414 ( .A(n12617), .Z(n12614) );
  HS65_LH_BFX4 U13415 ( .A(n12616), .Z(n12615) );
  HS65_LH_BFX4 U13416 ( .A(n12618), .Z(n12616) );
  HS65_LH_BFX4 U13417 ( .A(n12619), .Z(n12617) );
  HS65_LH_BFX4 U13418 ( .A(n12620), .Z(n12618) );
  HS65_LH_BFX4 U13419 ( .A(n12621), .Z(n12619) );
  HS65_LH_BFX4 U13420 ( .A(n12622), .Z(n12620) );
  HS65_LH_BFX4 U13421 ( .A(n12623), .Z(n12621) );
  HS65_LH_BFX4 U13422 ( .A(n12624), .Z(n12622) );
  HS65_LH_BFX4 U13423 ( .A(n12625), .Z(n12623) );
  HS65_LH_BFX4 U13424 ( .A(n12626), .Z(n12624) );
  HS65_LH_BFX4 U13425 ( .A(n12627), .Z(n12625) );
  HS65_LH_BFX4 U13426 ( .A(n12628), .Z(n12626) );
  HS65_LH_BFX4 U13427 ( .A(n12629), .Z(n12627) );
  HS65_LH_BFX4 U13428 ( .A(n12630), .Z(n12628) );
  HS65_LH_BFX4 U13429 ( .A(n12631), .Z(n12629) );
  HS65_LH_BFX4 U13430 ( .A(n12632), .Z(n12630) );
  HS65_LH_BFX4 U13431 ( .A(n12633), .Z(n12631) );
  HS65_LH_BFX4 U13432 ( .A(n12634), .Z(n12632) );
  HS65_LH_BFX4 U13433 ( .A(n12635), .Z(n12633) );
  HS65_LH_BFX4 U13434 ( .A(n12636), .Z(n12634) );
  HS65_LH_BFX4 U13435 ( .A(n12640), .Z(n12635) );
  HS65_LH_BFX4 U13436 ( .A(n12638), .Z(n12636) );
  HS65_LH_BFX4 U13437 ( .A(addr_to_iram_0), .Z(n12637) );
  HS65_LH_BFX4 U13438 ( .A(n12641), .Z(n12638) );
  HS65_LH_CNIVX3 U13439 ( .A(n14106), .Z(n12639) );
  HS65_LH_CNIVX3 U13440 ( .A(n12639), .Z(n12640) );
  HS65_LL_IVX2 U13441 ( .A(n17244), .Z(n14005) );
  HS65_LH_BFX4 U13442 ( .A(n12642), .Z(n12641) );
  HS65_LH_BFX4 U13443 ( .A(n12643), .Z(n12642) );
  HS65_LH_BFX4 U13444 ( .A(\u_DataPath/pc4_to_idexreg_i [2]), .Z(n12643) );
  HS65_LH_BFX4 U13445 ( .A(n12646), .Z(n12644) );
  HS65_LH_BFX4 U13446 ( .A(n12647), .Z(n12645) );
  HS65_LH_BFX4 U13447 ( .A(n12648), .Z(n12646) );
  HS65_LH_BFX4 U13448 ( .A(n12649), .Z(n12647) );
  HS65_LH_BFX4 U13449 ( .A(n12650), .Z(n12648) );
  HS65_LH_BFX4 U13450 ( .A(n12651), .Z(n12649) );
  HS65_LH_BFX4 U13451 ( .A(n12652), .Z(n12650) );
  HS65_LH_BFX4 U13452 ( .A(n12653), .Z(n12651) );
  HS65_LH_BFX4 U13453 ( .A(n12654), .Z(n12652) );
  HS65_LH_BFX4 U13454 ( .A(n12655), .Z(n12653) );
  HS65_LH_BFX4 U13455 ( .A(n12656), .Z(n12654) );
  HS65_LH_BFX4 U13456 ( .A(n12657), .Z(n12655) );
  HS65_LH_BFX4 U13457 ( .A(n12658), .Z(n12656) );
  HS65_LH_BFX4 U13458 ( .A(n12659), .Z(n12657) );
  HS65_LH_BFX4 U13459 ( .A(n12660), .Z(n12658) );
  HS65_LH_BFX4 U13460 ( .A(n12661), .Z(n12659) );
  HS65_LH_BFX4 U13461 ( .A(n12662), .Z(n12660) );
  HS65_LH_BFX4 U13462 ( .A(n12663), .Z(n12661) );
  HS65_LH_BFX4 U13463 ( .A(n12664), .Z(n12662) );
  HS65_LH_BFX4 U13464 ( .A(n12665), .Z(n12663) );
  HS65_LH_BFX4 U13465 ( .A(n12666), .Z(n12664) );
  HS65_LH_BFX4 U13466 ( .A(n12667), .Z(n12665) );
  HS65_LH_BFX4 U13467 ( .A(n12668), .Z(n12666) );
  HS65_LH_BFX4 U13468 ( .A(n12669), .Z(n12667) );
  HS65_LH_BFX4 U13469 ( .A(n12670), .Z(n12668) );
  HS65_LH_BFX4 U13470 ( .A(n14107), .Z(n12669) );
  HS65_LH_BFX4 U13471 ( .A(n12671), .Z(n12670) );
  HS65_LH_BFX4 U13472 ( .A(\u_DataPath/pc4_to_idexreg_i [3]), .Z(n12671) );
  HS65_LH_BFX4 U13473 ( .A(n12674), .Z(n12672) );
  HS65_LH_BFX4 U13474 ( .A(n12675), .Z(n12673) );
  HS65_LH_BFX4 U13475 ( .A(n12676), .Z(n12674) );
  HS65_LH_BFX4 U13476 ( .A(n12677), .Z(n12675) );
  HS65_LH_BFX4 U13477 ( .A(n12678), .Z(n12676) );
  HS65_LH_BFX4 U13478 ( .A(n12679), .Z(n12677) );
  HS65_LH_BFX4 U13479 ( .A(n12680), .Z(n12678) );
  HS65_LH_BFX4 U13480 ( .A(n12681), .Z(n12679) );
  HS65_LH_BFX4 U13481 ( .A(n12682), .Z(n12680) );
  HS65_LH_BFX4 U13482 ( .A(n12683), .Z(n12681) );
  HS65_LH_BFX4 U13483 ( .A(n12684), .Z(n12682) );
  HS65_LH_BFX4 U13484 ( .A(n12685), .Z(n12683) );
  HS65_LH_BFX4 U13485 ( .A(n12686), .Z(n12684) );
  HS65_LH_BFX4 U13486 ( .A(n12687), .Z(n12685) );
  HS65_LH_BFX4 U13487 ( .A(n12688), .Z(n12686) );
  HS65_LH_BFX4 U13488 ( .A(n12689), .Z(n12687) );
  HS65_LH_BFX4 U13489 ( .A(n12690), .Z(n12688) );
  HS65_LH_BFX4 U13490 ( .A(n12691), .Z(n12689) );
  HS65_LH_BFX4 U13491 ( .A(n12692), .Z(n12690) );
  HS65_LH_BFX4 U13492 ( .A(n12693), .Z(n12691) );
  HS65_LH_BFX4 U13493 ( .A(n12694), .Z(n12692) );
  HS65_LH_BFX4 U13494 ( .A(n12695), .Z(n12693) );
  HS65_LH_BFX4 U13495 ( .A(n12696), .Z(n12694) );
  HS65_LH_BFX4 U13496 ( .A(n12697), .Z(n12695) );
  HS65_LH_BFX4 U13497 ( .A(n12698), .Z(n12696) );
  HS65_LH_BFX4 U13498 ( .A(n12699), .Z(n12697) );
  HS65_LH_BFX4 U13499 ( .A(n12700), .Z(n12698) );
  HS65_LH_BFX4 U13500 ( .A(n12701), .Z(n12699) );
  HS65_LH_BFX4 U13501 ( .A(n12702), .Z(n12700) );
  HS65_LH_BFX4 U13502 ( .A(n12703), .Z(n12701) );
  HS65_LH_BFX4 U13503 ( .A(n12704), .Z(n12702) );
  HS65_LH_BFX4 U13504 ( .A(n12705), .Z(n12703) );
  HS65_LH_BFX4 U13505 ( .A(n12707), .Z(n12704) );
  HS65_LH_BFX4 U13506 ( .A(n12706), .Z(n12705) );
  HS65_LH_BFX4 U13507 ( .A(n12708), .Z(n12706) );
  HS65_LH_BFX4 U13508 ( .A(n12709), .Z(n12707) );
  HS65_LH_BFX4 U13509 ( .A(n12710), .Z(n12708) );
  HS65_LH_BFX4 U13510 ( .A(n12711), .Z(n12709) );
  HS65_LH_BFX4 U13511 ( .A(n12712), .Z(n12710) );
  HS65_LH_BFX4 U13512 ( .A(n12713), .Z(n12711) );
  HS65_LH_BFX4 U13513 ( .A(n12714), .Z(n12712) );
  HS65_LH_BFX4 U13514 ( .A(n14081), .Z(n12713) );
  HS65_LH_BFX4 U13515 ( .A(n12715), .Z(n12714) );
  HS65_LH_BFX4 U13516 ( .A(n12716), .Z(n12715) );
  HS65_LH_BFX4 U13517 ( .A(\u_DataPath/pc4_to_idexreg_i [4]), .Z(n12716) );
  HS65_LH_BFX4 U13518 ( .A(n17241), .Z(n12717) );
  HS65_LH_BFX4 U13519 ( .A(n12720), .Z(n12718) );
  HS65_LH_BFX4 U13520 ( .A(n12721), .Z(n12719) );
  HS65_LH_BFX4 U13521 ( .A(n12722), .Z(n12720) );
  HS65_LH_BFX4 U13522 ( .A(n12723), .Z(n12721) );
  HS65_LH_BFX4 U13523 ( .A(n12724), .Z(n12722) );
  HS65_LH_BFX4 U13524 ( .A(n12725), .Z(n12723) );
  HS65_LH_BFX4 U13525 ( .A(n12726), .Z(n12724) );
  HS65_LH_BFX4 U13526 ( .A(n12727), .Z(n12725) );
  HS65_LH_BFX4 U13527 ( .A(n12728), .Z(n12726) );
  HS65_LH_BFX4 U13528 ( .A(n12729), .Z(n12727) );
  HS65_LH_BFX4 U13529 ( .A(n12730), .Z(n12728) );
  HS65_LH_BFX4 U13530 ( .A(n12731), .Z(n12729) );
  HS65_LH_BFX4 U13531 ( .A(n12732), .Z(n12730) );
  HS65_LH_BFX4 U13532 ( .A(n12733), .Z(n12731) );
  HS65_LH_BFX4 U13533 ( .A(n12734), .Z(n12732) );
  HS65_LH_BFX4 U13534 ( .A(n12735), .Z(n12733) );
  HS65_LH_BFX4 U13535 ( .A(n12736), .Z(n12734) );
  HS65_LH_BFX4 U13536 ( .A(n12737), .Z(n12735) );
  HS65_LH_BFX4 U13537 ( .A(n12738), .Z(n12736) );
  HS65_LH_BFX4 U13538 ( .A(n12739), .Z(n12737) );
  HS65_LH_BFX4 U13539 ( .A(n12740), .Z(n12738) );
  HS65_LH_BFX4 U13540 ( .A(n12741), .Z(n12739) );
  HS65_LH_BFX4 U13541 ( .A(n12742), .Z(n12740) );
  HS65_LH_BFX4 U13542 ( .A(n12743), .Z(n12741) );
  HS65_LH_BFX4 U13543 ( .A(n12744), .Z(n12742) );
  HS65_LH_BFX4 U13544 ( .A(n12745), .Z(n12743) );
  HS65_LH_BFX4 U13545 ( .A(n12746), .Z(n12744) );
  HS65_LH_BFX4 U13546 ( .A(n12747), .Z(n12745) );
  HS65_LH_BFX4 U13547 ( .A(n12748), .Z(n12746) );
  HS65_LH_BFX4 U13548 ( .A(n12749), .Z(n12747) );
  HS65_LH_BFX4 U13549 ( .A(n12750), .Z(n12748) );
  HS65_LH_BFX4 U13550 ( .A(n12751), .Z(n12749) );
  HS65_LH_BFX4 U13551 ( .A(n12752), .Z(n12750) );
  HS65_LH_BFX4 U13552 ( .A(n12753), .Z(n12751) );
  HS65_LH_BFX4 U13553 ( .A(n12754), .Z(n12752) );
  HS65_LH_BFX4 U13554 ( .A(n12755), .Z(n12753) );
  HS65_LH_BFX4 U13555 ( .A(n12756), .Z(n12754) );
  HS65_LH_BFX4 U13556 ( .A(n12757), .Z(n12755) );
  HS65_LH_BFX4 U13557 ( .A(n12758), .Z(n12756) );
  HS65_LH_BFX4 U13558 ( .A(n15433), .Z(n12757) );
  HS65_LH_BFX4 U13559 ( .A(n12759), .Z(n12758) );
  HS65_LH_BFX4 U13560 ( .A(n12760), .Z(n12759) );
  HS65_LH_BFX4 U13561 ( .A(n12761), .Z(n12760) );
  HS65_LH_BFX4 U13562 ( .A(\u_DataPath/pc4_to_idexreg_i [5]), .Z(n12761) );
  HS65_LH_BFX4 U13563 ( .A(n17240), .Z(n12762) );
  HS65_LH_BFX4 U13564 ( .A(n12765), .Z(n12763) );
  HS65_LH_BFX4 U13565 ( .A(n12766), .Z(n12764) );
  HS65_LH_BFX4 U13566 ( .A(n12767), .Z(n12765) );
  HS65_LH_BFX4 U13567 ( .A(n12768), .Z(n12766) );
  HS65_LH_BFX4 U13568 ( .A(n12769), .Z(n12767) );
  HS65_LH_BFX4 U13569 ( .A(n12770), .Z(n12768) );
  HS65_LH_BFX4 U13570 ( .A(n12771), .Z(n12769) );
  HS65_LH_BFX4 U13571 ( .A(n12772), .Z(n12770) );
  HS65_LH_BFX4 U13572 ( .A(n12773), .Z(n12771) );
  HS65_LH_BFX4 U13573 ( .A(n12774), .Z(n12772) );
  HS65_LH_BFX4 U13574 ( .A(n12775), .Z(n12773) );
  HS65_LH_BFX4 U13575 ( .A(n12776), .Z(n12774) );
  HS65_LH_BFX4 U13576 ( .A(n12777), .Z(n12775) );
  HS65_LH_BFX4 U13577 ( .A(n12778), .Z(n12776) );
  HS65_LH_BFX4 U13578 ( .A(n12779), .Z(n12777) );
  HS65_LH_BFX4 U13579 ( .A(n12780), .Z(n12778) );
  HS65_LH_BFX4 U13580 ( .A(n12781), .Z(n12779) );
  HS65_LH_BFX4 U13581 ( .A(n12782), .Z(n12780) );
  HS65_LH_BFX4 U13582 ( .A(n12783), .Z(n12781) );
  HS65_LH_BFX4 U13583 ( .A(n12784), .Z(n12782) );
  HS65_LH_BFX4 U13584 ( .A(n12785), .Z(n12783) );
  HS65_LH_BFX4 U13585 ( .A(n12786), .Z(n12784) );
  HS65_LH_BFX4 U13586 ( .A(n12787), .Z(n12785) );
  HS65_LH_BFX4 U13587 ( .A(n12788), .Z(n12786) );
  HS65_LH_BFX4 U13588 ( .A(n12789), .Z(n12787) );
  HS65_LH_BFX4 U13589 ( .A(n12790), .Z(n12788) );
  HS65_LH_BFX4 U13590 ( .A(n12791), .Z(n12789) );
  HS65_LH_BFX4 U13591 ( .A(n12792), .Z(n12790) );
  HS65_LH_BFX4 U13592 ( .A(n12793), .Z(n12791) );
  HS65_LH_BFX4 U13593 ( .A(n12794), .Z(n12792) );
  HS65_LH_BFX4 U13594 ( .A(n12795), .Z(n12793) );
  HS65_LH_BFX4 U13595 ( .A(n12796), .Z(n12794) );
  HS65_LH_BFX4 U13596 ( .A(n12797), .Z(n12795) );
  HS65_LH_BFX4 U13597 ( .A(n12798), .Z(n12796) );
  HS65_LH_BFX4 U13598 ( .A(n12799), .Z(n12797) );
  HS65_LH_BFX4 U13599 ( .A(n12800), .Z(n12798) );
  HS65_LH_BFX4 U13600 ( .A(n12801), .Z(n12799) );
  HS65_LH_BFX4 U13601 ( .A(n14080), .Z(n12800) );
  HS65_LH_BFX4 U13602 ( .A(n12802), .Z(n12801) );
  HS65_LH_BFX4 U13603 ( .A(n12803), .Z(n12802) );
  HS65_LH_BFX4 U13604 ( .A(n12804), .Z(n12803) );
  HS65_LH_BFX4 U13605 ( .A(n12805), .Z(n12804) );
  HS65_LH_BFX4 U13606 ( .A(\u_DataPath/pc4_to_idexreg_i [6]), .Z(n12805) );
  HS65_LH_BFX4 U13607 ( .A(n17239), .Z(n12806) );
  HS65_LH_BFX4 U13608 ( .A(n12809), .Z(n12807) );
  HS65_LH_BFX4 U13609 ( .A(n12810), .Z(n12808) );
  HS65_LH_BFX4 U13610 ( .A(n12811), .Z(n12809) );
  HS65_LH_BFX4 U13611 ( .A(n12812), .Z(n12810) );
  HS65_LH_BFX4 U13612 ( .A(n12813), .Z(n12811) );
  HS65_LH_BFX4 U13613 ( .A(n12814), .Z(n12812) );
  HS65_LH_BFX4 U13614 ( .A(n12815), .Z(n12813) );
  HS65_LH_BFX4 U13615 ( .A(n12816), .Z(n12814) );
  HS65_LH_BFX4 U13616 ( .A(n12817), .Z(n12815) );
  HS65_LH_BFX4 U13617 ( .A(n12818), .Z(n12816) );
  HS65_LH_BFX4 U13618 ( .A(n12819), .Z(n12817) );
  HS65_LH_BFX4 U13619 ( .A(n12820), .Z(n12818) );
  HS65_LH_BFX4 U13620 ( .A(n12821), .Z(n12819) );
  HS65_LH_BFX4 U13621 ( .A(n12822), .Z(n12820) );
  HS65_LH_BFX4 U13622 ( .A(n12823), .Z(n12821) );
  HS65_LH_BFX4 U13623 ( .A(n12824), .Z(n12822) );
  HS65_LH_BFX4 U13624 ( .A(n12825), .Z(n12823) );
  HS65_LH_BFX4 U13625 ( .A(n12826), .Z(n12824) );
  HS65_LH_BFX4 U13626 ( .A(n12827), .Z(n12825) );
  HS65_LH_BFX4 U13627 ( .A(n12828), .Z(n12826) );
  HS65_LH_BFX4 U13628 ( .A(n12829), .Z(n12827) );
  HS65_LH_BFX4 U13629 ( .A(n12830), .Z(n12828) );
  HS65_LH_BFX4 U13630 ( .A(n12831), .Z(n12829) );
  HS65_LH_BFX4 U13631 ( .A(n12832), .Z(n12830) );
  HS65_LH_BFX4 U13632 ( .A(n12833), .Z(n12831) );
  HS65_LH_BFX4 U13633 ( .A(n12834), .Z(n12832) );
  HS65_LH_BFX4 U13634 ( .A(n12835), .Z(n12833) );
  HS65_LH_BFX4 U13635 ( .A(n12836), .Z(n12834) );
  HS65_LH_BFX4 U13636 ( .A(n12837), .Z(n12835) );
  HS65_LH_BFX4 U13637 ( .A(n12838), .Z(n12836) );
  HS65_LH_BFX4 U13638 ( .A(n12839), .Z(n12837) );
  HS65_LH_BFX4 U13639 ( .A(n12840), .Z(n12838) );
  HS65_LH_BFX4 U13640 ( .A(n12841), .Z(n12839) );
  HS65_LH_BFX4 U13641 ( .A(n12842), .Z(n12840) );
  HS65_LH_BFX4 U13642 ( .A(n12843), .Z(n12841) );
  HS65_LH_BFX4 U13643 ( .A(n12844), .Z(n12842) );
  HS65_LH_BFX4 U13644 ( .A(n12845), .Z(n12843) );
  HS65_LH_BFX4 U13645 ( .A(n12846), .Z(n12844) );
  HS65_LH_BFX4 U13646 ( .A(n12847), .Z(n12845) );
  HS65_LH_BFX4 U13647 ( .A(n15436), .Z(n12846) );
  HS65_LH_BFX4 U13648 ( .A(n12848), .Z(n12847) );
  HS65_LH_BFX4 U13649 ( .A(n12849), .Z(n12848) );
  HS65_LH_BFX4 U13650 ( .A(n12850), .Z(n12849) );
  HS65_LH_BFX4 U13651 ( .A(\u_DataPath/pc4_to_idexreg_i [7]), .Z(n12850) );
  HS65_LH_BFX4 U13652 ( .A(n12853), .Z(n12851) );
  HS65_LH_BFX4 U13653 ( .A(n12854), .Z(n12852) );
  HS65_LH_BFX4 U13654 ( .A(n12855), .Z(n12853) );
  HS65_LH_BFX4 U13655 ( .A(n12856), .Z(n12854) );
  HS65_LH_BFX4 U13656 ( .A(n12857), .Z(n12855) );
  HS65_LH_BFX4 U13657 ( .A(n12858), .Z(n12856) );
  HS65_LH_BFX4 U13658 ( .A(n12859), .Z(n12857) );
  HS65_LH_BFX4 U13659 ( .A(n12860), .Z(n12858) );
  HS65_LH_BFX4 U13660 ( .A(n12861), .Z(n12859) );
  HS65_LH_BFX4 U13661 ( .A(n12862), .Z(n12860) );
  HS65_LH_BFX4 U13662 ( .A(n12863), .Z(n12861) );
  HS65_LH_BFX4 U13663 ( .A(n12864), .Z(n12862) );
  HS65_LH_BFX4 U13664 ( .A(n12865), .Z(n12863) );
  HS65_LH_BFX4 U13665 ( .A(n12866), .Z(n12864) );
  HS65_LH_BFX4 U13666 ( .A(n12867), .Z(n12865) );
  HS65_LH_BFX4 U13667 ( .A(n12868), .Z(n12866) );
  HS65_LH_BFX4 U13668 ( .A(n12869), .Z(n12867) );
  HS65_LH_BFX4 U13669 ( .A(n12870), .Z(n12868) );
  HS65_LH_BFX4 U13670 ( .A(n12871), .Z(n12869) );
  HS65_LH_BFX4 U13671 ( .A(n12872), .Z(n12870) );
  HS65_LH_BFX4 U13672 ( .A(n12873), .Z(n12871) );
  HS65_LH_BFX4 U13673 ( .A(n12874), .Z(n12872) );
  HS65_LH_BFX4 U13674 ( .A(n12875), .Z(n12873) );
  HS65_LH_BFX4 U13675 ( .A(n12876), .Z(n12874) );
  HS65_LH_BFX4 U13676 ( .A(n12877), .Z(n12875) );
  HS65_LH_BFX4 U13677 ( .A(n12878), .Z(n12876) );
  HS65_LH_BFX4 U13678 ( .A(n12879), .Z(n12877) );
  HS65_LH_BFX4 U13679 ( .A(n12880), .Z(n12878) );
  HS65_LH_BFX4 U13680 ( .A(n12881), .Z(n12879) );
  HS65_LH_BFX4 U13681 ( .A(n12882), .Z(n12880) );
  HS65_LH_BFX4 U13682 ( .A(n12883), .Z(n12881) );
  HS65_LH_BFX4 U13683 ( .A(n12884), .Z(n12882) );
  HS65_LH_BFX4 U13684 ( .A(n12885), .Z(n12883) );
  HS65_LH_BFX4 U13685 ( .A(n12886), .Z(n12884) );
  HS65_LH_BFX4 U13686 ( .A(n12887), .Z(n12885) );
  HS65_LH_BFX4 U13687 ( .A(n12888), .Z(n12886) );
  HS65_LH_BFX4 U13688 ( .A(n12889), .Z(n12887) );
  HS65_LH_BFX4 U13689 ( .A(n12890), .Z(n12888) );
  HS65_LH_BFX4 U13690 ( .A(n12891), .Z(n12889) );
  HS65_LH_BFX4 U13691 ( .A(n12892), .Z(n12890) );
  HS65_LH_BFX4 U13692 ( .A(n14083), .Z(n12891) );
  HS65_LH_BFX4 U13693 ( .A(n12893), .Z(n12892) );
  HS65_LH_BFX4 U13694 ( .A(n12894), .Z(n12893) );
  HS65_LH_BFX4 U13695 ( .A(n12895), .Z(n12894) );
  HS65_LH_BFX4 U13696 ( .A(\u_DataPath/pc4_to_idexreg_i [8]), .Z(n12895) );
  HS65_LH_BFX4 U13697 ( .A(n17237), .Z(n12896) );
  HS65_LH_BFX4 U13698 ( .A(n12899), .Z(n12897) );
  HS65_LH_BFX4 U13699 ( .A(n12900), .Z(n12898) );
  HS65_LH_BFX4 U13700 ( .A(n12901), .Z(n12899) );
  HS65_LH_BFX4 U13701 ( .A(n12902), .Z(n12900) );
  HS65_LH_BFX4 U13702 ( .A(n12903), .Z(n12901) );
  HS65_LH_BFX4 U13703 ( .A(n12904), .Z(n12902) );
  HS65_LH_BFX4 U13704 ( .A(n12905), .Z(n12903) );
  HS65_LH_BFX4 U13705 ( .A(n12906), .Z(n12904) );
  HS65_LH_BFX4 U13706 ( .A(n12907), .Z(n12905) );
  HS65_LH_BFX4 U13707 ( .A(n12908), .Z(n12906) );
  HS65_LH_BFX4 U13708 ( .A(n12909), .Z(n12907) );
  HS65_LH_BFX4 U13709 ( .A(n12910), .Z(n12908) );
  HS65_LH_BFX4 U13710 ( .A(n12911), .Z(n12909) );
  HS65_LH_BFX4 U13711 ( .A(n12912), .Z(n12910) );
  HS65_LH_BFX4 U13712 ( .A(n12913), .Z(n12911) );
  HS65_LH_BFX4 U13713 ( .A(n12914), .Z(n12912) );
  HS65_LH_BFX4 U13714 ( .A(n12915), .Z(n12913) );
  HS65_LH_BFX4 U13715 ( .A(n12916), .Z(n12914) );
  HS65_LH_BFX4 U13716 ( .A(n12917), .Z(n12915) );
  HS65_LH_BFX4 U13717 ( .A(n12918), .Z(n12916) );
  HS65_LH_BFX4 U13718 ( .A(n12919), .Z(n12917) );
  HS65_LH_BFX4 U13719 ( .A(n12920), .Z(n12918) );
  HS65_LH_BFX4 U13720 ( .A(n12921), .Z(n12919) );
  HS65_LH_BFX4 U13721 ( .A(n12922), .Z(n12920) );
  HS65_LH_BFX4 U13722 ( .A(n12923), .Z(n12921) );
  HS65_LH_BFX4 U13723 ( .A(n12924), .Z(n12922) );
  HS65_LH_BFX4 U13724 ( .A(n12925), .Z(n12923) );
  HS65_LH_BFX4 U13725 ( .A(n12926), .Z(n12924) );
  HS65_LH_BFX4 U13726 ( .A(n12927), .Z(n12925) );
  HS65_LH_BFX4 U13727 ( .A(n12928), .Z(n12926) );
  HS65_LH_BFX4 U13728 ( .A(n12929), .Z(n12927) );
  HS65_LH_BFX4 U13729 ( .A(n12930), .Z(n12928) );
  HS65_LH_BFX4 U13730 ( .A(n12931), .Z(n12929) );
  HS65_LH_BFX4 U13731 ( .A(n12932), .Z(n12930) );
  HS65_LH_BFX4 U13732 ( .A(n12933), .Z(n12931) );
  HS65_LH_BFX4 U13733 ( .A(n12934), .Z(n12932) );
  HS65_LH_BFX4 U13734 ( .A(n12935), .Z(n12933) );
  HS65_LH_BFX4 U13735 ( .A(n12936), .Z(n12934) );
  HS65_LH_BFX4 U13736 ( .A(n12937), .Z(n12935) );
  HS65_LH_BFX4 U13737 ( .A(n15439), .Z(n12936) );
  HS65_LH_BFX4 U13738 ( .A(n12938), .Z(n12937) );
  HS65_LH_BFX4 U13739 ( .A(n12939), .Z(n12938) );
  HS65_LH_BFX4 U13740 ( .A(n12940), .Z(n12939) );
  HS65_LH_BFX4 U13741 ( .A(\u_DataPath/pc4_to_idexreg_i [9]), .Z(n12940) );
  HS65_LH_BFX4 U13742 ( .A(n12943), .Z(n12941) );
  HS65_LH_BFX4 U13743 ( .A(n12944), .Z(n12942) );
  HS65_LH_BFX4 U13744 ( .A(n12945), .Z(n12943) );
  HS65_LH_BFX4 U13745 ( .A(n12946), .Z(n12944) );
  HS65_LH_BFX4 U13746 ( .A(n12947), .Z(n12945) );
  HS65_LH_BFX4 U13747 ( .A(n12948), .Z(n12946) );
  HS65_LH_BFX4 U13748 ( .A(n12949), .Z(n12947) );
  HS65_LH_BFX4 U13749 ( .A(n12950), .Z(n12948) );
  HS65_LH_BFX4 U13750 ( .A(n12951), .Z(n12949) );
  HS65_LH_BFX4 U13751 ( .A(n12952), .Z(n12950) );
  HS65_LH_BFX4 U13752 ( .A(n12953), .Z(n12951) );
  HS65_LH_BFX4 U13753 ( .A(n12954), .Z(n12952) );
  HS65_LH_BFX4 U13754 ( .A(n12955), .Z(n12953) );
  HS65_LH_BFX4 U13755 ( .A(n12956), .Z(n12954) );
  HS65_LH_BFX4 U13756 ( .A(n12957), .Z(n12955) );
  HS65_LH_BFX4 U13757 ( .A(n12958), .Z(n12956) );
  HS65_LH_BFX4 U13758 ( .A(n12959), .Z(n12957) );
  HS65_LH_BFX4 U13759 ( .A(n12960), .Z(n12958) );
  HS65_LH_BFX4 U13760 ( .A(n12961), .Z(n12959) );
  HS65_LH_BFX4 U13761 ( .A(n12962), .Z(n12960) );
  HS65_LH_BFX4 U13762 ( .A(n12963), .Z(n12961) );
  HS65_LH_BFX4 U13763 ( .A(n12964), .Z(n12962) );
  HS65_LH_BFX4 U13764 ( .A(n12965), .Z(n12963) );
  HS65_LH_BFX4 U13765 ( .A(n12966), .Z(n12964) );
  HS65_LH_BFX4 U13766 ( .A(n12967), .Z(n12965) );
  HS65_LH_BFX4 U13767 ( .A(n12968), .Z(n12966) );
  HS65_LH_BFX4 U13768 ( .A(n12969), .Z(n12967) );
  HS65_LH_BFX4 U13769 ( .A(n12970), .Z(n12968) );
  HS65_LH_BFX4 U13770 ( .A(n12971), .Z(n12969) );
  HS65_LH_BFX4 U13771 ( .A(n12972), .Z(n12970) );
  HS65_LH_BFX4 U13772 ( .A(n12973), .Z(n12971) );
  HS65_LH_BFX4 U13773 ( .A(n12974), .Z(n12972) );
  HS65_LH_BFX4 U13774 ( .A(n12975), .Z(n12973) );
  HS65_LH_BFX4 U13775 ( .A(n12976), .Z(n12974) );
  HS65_LH_BFX4 U13776 ( .A(n12977), .Z(n12975) );
  HS65_LH_BFX4 U13777 ( .A(n12978), .Z(n12976) );
  HS65_LH_BFX4 U13778 ( .A(n12979), .Z(n12977) );
  HS65_LH_BFX4 U13779 ( .A(n12980), .Z(n12978) );
  HS65_LH_BFX4 U13780 ( .A(n12981), .Z(n12979) );
  HS65_LH_BFX4 U13781 ( .A(n12982), .Z(n12980) );
  HS65_LH_BFX4 U13782 ( .A(n14085), .Z(n12981) );
  HS65_LH_BFX4 U13783 ( .A(n12983), .Z(n12982) );
  HS65_LH_BFX4 U13784 ( .A(n12984), .Z(n12983) );
  HS65_LH_BFX4 U13785 ( .A(n12985), .Z(n12984) );
  HS65_LH_BFX4 U13786 ( .A(\u_DataPath/pc4_to_idexreg_i [10]), .Z(n12985) );
  HS65_LH_BFX4 U13787 ( .A(n17235), .Z(n12986) );
  HS65_LH_BFX4 U13788 ( .A(n12989), .Z(n12987) );
  HS65_LH_BFX4 U13789 ( .A(n12990), .Z(n12988) );
  HS65_LH_BFX4 U13790 ( .A(n12991), .Z(n12989) );
  HS65_LH_BFX4 U13791 ( .A(n12992), .Z(n12990) );
  HS65_LH_BFX4 U13792 ( .A(n12993), .Z(n12991) );
  HS65_LH_BFX4 U13793 ( .A(n12994), .Z(n12992) );
  HS65_LH_BFX4 U13794 ( .A(n12995), .Z(n12993) );
  HS65_LH_BFX4 U13795 ( .A(n12996), .Z(n12994) );
  HS65_LH_BFX4 U13796 ( .A(n12997), .Z(n12995) );
  HS65_LH_BFX4 U13797 ( .A(n12998), .Z(n12996) );
  HS65_LH_BFX4 U13798 ( .A(n12999), .Z(n12997) );
  HS65_LH_BFX4 U13799 ( .A(n13000), .Z(n12998) );
  HS65_LH_BFX4 U13800 ( .A(n13001), .Z(n12999) );
  HS65_LH_BFX4 U13801 ( .A(n13002), .Z(n13000) );
  HS65_LH_BFX4 U13802 ( .A(n13003), .Z(n13001) );
  HS65_LH_BFX4 U13803 ( .A(n13004), .Z(n13002) );
  HS65_LH_BFX4 U13804 ( .A(n13005), .Z(n13003) );
  HS65_LH_BFX4 U13805 ( .A(n13006), .Z(n13004) );
  HS65_LH_BFX4 U13806 ( .A(n13007), .Z(n13005) );
  HS65_LH_BFX4 U13807 ( .A(n13008), .Z(n13006) );
  HS65_LH_BFX4 U13808 ( .A(n13009), .Z(n13007) );
  HS65_LH_BFX4 U13809 ( .A(n13010), .Z(n13008) );
  HS65_LH_BFX4 U13810 ( .A(n13011), .Z(n13009) );
  HS65_LH_BFX4 U13811 ( .A(n13012), .Z(n13010) );
  HS65_LH_BFX4 U13812 ( .A(n13013), .Z(n13011) );
  HS65_LH_BFX4 U13813 ( .A(n13014), .Z(n13012) );
  HS65_LH_BFX4 U13814 ( .A(n13015), .Z(n13013) );
  HS65_LH_BFX4 U13815 ( .A(n13016), .Z(n13014) );
  HS65_LH_BFX4 U13816 ( .A(n13017), .Z(n13015) );
  HS65_LH_BFX4 U13817 ( .A(n13018), .Z(n13016) );
  HS65_LH_BFX4 U13818 ( .A(n13019), .Z(n13017) );
  HS65_LH_BFX4 U13819 ( .A(n13020), .Z(n13018) );
  HS65_LH_BFX4 U13820 ( .A(n13021), .Z(n13019) );
  HS65_LH_BFX4 U13821 ( .A(n13022), .Z(n13020) );
  HS65_LH_BFX4 U13822 ( .A(n13023), .Z(n13021) );
  HS65_LH_BFX4 U13823 ( .A(n13024), .Z(n13022) );
  HS65_LH_BFX4 U13824 ( .A(n13025), .Z(n13023) );
  HS65_LH_BFX4 U13825 ( .A(n13026), .Z(n13024) );
  HS65_LH_BFX4 U13826 ( .A(n13027), .Z(n13025) );
  HS65_LH_BFX4 U13827 ( .A(n15442), .Z(n13026) );
  HS65_LH_BFX4 U13828 ( .A(n13028), .Z(n13027) );
  HS65_LH_BFX4 U13829 ( .A(n13029), .Z(n13028) );
  HS65_LH_BFX4 U13830 ( .A(n13030), .Z(n13029) );
  HS65_LH_BFX4 U13831 ( .A(\u_DataPath/pc4_to_idexreg_i [11]), .Z(n13030) );
  HS65_LH_BFX4 U13832 ( .A(n13033), .Z(n13031) );
  HS65_LH_BFX4 U13833 ( .A(n13034), .Z(n13032) );
  HS65_LH_BFX4 U13834 ( .A(n13035), .Z(n13033) );
  HS65_LH_BFX4 U13835 ( .A(n13036), .Z(n13034) );
  HS65_LH_BFX4 U13836 ( .A(n13037), .Z(n13035) );
  HS65_LH_BFX4 U13837 ( .A(n13038), .Z(n13036) );
  HS65_LH_BFX4 U13838 ( .A(n13039), .Z(n13037) );
  HS65_LH_BFX4 U13839 ( .A(n13040), .Z(n13038) );
  HS65_LH_BFX4 U13840 ( .A(n13041), .Z(n13039) );
  HS65_LH_BFX4 U13841 ( .A(n13042), .Z(n13040) );
  HS65_LH_BFX4 U13842 ( .A(n13043), .Z(n13041) );
  HS65_LH_BFX4 U13843 ( .A(n13044), .Z(n13042) );
  HS65_LH_BFX4 U13844 ( .A(n13045), .Z(n13043) );
  HS65_LH_BFX4 U13845 ( .A(n13046), .Z(n13044) );
  HS65_LH_BFX4 U13846 ( .A(n13047), .Z(n13045) );
  HS65_LH_BFX4 U13847 ( .A(n13048), .Z(n13046) );
  HS65_LH_BFX4 U13848 ( .A(n13049), .Z(n13047) );
  HS65_LH_BFX4 U13849 ( .A(n13050), .Z(n13048) );
  HS65_LH_BFX4 U13850 ( .A(n13051), .Z(n13049) );
  HS65_LH_BFX4 U13851 ( .A(n13052), .Z(n13050) );
  HS65_LH_BFX4 U13852 ( .A(n13053), .Z(n13051) );
  HS65_LH_BFX4 U13853 ( .A(n13054), .Z(n13052) );
  HS65_LH_BFX4 U13854 ( .A(n13055), .Z(n13053) );
  HS65_LH_BFX4 U13855 ( .A(n13056), .Z(n13054) );
  HS65_LH_BFX4 U13856 ( .A(n13057), .Z(n13055) );
  HS65_LH_BFX4 U13857 ( .A(n13058), .Z(n13056) );
  HS65_LH_BFX4 U13858 ( .A(n13059), .Z(n13057) );
  HS65_LH_BFX4 U13859 ( .A(n13060), .Z(n13058) );
  HS65_LH_BFX4 U13860 ( .A(n13061), .Z(n13059) );
  HS65_LH_BFX4 U13861 ( .A(n13062), .Z(n13060) );
  HS65_LH_BFX4 U13862 ( .A(n13063), .Z(n13061) );
  HS65_LH_BFX4 U13863 ( .A(n13064), .Z(n13062) );
  HS65_LH_BFX4 U13864 ( .A(n13065), .Z(n13063) );
  HS65_LH_BFX4 U13865 ( .A(n13066), .Z(n13064) );
  HS65_LH_BFX4 U13866 ( .A(n13067), .Z(n13065) );
  HS65_LH_BFX4 U13867 ( .A(n13068), .Z(n13066) );
  HS65_LH_BFX4 U13868 ( .A(n13069), .Z(n13067) );
  HS65_LH_BFX4 U13869 ( .A(n13070), .Z(n13068) );
  HS65_LH_BFX4 U13870 ( .A(n13071), .Z(n13069) );
  HS65_LH_BFX4 U13871 ( .A(n13072), .Z(n13070) );
  HS65_LH_BFX4 U13872 ( .A(n14087), .Z(n13071) );
  HS65_LH_BFX4 U13873 ( .A(n13073), .Z(n13072) );
  HS65_LH_BFX4 U13874 ( .A(n13074), .Z(n13073) );
  HS65_LH_BFX4 U13875 ( .A(n13075), .Z(n13074) );
  HS65_LH_BFX4 U13876 ( .A(\u_DataPath/pc4_to_idexreg_i [12]), .Z(n13075) );
  HS65_LH_BFX4 U13877 ( .A(n17233), .Z(n13076) );
  HS65_LH_BFX4 U13878 ( .A(n13079), .Z(n13077) );
  HS65_LH_BFX4 U13879 ( .A(n13080), .Z(n13078) );
  HS65_LH_BFX4 U13880 ( .A(n13081), .Z(n13079) );
  HS65_LH_BFX4 U13881 ( .A(n13082), .Z(n13080) );
  HS65_LH_BFX4 U13882 ( .A(n13083), .Z(n13081) );
  HS65_LH_BFX4 U13883 ( .A(n13084), .Z(n13082) );
  HS65_LH_BFX4 U13884 ( .A(n13085), .Z(n13083) );
  HS65_LH_BFX4 U13885 ( .A(n13086), .Z(n13084) );
  HS65_LH_BFX4 U13886 ( .A(n13087), .Z(n13085) );
  HS65_LH_BFX4 U13887 ( .A(n13088), .Z(n13086) );
  HS65_LH_BFX4 U13888 ( .A(n13089), .Z(n13087) );
  HS65_LH_BFX4 U13889 ( .A(n13090), .Z(n13088) );
  HS65_LH_BFX4 U13890 ( .A(n13091), .Z(n13089) );
  HS65_LH_BFX4 U13891 ( .A(n13092), .Z(n13090) );
  HS65_LH_BFX4 U13892 ( .A(n13093), .Z(n13091) );
  HS65_LH_BFX4 U13893 ( .A(n13094), .Z(n13092) );
  HS65_LH_BFX4 U13894 ( .A(n13095), .Z(n13093) );
  HS65_LH_BFX4 U13895 ( .A(n13096), .Z(n13094) );
  HS65_LH_BFX4 U13896 ( .A(n13097), .Z(n13095) );
  HS65_LH_BFX4 U13897 ( .A(n13098), .Z(n13096) );
  HS65_LH_BFX4 U13898 ( .A(n13099), .Z(n13097) );
  HS65_LH_BFX4 U13899 ( .A(n13100), .Z(n13098) );
  HS65_LH_BFX4 U13900 ( .A(n13101), .Z(n13099) );
  HS65_LH_BFX4 U13901 ( .A(n13102), .Z(n13100) );
  HS65_LH_BFX4 U13902 ( .A(n13103), .Z(n13101) );
  HS65_LH_BFX4 U13903 ( .A(n13104), .Z(n13102) );
  HS65_LH_BFX4 U13904 ( .A(n13105), .Z(n13103) );
  HS65_LH_BFX4 U13905 ( .A(n13106), .Z(n13104) );
  HS65_LH_BFX4 U13906 ( .A(n13107), .Z(n13105) );
  HS65_LH_BFX4 U13907 ( .A(n13108), .Z(n13106) );
  HS65_LH_BFX4 U13908 ( .A(n13109), .Z(n13107) );
  HS65_LH_BFX4 U13909 ( .A(n13110), .Z(n13108) );
  HS65_LH_BFX4 U13910 ( .A(n13111), .Z(n13109) );
  HS65_LH_BFX4 U13911 ( .A(n13112), .Z(n13110) );
  HS65_LH_BFX4 U13912 ( .A(n13113), .Z(n13111) );
  HS65_LH_BFX4 U13913 ( .A(n13114), .Z(n13112) );
  HS65_LH_BFX4 U13914 ( .A(n13115), .Z(n13113) );
  HS65_LH_BFX4 U13915 ( .A(n13116), .Z(n13114) );
  HS65_LH_BFX4 U13916 ( .A(n13117), .Z(n13115) );
  HS65_LH_BFX4 U13917 ( .A(n15445), .Z(n13116) );
  HS65_LH_BFX4 U13918 ( .A(n13118), .Z(n13117) );
  HS65_LH_BFX4 U13919 ( .A(n13119), .Z(n13118) );
  HS65_LH_BFX4 U13920 ( .A(n13120), .Z(n13119) );
  HS65_LH_BFX4 U13921 ( .A(\u_DataPath/pc4_to_idexreg_i [13]), .Z(n13120) );
  HS65_LH_BFX4 U13922 ( .A(n13123), .Z(n13121) );
  HS65_LH_BFX4 U13923 ( .A(n13124), .Z(n13122) );
  HS65_LH_BFX4 U13924 ( .A(n13125), .Z(n13123) );
  HS65_LH_BFX4 U13925 ( .A(n13126), .Z(n13124) );
  HS65_LH_BFX4 U13926 ( .A(n13127), .Z(n13125) );
  HS65_LH_BFX4 U13927 ( .A(n13128), .Z(n13126) );
  HS65_LH_BFX4 U13928 ( .A(n13129), .Z(n13127) );
  HS65_LH_BFX4 U13929 ( .A(n13130), .Z(n13128) );
  HS65_LH_BFX4 U13930 ( .A(n13131), .Z(n13129) );
  HS65_LH_BFX4 U13931 ( .A(n13132), .Z(n13130) );
  HS65_LH_BFX4 U13932 ( .A(n13133), .Z(n13131) );
  HS65_LH_BFX4 U13933 ( .A(n13134), .Z(n13132) );
  HS65_LH_BFX4 U13934 ( .A(n13135), .Z(n13133) );
  HS65_LH_BFX4 U13935 ( .A(n13136), .Z(n13134) );
  HS65_LH_BFX4 U13936 ( .A(n13137), .Z(n13135) );
  HS65_LH_BFX4 U13937 ( .A(n13138), .Z(n13136) );
  HS65_LH_BFX4 U13938 ( .A(n13139), .Z(n13137) );
  HS65_LH_BFX4 U13939 ( .A(n13140), .Z(n13138) );
  HS65_LH_BFX4 U13940 ( .A(n13141), .Z(n13139) );
  HS65_LH_BFX4 U13941 ( .A(n13142), .Z(n13140) );
  HS65_LH_BFX4 U13942 ( .A(n13143), .Z(n13141) );
  HS65_LH_BFX4 U13943 ( .A(n13144), .Z(n13142) );
  HS65_LH_BFX4 U13944 ( .A(n13145), .Z(n13143) );
  HS65_LH_BFX4 U13945 ( .A(n13146), .Z(n13144) );
  HS65_LH_BFX4 U13946 ( .A(n13147), .Z(n13145) );
  HS65_LH_BFX4 U13947 ( .A(n13148), .Z(n13146) );
  HS65_LH_BFX4 U13948 ( .A(n13149), .Z(n13147) );
  HS65_LH_BFX4 U13949 ( .A(n13150), .Z(n13148) );
  HS65_LH_BFX4 U13950 ( .A(n13151), .Z(n13149) );
  HS65_LH_BFX4 U13951 ( .A(n13152), .Z(n13150) );
  HS65_LH_BFX4 U13952 ( .A(n13153), .Z(n13151) );
  HS65_LH_BFX4 U13953 ( .A(n13154), .Z(n13152) );
  HS65_LH_BFX4 U13954 ( .A(n13155), .Z(n13153) );
  HS65_LH_BFX4 U13955 ( .A(n13156), .Z(n13154) );
  HS65_LH_BFX4 U13956 ( .A(n13157), .Z(n13155) );
  HS65_LH_BFX4 U13957 ( .A(n13158), .Z(n13156) );
  HS65_LH_BFX4 U13958 ( .A(n13159), .Z(n13157) );
  HS65_LH_BFX4 U13959 ( .A(n13160), .Z(n13158) );
  HS65_LH_BFX4 U13960 ( .A(n13161), .Z(n13159) );
  HS65_LH_BFX4 U13961 ( .A(n13162), .Z(n13160) );
  HS65_LH_BFX4 U13962 ( .A(n14089), .Z(n13161) );
  HS65_LH_BFX4 U13963 ( .A(n13163), .Z(n13162) );
  HS65_LH_BFX4 U13964 ( .A(n13164), .Z(n13163) );
  HS65_LH_BFX4 U13965 ( .A(n13165), .Z(n13164) );
  HS65_LH_BFX4 U13966 ( .A(\u_DataPath/pc4_to_idexreg_i [14]), .Z(n13165) );
  HS65_LH_BFX4 U13967 ( .A(n17231), .Z(n13166) );
  HS65_LH_BFX4 U13968 ( .A(n13169), .Z(n13167) );
  HS65_LH_BFX4 U13969 ( .A(n13170), .Z(n13168) );
  HS65_LH_BFX4 U13970 ( .A(n13171), .Z(n13169) );
  HS65_LH_BFX4 U13971 ( .A(n13172), .Z(n13170) );
  HS65_LH_BFX4 U13972 ( .A(n13173), .Z(n13171) );
  HS65_LH_BFX4 U13973 ( .A(n13174), .Z(n13172) );
  HS65_LH_BFX4 U13974 ( .A(n13175), .Z(n13173) );
  HS65_LH_BFX4 U13975 ( .A(n13176), .Z(n13174) );
  HS65_LH_BFX4 U13976 ( .A(n13177), .Z(n13175) );
  HS65_LH_BFX4 U13977 ( .A(n13178), .Z(n13176) );
  HS65_LH_BFX4 U13978 ( .A(n13179), .Z(n13177) );
  HS65_LH_BFX4 U13979 ( .A(n13180), .Z(n13178) );
  HS65_LH_BFX4 U13980 ( .A(n13181), .Z(n13179) );
  HS65_LH_BFX4 U13981 ( .A(n13182), .Z(n13180) );
  HS65_LH_BFX4 U13982 ( .A(n13183), .Z(n13181) );
  HS65_LH_BFX4 U13983 ( .A(n13184), .Z(n13182) );
  HS65_LH_BFX4 U13984 ( .A(n13185), .Z(n13183) );
  HS65_LH_BFX4 U13985 ( .A(n13186), .Z(n13184) );
  HS65_LH_BFX4 U13986 ( .A(n13187), .Z(n13185) );
  HS65_LH_BFX4 U13987 ( .A(n13188), .Z(n13186) );
  HS65_LH_BFX4 U13988 ( .A(n13189), .Z(n13187) );
  HS65_LH_BFX4 U13989 ( .A(n13190), .Z(n13188) );
  HS65_LH_BFX4 U13990 ( .A(n13191), .Z(n13189) );
  HS65_LH_BFX4 U13991 ( .A(n13192), .Z(n13190) );
  HS65_LH_BFX4 U13992 ( .A(n13193), .Z(n13191) );
  HS65_LH_BFX4 U13993 ( .A(n13194), .Z(n13192) );
  HS65_LH_BFX4 U13994 ( .A(n13195), .Z(n13193) );
  HS65_LH_BFX4 U13995 ( .A(n13196), .Z(n13194) );
  HS65_LH_BFX4 U13996 ( .A(n13197), .Z(n13195) );
  HS65_LH_BFX4 U13997 ( .A(n13198), .Z(n13196) );
  HS65_LH_BFX4 U13998 ( .A(n13199), .Z(n13197) );
  HS65_LH_BFX4 U13999 ( .A(n13200), .Z(n13198) );
  HS65_LH_BFX4 U14000 ( .A(n13201), .Z(n13199) );
  HS65_LH_BFX4 U14001 ( .A(n13202), .Z(n13200) );
  HS65_LH_BFX4 U14002 ( .A(n13203), .Z(n13201) );
  HS65_LH_BFX4 U14003 ( .A(n13204), .Z(n13202) );
  HS65_LH_BFX4 U14004 ( .A(n13205), .Z(n13203) );
  HS65_LH_BFX4 U14005 ( .A(n13206), .Z(n13204) );
  HS65_LH_BFX4 U14006 ( .A(n13207), .Z(n13205) );
  HS65_LH_BFX4 U14007 ( .A(n15448), .Z(n13206) );
  HS65_LH_BFX4 U14008 ( .A(n13208), .Z(n13207) );
  HS65_LH_BFX4 U14009 ( .A(n13209), .Z(n13208) );
  HS65_LH_BFX4 U14010 ( .A(n13210), .Z(n13209) );
  HS65_LH_BFX4 U14011 ( .A(\u_DataPath/pc4_to_idexreg_i [15]), .Z(n13210) );
  HS65_LH_BFX4 U14012 ( .A(n13213), .Z(n13211) );
  HS65_LH_BFX4 U14013 ( .A(n13214), .Z(n13212) );
  HS65_LH_BFX4 U14014 ( .A(n13215), .Z(n13213) );
  HS65_LH_BFX4 U14015 ( .A(n13216), .Z(n13214) );
  HS65_LH_BFX4 U14016 ( .A(n13217), .Z(n13215) );
  HS65_LH_BFX4 U14017 ( .A(n13218), .Z(n13216) );
  HS65_LH_BFX4 U14018 ( .A(n13219), .Z(n13217) );
  HS65_LH_BFX4 U14019 ( .A(n13220), .Z(n13218) );
  HS65_LH_BFX4 U14020 ( .A(n13221), .Z(n13219) );
  HS65_LH_BFX4 U14021 ( .A(n13222), .Z(n13220) );
  HS65_LH_BFX4 U14022 ( .A(n13223), .Z(n13221) );
  HS65_LH_BFX4 U14023 ( .A(n13224), .Z(n13222) );
  HS65_LH_BFX4 U14024 ( .A(n13225), .Z(n13223) );
  HS65_LH_BFX4 U14025 ( .A(n13226), .Z(n13224) );
  HS65_LH_BFX4 U14026 ( .A(n13227), .Z(n13225) );
  HS65_LH_BFX4 U14027 ( .A(n13228), .Z(n13226) );
  HS65_LH_BFX4 U14028 ( .A(n13229), .Z(n13227) );
  HS65_LH_BFX4 U14029 ( .A(n13230), .Z(n13228) );
  HS65_LH_BFX4 U14030 ( .A(n13231), .Z(n13229) );
  HS65_LH_BFX4 U14031 ( .A(n13232), .Z(n13230) );
  HS65_LH_BFX4 U14032 ( .A(n13233), .Z(n13231) );
  HS65_LH_BFX4 U14033 ( .A(n13234), .Z(n13232) );
  HS65_LH_BFX4 U14034 ( .A(n13235), .Z(n13233) );
  HS65_LH_BFX4 U14035 ( .A(n13236), .Z(n13234) );
  HS65_LH_BFX4 U14036 ( .A(n13237), .Z(n13235) );
  HS65_LH_BFX4 U14037 ( .A(n13238), .Z(n13236) );
  HS65_LH_BFX4 U14038 ( .A(n13239), .Z(n13237) );
  HS65_LH_BFX4 U14039 ( .A(n13240), .Z(n13238) );
  HS65_LH_BFX4 U14040 ( .A(n13241), .Z(n13239) );
  HS65_LH_BFX4 U14041 ( .A(n13242), .Z(n13240) );
  HS65_LH_BFX4 U14042 ( .A(n13243), .Z(n13241) );
  HS65_LH_BFX4 U14043 ( .A(n13244), .Z(n13242) );
  HS65_LH_BFX4 U14044 ( .A(n13245), .Z(n13243) );
  HS65_LH_BFX4 U14045 ( .A(n13246), .Z(n13244) );
  HS65_LH_BFX4 U14046 ( .A(n13247), .Z(n13245) );
  HS65_LH_BFX4 U14047 ( .A(n13248), .Z(n13246) );
  HS65_LH_BFX4 U14048 ( .A(n13249), .Z(n13247) );
  HS65_LH_BFX4 U14049 ( .A(n13250), .Z(n13248) );
  HS65_LH_BFX4 U14050 ( .A(n13251), .Z(n13249) );
  HS65_LH_BFX4 U14051 ( .A(n13252), .Z(n13250) );
  HS65_LH_BFX4 U14052 ( .A(n14091), .Z(n13251) );
  HS65_LH_BFX4 U14053 ( .A(n13253), .Z(n13252) );
  HS65_LH_BFX4 U14054 ( .A(n13254), .Z(n13253) );
  HS65_LH_BFX4 U14055 ( .A(n13255), .Z(n13254) );
  HS65_LH_BFX4 U14056 ( .A(\u_DataPath/pc4_to_idexreg_i [16]), .Z(n13255) );
  HS65_LH_BFX4 U14057 ( .A(n17229), .Z(n13256) );
  HS65_LH_BFX4 U14058 ( .A(n13259), .Z(n13257) );
  HS65_LH_BFX4 U14060 ( .A(n13261), .Z(n13259) );
  HS65_LH_BFX4 U14061 ( .A(n13262), .Z(n13260) );
  HS65_LH_BFX4 U14062 ( .A(n13263), .Z(n13261) );
  HS65_LH_BFX4 U14063 ( .A(n13264), .Z(n13262) );
  HS65_LH_BFX4 U14064 ( .A(n13265), .Z(n13263) );
  HS65_LH_BFX4 U14065 ( .A(n13266), .Z(n13264) );
  HS65_LH_BFX4 U14066 ( .A(n13267), .Z(n13265) );
  HS65_LH_BFX4 U14067 ( .A(n13268), .Z(n13266) );
  HS65_LH_BFX4 U14068 ( .A(n13269), .Z(n13267) );
  HS65_LH_BFX4 U14069 ( .A(n13270), .Z(n13268) );
  HS65_LH_BFX4 U14070 ( .A(n13271), .Z(n13269) );
  HS65_LH_BFX4 U14071 ( .A(n13272), .Z(n13270) );
  HS65_LH_BFX4 U14072 ( .A(n13273), .Z(n13271) );
  HS65_LH_BFX4 U14073 ( .A(n13274), .Z(n13272) );
  HS65_LH_BFX4 U14074 ( .A(n13275), .Z(n13273) );
  HS65_LH_BFX4 U14075 ( .A(n13276), .Z(n13274) );
  HS65_LH_BFX4 U14076 ( .A(n13277), .Z(n13275) );
  HS65_LH_BFX4 U14077 ( .A(n13278), .Z(n13276) );
  HS65_LH_BFX4 U14078 ( .A(n13279), .Z(n13277) );
  HS65_LH_BFX4 U14079 ( .A(n13280), .Z(n13278) );
  HS65_LH_BFX4 U14080 ( .A(n13281), .Z(n13279) );
  HS65_LH_BFX4 U14081 ( .A(n13282), .Z(n13280) );
  HS65_LH_BFX4 U14082 ( .A(n13283), .Z(n13281) );
  HS65_LH_BFX4 U14083 ( .A(n13284), .Z(n13282) );
  HS65_LH_BFX4 U14084 ( .A(n13285), .Z(n13283) );
  HS65_LH_BFX4 U14085 ( .A(n13286), .Z(n13284) );
  HS65_LH_BFX4 U14086 ( .A(n13287), .Z(n13285) );
  HS65_LH_BFX4 U14087 ( .A(n13288), .Z(n13286) );
  HS65_LH_BFX4 U14088 ( .A(n13289), .Z(n13287) );
  HS65_LH_BFX4 U14089 ( .A(n13290), .Z(n13288) );
  HS65_LH_BFX4 U14090 ( .A(n13291), .Z(n13289) );
  HS65_LH_BFX4 U14091 ( .A(n13292), .Z(n13290) );
  HS65_LH_BFX4 U14092 ( .A(n13293), .Z(n13291) );
  HS65_LH_BFX4 U14093 ( .A(n13294), .Z(n13292) );
  HS65_LH_BFX4 U14094 ( .A(n13295), .Z(n13293) );
  HS65_LH_BFX4 U14095 ( .A(n13296), .Z(n13294) );
  HS65_LH_BFX4 U14096 ( .A(n13297), .Z(n13295) );
  HS65_LH_BFX4 U14097 ( .A(n15451), .Z(n13296) );
  HS65_LH_BFX4 U14098 ( .A(n13298), .Z(n13297) );
  HS65_LH_BFX4 U14099 ( .A(n13299), .Z(n13298) );
  HS65_LH_BFX4 U14100 ( .A(n13300), .Z(n13299) );
  HS65_LH_BFX4 U14101 ( .A(\u_DataPath/pc4_to_idexreg_i [17]), .Z(n13300) );
  HS65_LH_BFX4 U14103 ( .A(n13304), .Z(n13302) );
  HS65_LH_BFX4 U14105 ( .A(n13306), .Z(n13304) );
  HS65_LH_BFX4 U14107 ( .A(n13308), .Z(n13306) );
  HS65_LH_BFX4 U14109 ( .A(n13310), .Z(n13308) );
  HS65_LH_BFX4 U14111 ( .A(n13312), .Z(n13310) );
  HS65_LH_BFX4 U14112 ( .A(n13313), .Z(n13311) );
  HS65_LH_BFX4 U14113 ( .A(n13314), .Z(n13312) );
  HS65_LH_BFX4 U14114 ( .A(n13315), .Z(n13313) );
  HS65_LH_BFX4 U14115 ( .A(n13316), .Z(n13314) );
  HS65_LH_BFX4 U14116 ( .A(n13317), .Z(n13315) );
  HS65_LH_BFX4 U14117 ( .A(n13318), .Z(n13316) );
  HS65_LH_BFX4 U14118 ( .A(n13319), .Z(n13317) );
  HS65_LH_BFX4 U14119 ( .A(n13320), .Z(n13318) );
  HS65_LH_BFX4 U14120 ( .A(n13321), .Z(n13319) );
  HS65_LH_BFX4 U14121 ( .A(n13322), .Z(n13320) );
  HS65_LH_BFX4 U14122 ( .A(n13323), .Z(n13321) );
  HS65_LH_BFX4 U14123 ( .A(n13324), .Z(n13322) );
  HS65_LH_BFX4 U14124 ( .A(n13325), .Z(n13323) );
  HS65_LH_BFX4 U14125 ( .A(n13326), .Z(n13324) );
  HS65_LH_BFX4 U14126 ( .A(n13327), .Z(n13325) );
  HS65_LH_BFX4 U14127 ( .A(n13328), .Z(n13326) );
  HS65_LH_BFX4 U14128 ( .A(n13329), .Z(n13327) );
  HS65_LH_BFX4 U14129 ( .A(n13330), .Z(n13328) );
  HS65_LH_BFX4 U14130 ( .A(n13331), .Z(n13329) );
  HS65_LH_BFX4 U14131 ( .A(n13332), .Z(n13330) );
  HS65_LH_BFX4 U14132 ( .A(n13333), .Z(n13331) );
  HS65_LH_BFX4 U14133 ( .A(n13334), .Z(n13332) );
  HS65_LH_BFX4 U14134 ( .A(n13335), .Z(n13333) );
  HS65_LH_BFX4 U14135 ( .A(n13336), .Z(n13334) );
  HS65_LH_BFX4 U14136 ( .A(n13337), .Z(n13335) );
  HS65_LH_BFX4 U14137 ( .A(n13338), .Z(n13336) );
  HS65_LH_BFX4 U14138 ( .A(n13339), .Z(n13337) );
  HS65_LH_BFX4 U14139 ( .A(n13340), .Z(n13338) );
  HS65_LH_BFX4 U14140 ( .A(n13341), .Z(n13339) );
  HS65_LH_BFX4 U14141 ( .A(n13342), .Z(n13340) );
  HS65_LH_BFX4 U14142 ( .A(n14093), .Z(n13341) );
  HS65_LH_BFX4 U14143 ( .A(n13343), .Z(n13342) );
  HS65_LH_BFX4 U14144 ( .A(n13344), .Z(n13343) );
  HS65_LH_BFX4 U14145 ( .A(n13345), .Z(n13344) );
  HS65_LH_BFX4 U14146 ( .A(\u_DataPath/pc4_to_idexreg_i [18]), .Z(n13345) );
  HS65_LH_BFX4 U14147 ( .A(n17219), .Z(n13346) );
  HS65_LH_BFX4 U14148 ( .A(n13349), .Z(n13347) );
  HS65_LH_BFX4 U14150 ( .A(n13351), .Z(n13349) );
  HS65_LH_BFX4 U14152 ( .A(n13353), .Z(n13351) );
  HS65_LH_BFX4 U14154 ( .A(n13355), .Z(n13353) );
  HS65_LH_BFX4 U14156 ( .A(n13357), .Z(n13355) );
  HS65_LH_BFX4 U14158 ( .A(n13359), .Z(n13357) );
  HS65_LH_BFX4 U14160 ( .A(n13361), .Z(n13359) );
  HS65_LH_BFX4 U14162 ( .A(n13363), .Z(n13361) );
  HS65_LH_BFX4 U14164 ( .A(n13365), .Z(n13363) );
  HS65_LH_BFX4 U14166 ( .A(n13367), .Z(n13365) );
  HS65_LH_BFX4 U14168 ( .A(n13369), .Z(n13367) );
  HS65_LH_BFX4 U14170 ( .A(n13371), .Z(n13369) );
  HS65_LH_BFX4 U14172 ( .A(n13373), .Z(n13371) );
  HS65_LH_BFX4 U14174 ( .A(n13375), .Z(n13373) );
  HS65_LH_BFX4 U14176 ( .A(n13377), .Z(n13375) );
  HS65_LH_BFX4 U14178 ( .A(n13379), .Z(n13377) );
  HS65_LH_BFX4 U14180 ( .A(n13381), .Z(n13379) );
  HS65_LH_BFX4 U14182 ( .A(n13383), .Z(n13381) );
  HS65_LH_BFX4 U14184 ( .A(n13385), .Z(n13383) );
  HS65_LH_BFX4 U14186 ( .A(n13387), .Z(n13385) );
  HS65_LH_BFX4 U14188 ( .A(n13388), .Z(n13387) );
  HS65_LH_BFX4 U14189 ( .A(n13389), .Z(n13388) );
  HS65_LH_BFX4 U14190 ( .A(n13390), .Z(n13389) );
  HS65_LH_BFX4 U14191 ( .A(\u_DataPath/pc4_to_idexreg_i [27]), .Z(n13390) );
  HS65_LH_BFX4 U14193 ( .A(n13394), .Z(n13392) );
  HS65_LH_BFX4 U14195 ( .A(n13396), .Z(n13394) );
  HS65_LH_BFX4 U14197 ( .A(n13398), .Z(n13396) );
  HS65_LH_BFX4 U14199 ( .A(n13400), .Z(n13398) );
  HS65_LH_BFX4 U14201 ( .A(n13402), .Z(n13400) );
  HS65_LH_BFX4 U14203 ( .A(n13404), .Z(n13402) );
  HS65_LH_BFX4 U14205 ( .A(n13406), .Z(n13404) );
  HS65_LH_BFX4 U14207 ( .A(n13408), .Z(n13406) );
  HS65_LH_BFX4 U14209 ( .A(n13410), .Z(n13408) );
  HS65_LH_BFX4 U14211 ( .A(n13412), .Z(n13410) );
  HS65_LH_BFX4 U14213 ( .A(n13414), .Z(n13412) );
  HS65_LH_BFX4 U14215 ( .A(n13416), .Z(n13414) );
  HS65_LH_BFX4 U14217 ( .A(n13418), .Z(n13416) );
  HS65_LH_BFX4 U14219 ( .A(n13420), .Z(n13418) );
  HS65_LH_BFX4 U14221 ( .A(n13422), .Z(n13420) );
  HS65_LH_BFX4 U14223 ( .A(n13424), .Z(n13422) );
  HS65_LH_BFX4 U14225 ( .A(n13426), .Z(n13424) );
  HS65_LH_BFX4 U14227 ( .A(n13428), .Z(n13426) );
  HS65_LH_BFX4 U14229 ( .A(n13430), .Z(n13428) );
  HS65_LH_BFX4 U14231 ( .A(n13432), .Z(n13430) );
  HS65_LH_BFX4 U14233 ( .A(n13433), .Z(n13432) );
  HS65_LH_BFX4 U14234 ( .A(n13434), .Z(n13433) );
  HS65_LH_BFX4 U14235 ( .A(n13435), .Z(n13434) );
  HS65_LH_BFX4 U14236 ( .A(\u_DataPath/pc4_to_idexreg_i [28]), .Z(n13435) );
  HS65_LH_BFX4 U14237 ( .A(n17217), .Z(n13436) );
  HS65_LH_BFX4 U14238 ( .A(n13439), .Z(n13437) );
  HS65_LH_BFX4 U14240 ( .A(n13441), .Z(n13439) );
  HS65_LH_BFX4 U14242 ( .A(n13443), .Z(n13441) );
  HS65_LH_BFX4 U14244 ( .A(n13445), .Z(n13443) );
  HS65_LH_BFX4 U14246 ( .A(n13447), .Z(n13445) );
  HS65_LH_BFX4 U14248 ( .A(n13449), .Z(n13447) );
  HS65_LH_BFX4 U14250 ( .A(n13451), .Z(n13449) );
  HS65_LH_BFX4 U14252 ( .A(n13453), .Z(n13451) );
  HS65_LH_BFX4 U14254 ( .A(n13455), .Z(n13453) );
  HS65_LH_BFX4 U14256 ( .A(n13457), .Z(n13455) );
  HS65_LH_BFX4 U14258 ( .A(n13459), .Z(n13457) );
  HS65_LH_BFX4 U14260 ( .A(n13461), .Z(n13459) );
  HS65_LH_BFX4 U14262 ( .A(n13463), .Z(n13461) );
  HS65_LH_BFX4 U14264 ( .A(n13465), .Z(n13463) );
  HS65_LH_BFX4 U14266 ( .A(n13467), .Z(n13465) );
  HS65_LH_BFX4 U14268 ( .A(n13469), .Z(n13467) );
  HS65_LH_BFX4 U14270 ( .A(n13471), .Z(n13469) );
  HS65_LH_BFX4 U14272 ( .A(n13473), .Z(n13471) );
  HS65_LH_BFX4 U14274 ( .A(n13475), .Z(n13473) );
  HS65_LH_BFX4 U14276 ( .A(n13477), .Z(n13475) );
  HS65_LH_BFX4 U14278 ( .A(n13478), .Z(n13477) );
  HS65_LH_BFX4 U14279 ( .A(n13479), .Z(n13478) );
  HS65_LH_BFX4 U14280 ( .A(n13480), .Z(n13479) );
  HS65_LH_BFX4 U14281 ( .A(\u_DataPath/pc4_to_idexreg_i [29]), .Z(n13480) );
  HS65_LH_BFX4 U14283 ( .A(n13484), .Z(n13482) );
  HS65_LH_BFX4 U14285 ( .A(n13486), .Z(n13484) );
  HS65_LH_BFX4 U14287 ( .A(n13488), .Z(n13486) );
  HS65_LH_BFX4 U14289 ( .A(n13490), .Z(n13488) );
  HS65_LH_BFX4 U14291 ( .A(n13492), .Z(n13490) );
  HS65_LH_BFX4 U14293 ( .A(n13494), .Z(n13492) );
  HS65_LH_BFX4 U14295 ( .A(n13496), .Z(n13494) );
  HS65_LH_BFX4 U14297 ( .A(n13498), .Z(n13496) );
  HS65_LH_BFX4 U14299 ( .A(n13500), .Z(n13498) );
  HS65_LH_BFX4 U14301 ( .A(n13502), .Z(n13500) );
  HS65_LH_BFX4 U14303 ( .A(n13504), .Z(n13502) );
  HS65_LH_BFX4 U14305 ( .A(n13506), .Z(n13504) );
  HS65_LH_BFX4 U14307 ( .A(n13508), .Z(n13506) );
  HS65_LH_BFX4 U14309 ( .A(n13510), .Z(n13508) );
  HS65_LH_BFX4 U14311 ( .A(n13512), .Z(n13510) );
  HS65_LH_BFX4 U14313 ( .A(n13514), .Z(n13512) );
  HS65_LH_BFX4 U14315 ( .A(n13516), .Z(n13514) );
  HS65_LH_BFX4 U14317 ( .A(n13518), .Z(n13516) );
  HS65_LH_BFX4 U14319 ( .A(n13520), .Z(n13518) );
  HS65_LH_BFX4 U14321 ( .A(n13522), .Z(n13520) );
  HS65_LH_BFX4 U14323 ( .A(n13523), .Z(n13522) );
  HS65_LH_BFX4 U14324 ( .A(n13524), .Z(n13523) );
  HS65_LH_BFX4 U14325 ( .A(n13525), .Z(n13524) );
  HS65_LH_BFX4 U14326 ( .A(\u_DataPath/pc4_to_idexreg_i [30]), .Z(n13525) );
  HS65_LH_BFX4 U14327 ( .A(n11633), .Z(n13526) );
  HS65_LH_BFX4 U14328 ( .A(n10148), .Z(n13527) );
  HS65_LH_BFX4 U14329 ( .A(n10312), .Z(n13528) );
  HS65_LH_CNIVX3 U14331 ( .A(n9864), .Z(n13530) );
  HS65_LH_CNIVX3 U14332 ( .A(n13530), .Z(n13531) );
  HS65_LH_CNIVX3 U14333 ( .A(n13550), .Z(n13532) );
  HS65_LH_CNIVX3 U14334 ( .A(n13532), .Z(n13533) );
  HS65_LH_CNIVX3 U14337 ( .A(n9710), .Z(n13536) );
  HS65_LH_CNIVX3 U14338 ( .A(n13536), .Z(n13537) );
  HS65_LH_BFX4 U14339 ( .A(n11640), .Z(n13538) );
  HS65_LH_BFX4 U14340 ( .A(n12413), .Z(n13539) );
  HS65_LH_BFX4 U14341 ( .A(n13547), .Z(n13540) );
  HS65_LH_BFX4 U14342 ( .A(n13548), .Z(n13541) );
  HS65_LH_BFX4 U14343 ( .A(n13526), .Z(n13542) );
  HS65_LH_BFX4 U14347 ( .A(n13538), .Z(n13546) );
  HS65_LH_BFX4 U14348 ( .A(n13556), .Z(n13547) );
  HS65_LH_BFX4 U14349 ( .A(n13558), .Z(n13548) );
  HS65_LH_BFX4 U14350 ( .A(n13542), .Z(n13549) );
  HS65_LH_BFX4 U14351 ( .A(n13552), .Z(n13550) );
  HS65_LH_CNIVX3 U14352 ( .A(n13561), .Z(n13551) );
  HS65_LH_CNIVX3 U14353 ( .A(n13551), .Z(n13552) );
  HS65_LH_BFX4 U14357 ( .A(n13565), .Z(n13556) );
  HS65_LH_BFX4 U14358 ( .A(n13546), .Z(n13557) );
  HS65_LH_BFX4 U14359 ( .A(n13567), .Z(n13558) );
  HS65_LH_BFX4 U14360 ( .A(n13549), .Z(n13559) );
  HS65_LH_CNIVX3 U14361 ( .A(n13570), .Z(n13560) );
  HS65_LH_CNIVX3 U14362 ( .A(n13560), .Z(n13561) );
  HS65_LH_BFX4 U14366 ( .A(n13574), .Z(n13565) );
  HS65_LH_BFX4 U14367 ( .A(n13557), .Z(n13566) );
  HS65_LH_BFX4 U14368 ( .A(n13576), .Z(n13567) );
  HS65_LH_BFX4 U14369 ( .A(n13559), .Z(n13568) );
  HS65_LH_CNIVX3 U14370 ( .A(n10480), .Z(n13569) );
  HS65_LH_CNIVX3 U14371 ( .A(n13569), .Z(n13570) );
  HS65_LH_BFX4 U14375 ( .A(n13582), .Z(n13574) );
  HS65_LH_BFX4 U14376 ( .A(n13566), .Z(n13575) );
  HS65_LH_BFX4 U14377 ( .A(n13583), .Z(n13576) );
  HS65_LH_CNIVX3 U14378 ( .A(n13539), .Z(n13577) );
  HS65_LH_CNIVX3 U14379 ( .A(n13577), .Z(n13578) );
  HS65_LH_BFX4 U14380 ( .A(n13568), .Z(n13579) );
  HS65_LH_BFX4 U14383 ( .A(n13589), .Z(n13582) );
  HS65_LH_BFX4 U14384 ( .A(n15478), .Z(n13583) );
  HS65_LH_BFX4 U14385 ( .A(n13575), .Z(n13584) );
  HS65_LH_BFX4 U14386 ( .A(n10289), .Z(n13585) );
  HS65_LH_BFX4 U14387 ( .A(n13579), .Z(n13586) );
  HS65_LH_BFX4 U14388 ( .A(n11628), .Z(n13587) );
  HS65_LH_BFX4 U14390 ( .A(n13596), .Z(n13589) );
  HS65_LH_BFX4 U14391 ( .A(n13584), .Z(n13590) );
  HS65_LH_BFX4 U14392 ( .A(n13593), .Z(n13591) );
  HS65_LH_CNIVX3 U14393 ( .A(n13607), .Z(n13592) );
  HS65_LH_CNIVX3 U14394 ( .A(n13592), .Z(n13593) );
  HS65_LH_BFX4 U14395 ( .A(n13586), .Z(n13594) );
  HS65_LH_BFX4 U14397 ( .A(n13599), .Z(n13596) );
  HS65_LH_BFX4 U14398 ( .A(n13590), .Z(n13597) );
  HS65_LH_BFX4 U14400 ( .A(n13603), .Z(n13599) );
  HS65_LH_BFX4 U14401 ( .A(n13597), .Z(n13600) );
  HS65_LH_BFX4 U14402 ( .A(n13587), .Z(n13601) );
  HS65_LH_BFX4 U14404 ( .A(n13609), .Z(n13603) );
  HS65_LH_BFX4 U14405 ( .A(n13600), .Z(n13604) );
  HS65_LH_BFX4 U14406 ( .A(n13601), .Z(n13605) );
  HS65_LH_CNIVX3 U14407 ( .A(n13605), .Z(n13606) );
  HS65_LH_CNIVX3 U14408 ( .A(n13606), .Z(n13607) );
  HS65_LH_BFX4 U14410 ( .A(n13614), .Z(n13609) );
  HS65_LH_BFX4 U14411 ( .A(n13604), .Z(n13610) );
  HS65_LH_CNIVX3 U14413 ( .A(n13618), .Z(n13612) );
  HS65_LH_CNIVX3 U14414 ( .A(n13612), .Z(n13613) );
  HS65_LH_BFX4 U14415 ( .A(n13616), .Z(n13614) );
  HS65_LH_BFX4 U14417 ( .A(n13619), .Z(n13616) );
  HS65_LH_BFX4 U14419 ( .A(n13622), .Z(n13618) );
  HS65_LH_BFX4 U14420 ( .A(n13621), .Z(n13619) );
  HS65_LH_BFX4 U14422 ( .A(n13624), .Z(n13621) );
  HS65_LH_BFX4 U14423 ( .A(n13874), .Z(n13622) );
  HS65_LH_BFX4 U14425 ( .A(n13626), .Z(n13624) );
  HS65_LH_BFX4 U14427 ( .A(n13628), .Z(n13626) );
  HS65_LH_BFX4 U14429 ( .A(n13630), .Z(n13628) );
  HS65_LH_BFX4 U14431 ( .A(n13632), .Z(n13630) );
  HS65_LH_BFX4 U14433 ( .A(n13633), .Z(n13632) );
  HS65_LH_BFX4 U14434 ( .A(n13635), .Z(n13633) );
  HS65_LH_BFX4 U14436 ( .A(n13636), .Z(n13635) );
  HS65_LH_BFX4 U14437 ( .A(n13637), .Z(n13636) );
  HS65_LH_BFX4 U14438 ( .A(\u_DataPath/pc4_to_idexreg_i [31]), .Z(n13637) );
  HS65_LH_BFX4 U14440 ( .A(n10453), .Z(n13639) );
  HS65_LH_BFX4 U14441 ( .A(n13653), .Z(n13640) );
  HS65_LH_BFX4 U14442 ( .A(n13655), .Z(n13641) );
  HS65_LH_BFX4 U14443 ( .A(n13656), .Z(n13642) );
  HS65_LH_BFX4 U14444 ( .A(n12483), .Z(n13643) );
  HS65_LH_BFX4 U14445 ( .A(\u_DataPath/immediate_ext_dec_i [3]), .Z(n13644) );
  HS65_LH_BFX4 U14446 ( .A(n10450), .Z(n13645) );
  HS65_LH_BFX4 U14447 ( .A(n13659), .Z(n13646) );
  HS65_LH_BFX4 U14448 ( .A(n11915), .Z(n13647) );
  HS65_LH_BFX4 U14449 ( .A(n11919), .Z(n13648) );
  HS65_LH_BFX4 U14450 ( .A(n13662), .Z(n13649) );
  HS65_LH_BFX4 U14451 ( .A(n13663), .Z(n13650) );
  HS65_LH_BFX4 U14453 ( .A(n13665), .Z(n13652) );
  HS65_LH_BFX4 U14454 ( .A(n13666), .Z(n13653) );
  HS65_LH_BFX4 U14455 ( .A(n13667), .Z(n13654) );
  HS65_LH_BFX4 U14456 ( .A(n13670), .Z(n13655) );
  HS65_LH_BFX4 U14457 ( .A(n13671), .Z(n13656) );
  HS65_LH_BFX4 U14458 ( .A(n13644), .Z(n13657) );
  HS65_LH_BFX4 U14459 ( .A(n13645), .Z(n13658) );
  HS65_LH_BFX4 U14460 ( .A(n13672), .Z(n13659) );
  HS65_LH_BFX4 U14461 ( .A(n13647), .Z(n13660) );
  HS65_LH_BFX4 U14462 ( .A(n13648), .Z(n13661) );
  HS65_LH_BFX4 U14463 ( .A(n13675), .Z(n13662) );
  HS65_LH_BFX4 U14464 ( .A(n13676), .Z(n13663) );
  HS65_LH_BFX4 U14466 ( .A(n13678), .Z(n13665) );
  HS65_LH_BFX4 U14467 ( .A(n13679), .Z(n13666) );
  HS65_LH_BFX4 U14468 ( .A(n13680), .Z(n13667) );
  HS65_LH_BFX4 U14469 ( .A(n13657), .Z(n13668) );
  HS65_LH_BFX4 U14470 ( .A(n13658), .Z(n13669) );
  HS65_LH_BFX4 U14471 ( .A(n13684), .Z(n13670) );
  HS65_LH_BFX4 U14472 ( .A(n13685), .Z(n13671) );
  HS65_LH_BFX4 U14473 ( .A(n13683), .Z(n13672) );
  HS65_LH_BFX4 U14474 ( .A(n13660), .Z(n13673) );
  HS65_LH_BFX4 U14475 ( .A(n13661), .Z(n13674) );
  HS65_LH_BFX4 U14476 ( .A(n13688), .Z(n13675) );
  HS65_LH_BFX4 U14477 ( .A(n13689), .Z(n13676) );
  HS65_LH_BFX4 U14479 ( .A(n13691), .Z(n13678) );
  HS65_LH_BFX4 U14480 ( .A(n13692), .Z(n13679) );
  HS65_LH_BFX4 U14481 ( .A(n13693), .Z(n13680) );
  HS65_LH_BFX4 U14482 ( .A(n13668), .Z(n13681) );
  HS65_LH_BFX4 U14483 ( .A(n13669), .Z(n13682) );
  HS65_LH_BFX4 U14484 ( .A(n13696), .Z(n13683) );
  HS65_LH_BFX4 U14485 ( .A(n13698), .Z(n13684) );
  HS65_LH_BFX4 U14486 ( .A(n13699), .Z(n13685) );
  HS65_LH_BFX4 U14487 ( .A(n13673), .Z(n13686) );
  HS65_LH_BFX4 U14488 ( .A(n13674), .Z(n13687) );
  HS65_LH_BFX4 U14489 ( .A(n13701), .Z(n13688) );
  HS65_LH_BFX4 U14490 ( .A(n13702), .Z(n13689) );
  HS65_LH_BFX4 U14492 ( .A(n13704), .Z(n13691) );
  HS65_LH_BFX4 U14493 ( .A(n13705), .Z(n13692) );
  HS65_LH_BFX4 U14494 ( .A(n13706), .Z(n13693) );
  HS65_LH_BFX4 U14495 ( .A(n13681), .Z(n13694) );
  HS65_LH_BFX4 U14496 ( .A(n13682), .Z(n13695) );
  HS65_LH_BFX4 U14497 ( .A(n13709), .Z(n13696) );
  HS65_LH_BFX4 U14498 ( .A(n13686), .Z(n13697) );
  HS65_LH_BFX4 U14499 ( .A(n13711), .Z(n13698) );
  HS65_LH_BFX4 U14500 ( .A(n13712), .Z(n13699) );
  HS65_LH_BFX4 U14501 ( .A(n13687), .Z(n13700) );
  HS65_LH_BFX4 U14502 ( .A(n13714), .Z(n13701) );
  HS65_LH_BFX4 U14503 ( .A(n13715), .Z(n13702) );
  HS65_LH_BFX4 U14505 ( .A(n13717), .Z(n13704) );
  HS65_LH_BFX4 U14506 ( .A(n13718), .Z(n13705) );
  HS65_LH_BFX4 U14507 ( .A(n13719), .Z(n13706) );
  HS65_LH_BFX4 U14508 ( .A(n13694), .Z(n13707) );
  HS65_LH_BFX4 U14509 ( .A(n13695), .Z(n13708) );
  HS65_LH_BFX4 U14510 ( .A(n13722), .Z(n13709) );
  HS65_LH_BFX4 U14511 ( .A(n13697), .Z(n13710) );
  HS65_LH_BFX4 U14512 ( .A(n13724), .Z(n13711) );
  HS65_LH_BFX4 U14513 ( .A(n13725), .Z(n13712) );
  HS65_LH_BFX4 U14514 ( .A(n13700), .Z(n13713) );
  HS65_LH_BFX4 U14515 ( .A(n13726), .Z(n13714) );
  HS65_LH_BFX4 U14516 ( .A(n13728), .Z(n13715) );
  HS65_LH_BFX4 U14518 ( .A(n13730), .Z(n13717) );
  HS65_LH_BFX4 U14519 ( .A(n13731), .Z(n13718) );
  HS65_LH_BFX4 U14520 ( .A(n13732), .Z(n13719) );
  HS65_LH_BFX4 U14521 ( .A(n13707), .Z(n13720) );
  HS65_LH_BFX4 U14522 ( .A(n13708), .Z(n13721) );
  HS65_LH_BFX4 U14523 ( .A(n13735), .Z(n13722) );
  HS65_LH_BFX4 U14524 ( .A(n13710), .Z(n13723) );
  HS65_LH_BFX4 U14525 ( .A(n13738), .Z(n13724) );
  HS65_LH_BFX4 U14526 ( .A(n13739), .Z(n13725) );
  HS65_LH_BFX4 U14527 ( .A(n13737), .Z(n13726) );
  HS65_LH_BFX4 U14528 ( .A(n13713), .Z(n13727) );
  HS65_LH_BFX4 U14529 ( .A(n13741), .Z(n13728) );
  HS65_LH_BFX4 U14531 ( .A(n13743), .Z(n13730) );
  HS65_LH_BFX4 U14532 ( .A(n13744), .Z(n13731) );
  HS65_LH_BFX4 U14533 ( .A(n13745), .Z(n13732) );
  HS65_LH_BFX4 U14534 ( .A(n13720), .Z(n13733) );
  HS65_LH_BFX4 U14535 ( .A(n13721), .Z(n13734) );
  HS65_LH_BFX4 U14536 ( .A(n13748), .Z(n13735) );
  HS65_LH_BFX4 U14537 ( .A(n13723), .Z(n13736) );
  HS65_LH_BFX4 U14538 ( .A(n13750), .Z(n13737) );
  HS65_LH_BFX4 U14539 ( .A(n13751), .Z(n13738) );
  HS65_LH_BFX4 U14540 ( .A(n13752), .Z(n13739) );
  HS65_LH_BFX4 U14541 ( .A(n13727), .Z(n13740) );
  HS65_LH_BFX4 U14542 ( .A(n13753), .Z(n13741) );
  HS65_LH_BFX4 U14544 ( .A(n13756), .Z(n13743) );
  HS65_LH_BFX4 U14545 ( .A(n13757), .Z(n13744) );
  HS65_LH_BFX4 U14546 ( .A(n13758), .Z(n13745) );
  HS65_LH_BFX4 U14547 ( .A(n13733), .Z(n13746) );
  HS65_LH_BFX4 U14548 ( .A(n13734), .Z(n13747) );
  HS65_LH_BFX4 U14549 ( .A(n13762), .Z(n13748) );
  HS65_LH_BFX4 U14550 ( .A(n13736), .Z(n13749) );
  HS65_LH_BFX4 U14551 ( .A(n13763), .Z(n13750) );
  HS65_LH_BFX4 U14552 ( .A(n13766), .Z(n13751) );
  HS65_LH_BFX4 U14553 ( .A(n13767), .Z(n13752) );
  HS65_LH_BFX4 U14554 ( .A(n13764), .Z(n13753) );
  HS65_LH_BFX4 U14556 ( .A(n13740), .Z(n13755) );
  HS65_LH_BFX4 U14557 ( .A(n13768), .Z(n13756) );
  HS65_LH_BFX4 U14558 ( .A(n13770), .Z(n13757) );
  HS65_LH_BFX4 U14559 ( .A(n13771), .Z(n13758) );
  HS65_LH_BFX4 U14560 ( .A(n13746), .Z(n13759) );
  HS65_LH_BFX4 U14561 ( .A(n13749), .Z(n13760) );
  HS65_LH_BFX4 U14562 ( .A(n13747), .Z(n13761) );
  HS65_LH_BFX4 U14563 ( .A(n13775), .Z(n13762) );
  HS65_LH_BFX4 U14564 ( .A(n13776), .Z(n13763) );
  HS65_LH_BFX4 U14565 ( .A(n13777), .Z(n13764) );
  HS65_LH_BFX4 U14567 ( .A(n13780), .Z(n13766) );
  HS65_LH_BFX4 U14568 ( .A(n13781), .Z(n13767) );
  HS65_LH_BFX4 U14569 ( .A(n13779), .Z(n13768) );
  HS65_LH_BFX4 U14570 ( .A(n13755), .Z(n13769) );
  HS65_LH_BFX4 U14571 ( .A(n13783), .Z(n13770) );
  HS65_LH_BFX4 U14572 ( .A(n13784), .Z(n13771) );
  HS65_LH_BFX4 U14573 ( .A(n13759), .Z(n13772) );
  HS65_LH_BFX4 U14574 ( .A(n13760), .Z(n13773) );
  HS65_LH_BFX4 U14575 ( .A(n13761), .Z(n13774) );
  HS65_LH_BFX4 U14576 ( .A(n13788), .Z(n13775) );
  HS65_LH_BFX4 U14577 ( .A(n13789), .Z(n13776) );
  HS65_LH_BFX4 U14578 ( .A(n13790), .Z(n13777) );
  HS65_LH_BFX4 U14580 ( .A(n13792), .Z(n13779) );
  HS65_LH_BFX4 U14581 ( .A(n13793), .Z(n13780) );
  HS65_LH_BFX4 U14582 ( .A(n13794), .Z(n13781) );
  HS65_LH_BFX4 U14583 ( .A(n13769), .Z(n13782) );
  HS65_LH_BFX4 U14584 ( .A(n13796), .Z(n13783) );
  HS65_LH_BFX4 U14585 ( .A(n13797), .Z(n13784) );
  HS65_LH_BFX4 U14586 ( .A(n13772), .Z(n13785) );
  HS65_LH_BFX4 U14587 ( .A(n13773), .Z(n13786) );
  HS65_LH_BFX4 U14588 ( .A(n13774), .Z(n13787) );
  HS65_LH_BFX4 U14589 ( .A(n13802), .Z(n13788) );
  HS65_LH_BFX4 U14590 ( .A(n13801), .Z(n13789) );
  HS65_LH_BFX4 U14591 ( .A(n13803), .Z(n13790) );
  HS65_LH_BFX4 U14593 ( .A(n13805), .Z(n13792) );
  HS65_LH_BFX4 U14594 ( .A(n13806), .Z(n13793) );
  HS65_LH_BFX4 U14595 ( .A(n13807), .Z(n13794) );
  HS65_LH_BFX4 U14596 ( .A(n13782), .Z(n13795) );
  HS65_LH_BFX4 U14597 ( .A(n13809), .Z(n13796) );
  HS65_LH_BFX4 U14598 ( .A(n13810), .Z(n13797) );
  HS65_LH_BFX4 U14599 ( .A(n13785), .Z(n13798) );
  HS65_LH_BFX4 U14600 ( .A(n13786), .Z(n13799) );
  HS65_LH_BFX4 U14601 ( .A(n13787), .Z(n13800) );
  HS65_LH_BFX4 U14602 ( .A(n13813), .Z(n13801) );
  HS65_LH_BFX4 U14603 ( .A(n13815), .Z(n13802) );
  HS65_LH_BFX4 U14604 ( .A(n13816), .Z(n13803) );
  HS65_LH_BFX4 U14606 ( .A(n13818), .Z(n13805) );
  HS65_LH_BFX4 U14607 ( .A(n13819), .Z(n13806) );
  HS65_LH_BFX4 U14608 ( .A(n13820), .Z(n13807) );
  HS65_LH_BFX4 U14609 ( .A(n13795), .Z(n13808) );
  HS65_LH_BFX4 U14610 ( .A(n13822), .Z(n13809) );
  HS65_LH_BFX4 U14611 ( .A(n13823), .Z(n13810) );
  HS65_LH_BFX4 U14612 ( .A(n13798), .Z(n13811) );
  HS65_LH_BFX4 U14613 ( .A(n13799), .Z(n13812) );
  HS65_LH_BFX4 U14614 ( .A(n13826), .Z(n13813) );
  HS65_LH_BFX4 U14615 ( .A(n13800), .Z(n13814) );
  HS65_LH_BFX4 U14616 ( .A(n13831), .Z(n13815) );
  HS65_LH_BFX4 U14617 ( .A(n13827), .Z(n13816) );
  HS65_LH_BFX4 U14619 ( .A(n13830), .Z(n13818) );
  HS65_LH_BFX4 U14620 ( .A(n13832), .Z(n13819) );
  HS65_LH_BFX4 U14621 ( .A(n13833), .Z(n13820) );
  HS65_LH_BFX4 U14622 ( .A(n13808), .Z(n13821) );
  HS65_LH_BFX4 U14623 ( .A(n13835), .Z(n13822) );
  HS65_LH_BFX4 U14624 ( .A(n13836), .Z(n13823) );
  HS65_LH_BFX4 U14625 ( .A(n13811), .Z(n13824) );
  HS65_LH_BFX4 U14626 ( .A(n13812), .Z(n13825) );
  HS65_LH_BFX4 U14627 ( .A(n13839), .Z(n13826) );
  HS65_LH_BFX4 U14628 ( .A(n13842), .Z(n13827) );
  HS65_LH_BFX4 U14629 ( .A(n13814), .Z(n13828) );
  HS65_LH_BFX4 U14631 ( .A(n13841), .Z(n13830) );
  HS65_LH_BFX4 U14632 ( .A(n13844), .Z(n13831) );
  HS65_LH_BFX4 U14633 ( .A(n13845), .Z(n13832) );
  HS65_LH_BFX4 U14634 ( .A(n13846), .Z(n13833) );
  HS65_LH_BFX4 U14635 ( .A(n13821), .Z(n13834) );
  HS65_LH_BFX4 U14636 ( .A(n13847), .Z(n13835) );
  HS65_LH_BFX4 U14637 ( .A(n13848), .Z(n13836) );
  HS65_LH_BFX4 U14638 ( .A(n13824), .Z(n13837) );
  HS65_LH_BFX4 U14639 ( .A(n13825), .Z(n13838) );
  HS65_LH_BFX4 U14640 ( .A(n13852), .Z(n13839) );
  HS65_LH_BFX4 U14642 ( .A(n13854), .Z(n13841) );
  HS65_LH_BFX4 U14643 ( .A(n13855), .Z(n13842) );
  HS65_LH_BFX4 U14644 ( .A(n13828), .Z(n13843) );
  HS65_LH_BFX4 U14645 ( .A(n13857), .Z(n13844) );
  HS65_LH_BFX4 U14646 ( .A(n13860), .Z(n13845) );
  HS65_LH_BFX4 U14647 ( .A(n13861), .Z(n13846) );
  HS65_LH_BFX4 U14648 ( .A(n13858), .Z(n13847) );
  HS65_LH_BFX4 U14649 ( .A(n13859), .Z(n13848) );
  HS65_LH_BFX4 U14650 ( .A(n13834), .Z(n13849) );
  HS65_LH_BFX4 U14651 ( .A(n13837), .Z(n13850) );
  HS65_LH_BFX4 U14652 ( .A(n13838), .Z(n13851) );
  HS65_LH_BFX4 U14653 ( .A(n13865), .Z(n13852) );
  HS65_LH_BFX4 U14655 ( .A(n13867), .Z(n13854) );
  HS65_LH_BFX4 U14656 ( .A(n13868), .Z(n13855) );
  HS65_LH_BFX4 U14657 ( .A(n13843), .Z(n13856) );
  HS65_LH_BFX4 U14658 ( .A(n13870), .Z(n13857) );
  HS65_LH_BFX4 U14659 ( .A(n12488), .Z(n13858) );
  HS65_LH_BFX4 U14660 ( .A(n13873), .Z(n13859) );
  HS65_LH_BFX4 U14661 ( .A(n13871), .Z(n13860) );
  HS65_LH_BFX4 U14662 ( .A(n13872), .Z(n13861) );
  HS65_LH_BFX4 U14663 ( .A(n13850), .Z(n13862) );
  HS65_LH_BFX4 U14664 ( .A(n13849), .Z(n13863) );
  HS65_LH_BFX4 U14665 ( .A(n13851), .Z(n13864) );
  HS65_LH_BFX4 U14666 ( .A(n13880), .Z(n13865) );
  HS65_LH_BFX4 U14668 ( .A(n13881), .Z(n13867) );
  HS65_LH_BFX4 U14669 ( .A(n13882), .Z(n13868) );
  HS65_LH_BFX4 U14670 ( .A(n13856), .Z(n13869) );
  HS65_LH_BFX4 U14671 ( .A(n14044), .Z(n13870) );
  HS65_LH_BFX4 U14672 ( .A(n11648), .Z(n13871) );
  HS65_LH_BFX4 U14673 ( .A(n9478), .Z(n13872) );
  HS65_LH_BFX4 U14674 ( .A(n13643), .Z(n13873) );
  HS65_LH_BFX4 U14675 ( .A(n13610), .Z(n13874) );
  HS65_LH_BFX4 U14676 ( .A(n13862), .Z(n13875) );
  HS65_LH_BFX4 U14677 ( .A(n13863), .Z(n13876) );
  HS65_LH_BFX4 U14678 ( .A(n13864), .Z(n13877) );
  HS65_LH_CNIVX3 U14679 ( .A(n13869), .Z(n13878) );
  HS65_LH_CNIVX3 U14680 ( .A(n13878), .Z(n13879) );
  HS65_LH_BFX4 U14681 ( .A(n11643), .Z(n13880) );
  HS65_LH_BFX4 U14682 ( .A(opcode_i[4]), .Z(n13881) );
  HS65_LH_BFX4 U14683 ( .A(n14060), .Z(n13882) );
  HS65_LH_BFX4 U14684 ( .A(n13875), .Z(n13883) );
  HS65_LH_CNIVX3 U14685 ( .A(n13877), .Z(n13884) );
  HS65_LH_CNIVX3 U14686 ( .A(n13884), .Z(n13885) );
  HS65_LH_CNIVX3 U14687 ( .A(n13876), .Z(n13886) );
  HS65_LH_CNIVX3 U14688 ( .A(n13886), .Z(n13887) );
  HS65_LH_BFX4 U14689 ( .A(n13883), .Z(n13888) );
  HS65_LH_CNIVX3 U14690 ( .A(n13888), .Z(n13889) );
  HS65_LH_CNIVX3 U14691 ( .A(n13889), .Z(n13890) );
  HS65_LH_IVX13 U14693 ( .A(n14027), .Z(n13893) );
  HS65_LH_IVX2 U14694 ( .A(n15069), .Z(n15245) );
  HS65_LH_NOR2X2 U14695 ( .A(n15789), .B(n15787), .Z(n16359) );
  HS65_LL_NAND2X7 U14696 ( .A(n15168), .B(n1113), .Z(n16503) );
  HS65_LH_NOR2X2 U14697 ( .A(n15781), .B(n15780), .Z(n16460) );
  HS65_LH_NOR2X2 U14698 ( .A(n15772), .B(n15781), .Z(n16399) );
  HS65_LH_NOR2X2 U14699 ( .A(n15772), .B(n15789), .Z(n16341) );
  HS65_LL_NAND2X7 U14700 ( .A(n12291), .B(n1912), .Z(n15786) );
  HS65_LH_NOR2X2 U14701 ( .A(n16490), .B(n16497), .Z(n17164) );
  HS65_LH_IVX13 U14702 ( .A(n15651), .Z(n13941) );
  HS65_LL_NAND2X7 U14703 ( .A(n13578), .B(n1113), .Z(n16505) );
  HS65_LH_NOR2X2 U14704 ( .A(n16488), .B(n16497), .Z(n17091) );
  HS65_LH_IVX13 U14705 ( .A(n12762), .Z(n13971) );
  HS65_LH_IVX13 U14706 ( .A(n4273), .Z(n13973) );
  HS65_LH_IVX13 U14707 ( .A(n17242), .Z(n13975) );
  HS65_LH_IVX13 U14708 ( .A(n17236), .Z(n13977) );
  HS65_LH_IVX13 U14709 ( .A(n17238), .Z(n13979) );
  HS65_LH_IVX13 U14710 ( .A(n17232), .Z(n13981) );
  HS65_LH_IVX13 U14711 ( .A(n17234), .Z(n13983) );
  HS65_LH_IVX13 U14712 ( .A(n17228), .Z(n13985) );
  HS65_LH_IVX13 U14713 ( .A(n17230), .Z(n13987) );
  HS65_LH_IVX13 U14714 ( .A(n17224), .Z(n13989) );
  HS65_LH_IVX13 U14715 ( .A(n17226), .Z(n13991) );
  HS65_LH_IVX13 U14716 ( .A(n17220), .Z(n13993) );
  HS65_LH_IVX13 U14717 ( .A(n17222), .Z(n13995) );
  HS65_LH_IVX13 U14718 ( .A(n17216), .Z(n13997) );
  HS65_LH_IVX13 U14719 ( .A(n17218), .Z(n13999) );
  HS65_LL_NAND3X5 U14720 ( .A(n15711), .B(n15714), .C(n15713), .Z(n105) );
  HS65_LL_OAI21X18 U14721 ( .A(n17324), .B(n99), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N131 ) );
  HS65_LL_OAI21X18 U14722 ( .A(n17324), .B(n101), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N139 ) );
  HS65_LL_IVX27 U14723 ( .A(n14005), .Z(addr_to_iram_0) );
  HS65_LL_OAI21X18 U14725 ( .A(n17323), .B(n104), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N141 ) );
  HS65_LL_OAI21X18 U14726 ( .A(n17323), .B(n101), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N133 ) );
  HS65_LL_OAI21X18 U14727 ( .A(n99), .B(n17323), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N125 ) );
  HS65_LL_OAI21X18 U14728 ( .A(n17323), .B(n113), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N149 ) );
  HS65_LL_NAND3X5 U14729 ( .A(n15711), .B(
        \u_DataPath/regfile_addr_out_towb_i [2]), .C(n15710), .Z(n108) );
  HS65_LL_OAI21X18 U14730 ( .A(n17322), .B(n113), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N153 ) );
  HS65_LL_OAI21X18 U14731 ( .A(n17322), .B(n101), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N137 ) );
  HS65_LL_OAI21X18 U14732 ( .A(n17322), .B(n104), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N145 ) );
  HS65_LL_OAI21X12 U14733 ( .A(n99), .B(n17322), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N129 ) );
  HS65_LL_NAND3X5 U14734 ( .A(n15711), .B(n15713), .C(n15710), .Z(n112) );
  HS65_LL_NOR2AX25 U14735 ( .A(\u_DataPath/mem_writedata_out_i [28]), .B(
        n14072), .Z(\Data_in[28]_snps_wire ) );
  HS65_LL_OAI21X12 U14736 ( .A(n99), .B(n17321), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N130 ) );
  HS65_LL_OAI21X12 U14737 ( .A(n17321), .B(n113), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N154 ) );
  HS65_LL_OAI21X18 U14738 ( .A(n17321), .B(n101), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N138 ) );
  HS65_LL_OAI21X18 U14739 ( .A(n17321), .B(n104), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N146 ) );
  HS65_LL_NAND3X5 U14740 ( .A(n15714), .B(n15713), .C(n15712), .Z(n114) );
  HS65_LL_IVX2 U14741 ( .A(n15151), .Z(n15522) );
  HS65_LL_NOR2AX25 U14742 ( .A(\u_DataPath/mem_writedata_out_i [31]), .B(
        n14072), .Z(\Data_in[31]_snps_wire ) );
  HS65_LL_AND2ABX18 U14743 ( .A(n15700), .B(n15662), .Z(
        \Address_toRAM[8]_snps_wire ) );
  HS65_LL_OAI21X12 U14744 ( .A(n17320), .B(n104), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N140 ) );
  HS65_LL_OAI21X12 U14745 ( .A(n17320), .B(n113), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N148 ) );
  HS65_LL_OAI21X18 U14746 ( .A(n17320), .B(n99), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N92 ) );
  HS65_LL_OAI21X18 U14747 ( .A(n17320), .B(n101), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N132 ) );
  HS65_LL_NAND3X5 U14748 ( .A(n15712), .B(n15710), .C(n15669), .Z(n107) );
  HS65_LL_OAI21X12 U14749 ( .A(n17325), .B(n104), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N142 ) );
  HS65_LL_OAI21X12 U14750 ( .A(n17325), .B(n113), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N150 ) );
  HS65_LL_OAI21X12 U14751 ( .A(n17325), .B(n101), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N134 ) );
  HS65_LL_OAI21X12 U14752 ( .A(n99), .B(n17325), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N126 ) );
  HS65_LL_NOR2AX25 U14753 ( .A(\u_DataPath/mem_writedata_out_i [27]), .B(
        n14072), .Z(\Data_in[27]_snps_wire ) );
  HS65_LL_OR3ABCX35 U14754 ( .A(n14077), .B(n14070), .C(n14048), .Z(n14072) );
  HS65_LH_IVX13 U14755 ( .A(n15705), .Z(n14010) );
  HS65_LL_OAI21X12 U14756 ( .A(n17319), .B(n101), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N135 ) );
  HS65_LL_OAI21X12 U14757 ( .A(n99), .B(n17319), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N127 ) );
  HS65_LL_OAI21X12 U14758 ( .A(n17319), .B(n113), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N151 ) );
  HS65_LL_OAI21X12 U14759 ( .A(n17319), .B(n104), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N143 ) );
  HS65_LL_NAND3X5 U14760 ( .A(\u_DataPath/regfile_addr_out_towb_i [2]), .B(
        n15711), .C(n15714), .Z(n110) );
  HS65_LH_IVX13 U14761 ( .A(n15674), .Z(n14012) );
  HS65_LH_IVX13 U14762 ( .A(n15692), .Z(n14014) );
  HS65_LH_IVX13 U14763 ( .A(n15687), .Z(n14016) );
  HS65_LH_IVX13 U14764 ( .A(n15690), .Z(n14018) );
  HS65_LH_IVX13 U14765 ( .A(n15693), .Z(n14020) );
  HS65_LH_IVX13 U14766 ( .A(n15695), .Z(n14022) );
  HS65_LH_IVX13 U14767 ( .A(n15691), .Z(n14024) );
  HS65_LL_NOR2X6 U14768 ( .A(\u_DataPath/cw_towb_i [1]), .B(n9540), .Z(n1907)
         );
  HS65_LL_NAND2X7 U14769 ( .A(n12382), .B(n15168), .Z(n16507) );
  HS65_LL_NOR2X6 U14770 ( .A(n16507), .B(n16508), .Z(n17131) );
  HS65_LL_NOR2X6 U14771 ( .A(n16503), .B(n16508), .Z(n17182) );
  HS65_LL_NAND2X7 U14772 ( .A(n14966), .B(n15411), .Z(n15414) );
  HS65_LH_CNIVX3 U14773 ( .A(n10719), .Z(n14047) );
  HS65_LH_CNIVX3 U14774 ( .A(n10683), .Z(n14048) );
  HS65_LH_OA12X4 U14775 ( .A(n15449), .B(addr_to_iram_16), .C(n15453), .Z(
        n14093) );
  HS65_LH_IVX2 U14776 ( .A(n14880), .Z(n14559) );
  HS65_LH_OA12X4 U14777 ( .A(n15440), .B(addr_to_iram_10), .C(n15444), .Z(
        n14087) );
  HS65_LH_IVX2 U14778 ( .A(n14730), .Z(n14734) );
  HS65_LH_IVX2 U14779 ( .A(n14843), .Z(n14627) );
  HS65_LH_OA12X4 U14780 ( .A(n14799), .B(n6703), .C(n14450), .Z(n14451) );
  HS65_LH_OA12X4 U14781 ( .A(n15437), .B(addr_to_iram_8), .C(n15441), .Z(
        n14085) );
  HS65_LH_OA12X4 U14782 ( .A(n14963), .B(n8363), .C(n14962), .Z(n14964) );
  HS65_LH_OA12X4 U14783 ( .A(n15434), .B(addr_to_iram_6), .C(n15438), .Z(
        n14083) );
  HS65_LH_OA12X4 U14784 ( .A(n15431), .B(n14059), .C(n15435), .Z(n14080) );
  HS65_LH_OA12X4 U14785 ( .A(n15160), .B(n9020), .C(n15159), .Z(n15161) );
  HS65_LH_AOI21X2 U14786 ( .A(n14941), .B(n14720), .C(n15160), .Z(n14721) );
  HS65_LH_CB4I1X4 U14787 ( .A(\u_DataPath/pc_4_to_ex_i [3]), .B(n8860), .C(
        \u_DataPath/pc_4_to_ex_i [4]), .D(n14941), .Z(n14942) );
  HS65_LH_CNIVX3 U14788 ( .A(\u_DataPath/dataOut_exe_i [8]), .Z(n15646) );
  HS65_LH_CNIVX3 U14789 ( .A(n6170), .Z(n15698) );
  HS65_LH_BFX4 U14790 ( .A(n12425), .Z(n14056) );
  HS65_LH_BFX4 U14791 ( .A(n12381), .Z(n14055) );
  HS65_LH_BFX4 U14792 ( .A(n12452), .Z(n14057) );
  HS65_LH_BFX4 U14793 ( .A(\u_DataPath/jaddr_i [19]), .Z(n14054) );
  HS65_LH_BFX4 U14794 ( .A(n12479), .Z(n14058) );
  HS65_LH_BFX4 U14795 ( .A(n10379), .Z(n14045) );
  HS65_LH_BFX4 U14796 ( .A(n10749), .Z(n14038) );
  HS65_LH_BFX4 U14797 ( .A(n12290), .Z(n14052) );
  HS65_LH_OAI211X1 U14798 ( .A(n14534), .B(n15080), .C(n14316), .D(n14327), 
        .Z(n15556) );
  HS65_LH_OA12X4 U14800 ( .A(n14654), .B(n17549), .C(n15388), .Z(n14510) );
  HS65_LH_OAI211X1 U14801 ( .A(n15386), .B(n17472), .C(n15384), .D(n15383), 
        .Z(n15542) );
  HS65_LH_OA12X4 U14802 ( .A(n14875), .B(n17914), .C(n14874), .Z(n14876) );
  HS65_LH_OA12X4 U14803 ( .A(n14748), .B(n17963), .C(n14481), .Z(n14482) );
  HS65_LH_OAI211X1 U14804 ( .A(n33728), .B(n15214), .C(n14939), .D(n14938), 
        .Z(n15541) );
  HS65_LH_CBI4I1X3 U14805 ( .A(n14428), .B(n17638), .C(n15196), .D(n14427), 
        .Z(n15537) );
  HS65_LH_OA12X4 U14806 ( .A(n14839), .B(n17543), .C(n14838), .Z(n14840) );
  HS65_LH_OA12X4 U14807 ( .A(n14906), .B(n17906), .C(n14905), .Z(n14907) );
  HS65_LH_OA12X4 U14808 ( .A(n14988), .B(n17892), .C(n14987), .Z(n14989) );
  HS65_LH_OA12X4 U14809 ( .A(n17465), .B(n17872), .C(n15122), .Z(n15124) );
  HS65_LH_OA12X4 U14810 ( .A(n15015), .B(\u_DataPath/pc_4_to_ex_i [16]), .C(
        n15053), .Z(n15016) );
  HS65_LH_OA12X4 U14811 ( .A(n14604), .B(n6189), .C(n14329), .Z(n14307) );
  HS65_LH_IVX2 U14812 ( .A(n14921), .Z(n14918) );
  HS65_LH_OA12X4 U14813 ( .A(n14542), .B(\u_DataPath/pc_4_to_ex_i [12]), .C(
        n14606), .Z(n14543) );
  HS65_LH_IVX2 U14814 ( .A(n14550), .Z(n14997) );
  HS65_LH_IVX2 U14815 ( .A(n15099), .Z(n15096) );
  HS65_LH_IVX2 U14816 ( .A(n14494), .Z(n14642) );
  HS65_LH_IVX2 U14817 ( .A(n14817), .Z(n14822) );
  HS65_LH_AOI21X2 U14818 ( .A(n14450), .B(n14356), .C(n14542), .Z(n14357) );
  HS65_LH_IVX2 U14819 ( .A(n17253), .Z(n14033) );
  HS65_LH_IVX2 U14820 ( .A(n17256), .Z(n14545) );
  HS65_LH_IVX2 U14821 ( .A(n17252), .Z(n14358) );
  HS65_LH_AOI21X2 U14822 ( .A(n14962), .B(n14800), .C(n14799), .Z(n14801) );
  HS65_LH_OAI212X3 U14823 ( .A(n17492), .B(n40255), .C(n17624), .D(n17728), 
        .E(n15482), .Z(n15483) );
  HS65_LH_AOI21X2 U14824 ( .A(n15159), .B(n14576), .C(n14963), .Z(n14577) );
  HS65_LH_AOI21X2 U14825 ( .A(n15641), .B(n14111), .C(n15640), .Z(n15642) );
  HS65_LH_AOI21X2 U14826 ( .A(n14111), .B(n15165), .C(n15164), .Z(n15166) );
  HS65_LH_AOI21X2 U14827 ( .A(n15432), .B(n4322), .C(n15431), .Z(n15433) );
  HS65_LH_CNIVX3 U14828 ( .A(\u_DataPath/dataOut_exe_i [20]), .Z(n15697) );
  HS65_LH_IVX2 U14829 ( .A(\u_DataPath/dataOut_exe_i [25]), .Z(n14747) );
  HS65_LH_CNIVX3 U14831 ( .A(addr_to_iram_23), .Z(n14100) );
  HS65_LH_CNIVX3 U14832 ( .A(addr_to_iram_21), .Z(n14098) );
  HS65_LH_BFX4 U14833 ( .A(\u_DataPath/cw_to_ex_i [15]), .Z(n14049) );
  HS65_LH_CNIVX3 U14834 ( .A(addr_to_iram_19), .Z(n14096) );
  HS65_LH_CNIVX3 U14835 ( .A(n13594), .Z(n14046) );
  HS65_LH_CNIVX3 U14836 ( .A(addr_to_iram_27), .Z(n14104) );
  HS65_LH_CNIVX3 U14837 ( .A(addr_to_iram_25), .Z(n14102) );
  HS65_LH_BFX4 U14838 ( .A(\u_DataPath/u_idexreg/N21 ), .Z(n14043) );
  HS65_LH_BFX4 U14839 ( .A(n10446), .Z(n14060) );
  HS65_LH_CNIVX3 U14840 ( .A(addr_to_iram_17), .Z(n14094) );
  HS65_LH_OAI211X1 U14841 ( .A(n14873), .B(n14872), .C(n14871), .D(n14870), 
        .Z(n15568) );
  HS65_LH_NAND3X2 U14842 ( .A(n14508), .B(n14500), .C(n14507), .Z(n15567) );
  HS65_LH_AOI211X1 U14843 ( .A(n14930), .B(n14869), .C(n14575), .D(n14574), 
        .Z(n15548) );
  HS65_LH_AOI21X2 U14844 ( .A(n14874), .B(n40650), .C(n14654), .Z(n14656) );
  HS65_LH_AOI21X2 U14845 ( .A(n15468), .B(n18029), .C(n15467), .Z(n15469) );
  HS65_LH_AOI21X2 U14846 ( .A(n14481), .B(n40472), .C(n14875), .Z(n14300) );
  HS65_LH_AOI21X2 U14847 ( .A(n15465), .B(n18034), .C(n15464), .Z(n15466) );
  HS65_LH_AOI21X2 U14848 ( .A(n14838), .B(n17594), .C(n14748), .Z(n14750) );
  HS65_LH_AOI21X2 U14849 ( .A(n17481), .B(n18039), .C(n15461), .Z(n15463) );
  HS65_LH_AOI21X2 U14850 ( .A(n14905), .B(n17595), .C(n14839), .Z(n14485) );
  HS65_LH_AOI21X2 U14851 ( .A(n15459), .B(n3798), .C(n15458), .Z(n15460) );
  HS65_LH_AOI21X2 U14852 ( .A(n14987), .B(n17596), .C(n14906), .Z(n14697) );
  HS65_LH_AOI21X2 U14853 ( .A(n15456), .B(n3695), .C(n15455), .Z(n15457) );
  HS65_LH_AOI21X2 U14854 ( .A(n15122), .B(n17597), .C(n14988), .Z(n14381) );
  HS65_LH_AOI21X2 U14855 ( .A(n15453), .B(n3592), .C(n15452), .Z(n15454) );
  HS65_LH_NAND2X2 U14856 ( .A(n14283), .B(n14910), .Z(n15248) );
  HS65_LH_AOI21X2 U14857 ( .A(n17466), .B(n17598), .C(n17465), .Z(n15054) );
  HS65_LH_AOI21X2 U14858 ( .A(n15450), .B(n3489), .C(n15449), .Z(n15451) );
  HS65_LH_AOI21X2 U14859 ( .A(n14329), .B(n6311), .C(n15015), .Z(n14330) );
  HS65_LH_AOI21X2 U14860 ( .A(n15447), .B(n3386), .C(n15446), .Z(n15448) );
  HS65_LH_AOI21X2 U14861 ( .A(n14606), .B(n14605), .C(n14604), .Z(n14607) );
  HS65_LH_AOI21X2 U14862 ( .A(n15444), .B(n3283), .C(n15443), .Z(n15445) );
  HS65_LH_IVX2 U14863 ( .A(n15062), .Z(n15324) );
  HS65_LH_IVX2 U14864 ( .A(n14852), .Z(n14850) );
  HS65_LH_AOI21X2 U14865 ( .A(n15441), .B(n3180), .C(n15440), .Z(n15442) );
  HS65_LH_IVX2 U14866 ( .A(n17254), .Z(n14583) );
  HS65_LH_IVX2 U14867 ( .A(n17989), .Z(n14035) );
  HS65_LH_AOI21X2 U14868 ( .A(n15438), .B(n3077), .C(n15437), .Z(n15439) );
  HS65_LH_OAI212X3 U14869 ( .A(n17650), .B(n17585), .C(n17622), .D(n17648), 
        .E(n15489), .Z(n15490) );
  HS65_LH_AOI21X2 U14870 ( .A(n15435), .B(n2974), .C(n15434), .Z(n15436) );
  HS65_LH_NAND2X2 U14871 ( .A(n17629), .B(n15476), .Z(n15707) );
  HS65_LH_CNIVX3 U14872 ( .A(n10911), .Z(n14050) );
  HS65_LH_CNIVX3 U14873 ( .A(\u_DataPath/dataOut_exe_i [12]), .Z(n15660) );
  HS65_LH_CNIVX3 U14874 ( .A(\u_DataPath/dataOut_exe_i [13]), .Z(n15644) );
  HS65_LH_CNIVX3 U14875 ( .A(\u_DataPath/dataOut_exe_i [15]), .Z(n14328) );
  HS65_LH_CNIVX3 U14876 ( .A(\u_DataPath/dataOut_exe_i [16]), .Z(n14990) );
  HS65_LH_CNIVX3 U14877 ( .A(\u_DataPath/dataOut_exe_i [17]), .Z(n15017) );
  HS65_LH_CNIVX3 U14878 ( .A(\u_DataPath/dataOut_exe_i [18]), .Z(n15094) );
  HS65_LH_CNIVX3 U14879 ( .A(\u_DataPath/dataOut_exe_i [19]), .Z(n14379) );
  HS65_LH_CNIVX3 U14880 ( .A(\u_DataPath/dataOut_exe_i [21]), .Z(n14695) );
  HS65_LH_CNIVX3 U14881 ( .A(\u_DataPath/dataOut_exe_i [22]), .Z(n14877) );
  HS65_LH_IVX2 U14883 ( .A(\u_DataPath/dataOut_exe_i [24]), .Z(n14802) );
  HS65_LH_IVX2 U14884 ( .A(n33776), .Z(n14452) );
  HS65_LH_IVX2 U14885 ( .A(n33771), .Z(n14213) );
  HS65_LH_IVX2 U14887 ( .A(n33654), .Z(n14653) );
  HS65_LH_CNIVX3 U14889 ( .A(addr_to_iram_5), .Z(n14082) );
  HS65_LH_CNIVX3 U14890 ( .A(addr_to_iram_7), .Z(n14084) );
  HS65_LH_CNIVX3 U14891 ( .A(addr_to_iram_9), .Z(n14086) );
  HS65_LH_CNIVX3 U14892 ( .A(addr_to_iram_11), .Z(n14088) );
  HS65_LH_CNIVX3 U14893 ( .A(addr_to_iram_13), .Z(n14090) );
  HS65_LH_CNIVX3 U14894 ( .A(addr_to_iram_15), .Z(n14092) );
  HS65_LH_BFX4 U14895 ( .A(n11877), .Z(n14051) );
  HS65_LH_CNIVX3 U14896 ( .A(\u_DataPath/dataOut_exe_i [3]), .Z(n14405) );
  HS65_LH_CNIVX3 U14897 ( .A(\u_DataPath/dataOut_exe_i [4]), .Z(n15658) );
  HS65_LH_CNIVX3 U14898 ( .A(\u_DataPath/dataOut_exe_i [5]), .Z(n15650) );
  HS65_LH_CNIVX3 U14899 ( .A(\u_DataPath/dataOut_exe_i [9]), .Z(n15656) );
  HS65_LH_CNIVX3 U14900 ( .A(\u_DataPath/dataOut_exe_i [10]), .Z(n15662) );
  HS65_LH_CNIVX3 U14901 ( .A(\u_DataPath/dataOut_exe_i [7]), .Z(n15648) );
  HS65_LH_CNIVX3 U14902 ( .A(\u_DataPath/dataOut_exe_i [11]), .Z(n15654) );
  HS65_LH_CNIVX3 U14903 ( .A(\u_DataPath/dataOut_exe_i [2]), .Z(n15699) );
  HS65_LH_OAI212X3 U14904 ( .A(n17464), .B(n17309), .C(n17588), .D(n17274), 
        .E(n17280), .Z(n15577) );
  HS65_LH_AOI21X2 U14905 ( .A(n14900), .B(n14426), .C(n14402), .Z(n15558) );
  HS65_LH_IVX2 U14906 ( .A(n14709), .Z(n15268) );
  HS65_LH_IVX2 U14907 ( .A(n15032), .Z(n15018) );
  HS65_LH_IVX2 U14908 ( .A(n15507), .Z(n15246) );
  HS65_LH_IVX2 U14909 ( .A(n32851), .Z(n14032) );
  HS65_LH_NOR3X1 U14910 ( .A(n10482), .B(n10483), .C(n11636), .Z(n15478) );
  HS65_LH_CNIVX3 U14911 ( .A(n12324), .Z(n14053) );
  HS65_LH_BFX4 U14912 ( .A(n10320), .Z(n14044) );
  HS65_LH_CNIVX3 U14913 ( .A(addr_to_iram_3), .Z(n14079) );
  HS65_LH_NOR3X1 U14914 ( .A(n15577), .B(n17317), .C(n15575), .Z(n15578) );
  HS65_LH_AOI211X1 U14915 ( .A(n15042), .B(n15381), .C(n15014), .D(n15013), 
        .Z(n15557) );
  HS65_LH_AOI21X2 U14916 ( .A(n14930), .B(n15421), .C(n14355), .Z(n15552) );
  HS65_LH_OAI222X2 U14917 ( .A(n37585), .B(n17618), .C(n14273), .D(n17344), 
        .E(n17616), .F(n17264), .Z(n14255) );
  HS65_LH_OAI222X2 U14918 ( .A(n36008), .B(n17618), .C(n14273), .D(n32281), 
        .E(n17616), .F(n33749), .Z(n14254) );
  HS65_LH_OAI222X2 U14919 ( .A(n35907), .B(n17617), .C(n14273), .D(n32258), 
        .E(n17615), .F(\u_DataPath/dataOut_exe_i [24]), .Z(n14253) );
  HS65_LH_OAI222X2 U14920 ( .A(n37932), .B(n17618), .C(n14273), .D(n17867), 
        .E(n17615), .F(n17859), .Z(n14215) );
  HS65_LH_OAI212X3 U14921 ( .A(n17518), .B(n17704), .C(n17619), .D(n34391), 
        .E(n17844), .Z(n15177) );
  HS65_LH_AOI212X2 U14922 ( .A(n17506), .B(n17728), .C(n17709), .D(n17508), 
        .E(n15178), .Z(n15182) );
  HS65_LH_AOI212X2 U14923 ( .A(n14042), .B(\u_DataPath/rs_ex_i [3]), .C(
        \u_DataPath/u_idexreg/N56 ), .D(n14050), .E(n14135), .Z(n14138) );
  HS65_LH_AOI212X2 U14924 ( .A(n14041), .B(\u_DataPath/rs_ex_i [2]), .C(
        \u_DataPath/rs_ex_i [1]), .D(n14040), .E(n14136), .Z(n14137) );
  HS65_LH_CNIVX3 U14925 ( .A(\u_DataPath/dataOut_exe_i [6]), .Z(n15652) );
  HS65_LH_CNIVX3 U14926 ( .A(n10592), .Z(n14067) );
  HS65_LH_CNIVX3 U14927 ( .A(n9568), .Z(n14039) );
  HS65_LH_IVX2 U14929 ( .A(n14521), .Z(n14031) );
  HS65_LH_IVX2 U14930 ( .A(n18016), .Z(n14029) );
  HS65_LH_OAI222X2 U14931 ( .A(n37340), .B(n17617), .C(n14273), .D(n32236), 
        .E(n17615), .F(\u_DataPath/dataOut_exe_i [25]), .Z(n14252) );
  HS65_LH_AOI212X2 U14933 ( .A(n17480), .B(n17707), .C(n17628), .D(n17702), 
        .E(n15180), .Z(n15181) );
  HS65_LH_CNIVX3 U14934 ( .A(n12490), .Z(n258) );
  HS65_LH_IVX2 U14935 ( .A(\u_DataPath/dataOut_exe_i [31]), .Z(n15387) );
  HS65_LH_NAND3AX3 U14936 ( .A(n35243), .B(n39446), .C(n39444), .Z(n15491) );
  HS65_LH_IVX2 U14937 ( .A(n17249), .Z(n14036) );
  HS65_LH_IVX2 U14938 ( .A(n15337), .Z(n15163) );
  HS65_LH_CBI4I1X3 U14940 ( .A(n15186), .B(n10704), .C(n15185), .D(n15703), 
        .Z(n288) );
  HS65_LH_CNIVX3 U14941 ( .A(n8860), .Z(n14110) );
  HS65_LH_CBI4I6X2 U14942 ( .A(n17463), .B(n17462), .C(n17308), .D(n15425), 
        .Z(n15572) );
  HS65_LH_OAI21X2 U14943 ( .A(n14694), .B(n14693), .C(n14692), .Z(n15576) );
  HS65_LH_OAI21X2 U14944 ( .A(n15217), .B(n15051), .C(n15050), .Z(n15559) );
  HS65_LH_OAI211X1 U14945 ( .A(n14474), .B(n15080), .C(n14435), .D(n14434), 
        .Z(n14436) );
  HS65_LH_OA12X4 U14946 ( .A(n15464), .B(n18118), .C(n15468), .Z(n14103) );
  HS65_LH_OA12X4 U14947 ( .A(n15461), .B(n18116), .C(n15465), .Z(n14101) );
  HS65_LH_AOI21X2 U14948 ( .A(n17314), .B(n14788), .C(n14787), .Z(n14789) );
  HS65_LH_OA12X4 U14949 ( .A(n17482), .B(n18114), .C(n17481), .Z(n14099) );
  HS65_LH_OA12X4 U14951 ( .A(n15455), .B(addr_to_iram_20), .C(n15459), .Z(
        n14097) );
  HS65_LH_OA12X4 U14952 ( .A(n15452), .B(addr_to_iram_18), .C(n15456), .Z(
        n14095) );
  HS65_LH_OAI211X1 U14953 ( .A(n33045), .B(n14358), .C(n17314), .D(n14279), 
        .Z(n14359) );
  HS65_LH_MX41X4 U14954 ( .D0(n17433), .S0(n17573), .D1(n17206), .S1(n17576), 
        .D2(n17514), .S2(n17305), .D3(n17444), .S3(n17302), .Z(n197) );
  HS65_LH_OAI222X2 U14955 ( .A(n38185), .B(n17617), .C(n14273), .D(n32214), 
        .E(n17615), .F(n33776), .Z(n14251) );
  HS65_LH_OAI222X2 U14956 ( .A(n37666), .B(n17618), .C(n14273), .D(n17337), 
        .E(n17616), .F(n17372), .Z(n14258) );
  HS65_LH_BFX4 U14957 ( .A(n14210), .Z(n14034) );
  HS65_LH_NOR2X2 U14958 ( .A(n13646), .B(n13879), .Z(n15748) );
  HS65_LH_NAND2X2 U14959 ( .A(n13887), .B(n15429), .Z(n236) );
  HS65_LH_AOI212X2 U14960 ( .A(n14652), .B(n14651), .C(n15187), .D(n14650), 
        .E(n14649), .Z(n15551) );
  HS65_LH_OAI21X2 U14961 ( .A(n33693), .B(n33687), .C(n14960), .Z(n15549) );
  HS65_LH_CBI4I6X2 U14962 ( .A(n15206), .B(n14603), .C(n14602), .D(n14601), 
        .Z(n15546) );
  HS65_LH_NOR4ABX2 U14963 ( .A(n14249), .B(n15098), .C(n14248), .D(n14247), 
        .Z(n14250) );
  HS65_LH_NOR4ABX2 U14964 ( .A(n14499), .B(n14498), .C(n14497), .D(n14496), 
        .Z(n14500) );
  HS65_LH_IVX2 U14966 ( .A(n17260), .Z(n14030) );
  HS65_LH_OAI222X2 U14967 ( .A(n17611), .B(n17940), .C(n17631), .D(n33654), 
        .E(n17610), .F(n17361), .Z(n14521) );
  HS65_LH_OAI222X2 U14968 ( .A(n14141), .B(n8318), .C(n14239), .D(
        \u_DataPath/dataOut_exe_i [8]), .E(n14238), .F(n4737), .Z(n15240) );
  HS65_LH_AOI21X2 U14969 ( .A(n17514), .B(n17566), .C(n17296), .Z(n195) );
  HS65_LH_OAI222X2 U14970 ( .A(n38105), .B(n17617), .C(n17614), .D(n17334), 
        .E(n17615), .F(n17263), .Z(n14259) );
  HS65_LH_OAI222X2 U14971 ( .A(n36776), .B(n17617), .C(n17614), .D(n17351), 
        .E(n17615), .F(n17292), .Z(n14266) );
  HS65_LH_OAI222X2 U14972 ( .A(n36435), .B(n17617), .C(n17614), .D(n17352), 
        .E(n17615), .F(n17367), .Z(n14264) );
  HS65_LH_OAI222X2 U14973 ( .A(n36720), .B(n17617), .C(n14273), .D(n17350), 
        .E(n17615), .F(n17290), .Z(n14268) );
  HS65_LH_OAI222X2 U14974 ( .A(n38385), .B(n17617), .C(n14273), .D(n17354), 
        .E(n17615), .F(n17287), .Z(n14222) );
  HS65_LH_OAI222X2 U14975 ( .A(n36130), .B(n17617), .C(n17614), .D(n17345), 
        .E(n17615), .F(n17364), .Z(n14270) );
  HS65_LH_OAI222X2 U14976 ( .A(n36661), .B(n17617), .C(n14273), .D(n17348), 
        .E(n17615), .F(n17366), .Z(n14269) );
  HS65_LH_OAI222X2 U14977 ( .A(n37261), .B(n17617), .C(n17614), .D(n17330), 
        .E(n17615), .F(n17370), .Z(n14262) );
  HS65_LH_NOR2X2 U14978 ( .A(n13890), .B(n236), .Z(n274) );
  HS65_LH_AOI211X1 U14979 ( .A(n17648), .B(n17508), .C(n15174), .D(n15173), 
        .Z(n15175) );
  HS65_LH_OA12X4 U14980 ( .A(n15446), .B(addr_to_iram_14), .C(n15450), .Z(
        n14091) );
  HS65_LH_NOR2X2 U14981 ( .A(n11644), .B(n1101), .Z(n196) );
  HS65_LH_OA12X4 U14982 ( .A(n15443), .B(addr_to_iram_12), .C(n15447), .Z(
        n14089) );
  HS65_LH_CNIVX3 U14983 ( .A(n9652), .Z(n14040) );
  HS65_LH_CNIVX3 U14984 ( .A(n9803), .Z(n14042) );
  HS65_LH_CNIVX3 U14985 ( .A(n10156), .Z(n14106) );
  HS65_LH_CNIVX3 U14986 ( .A(\u_DataPath/pc_4_to_ex_i [13]), .Z(n14605) );
  HS65_LH_OAI211X1 U14987 ( .A(n33880), .B(n15505), .C(n15504), .D(n15503), 
        .Z(n15534) );
  HS65_LH_NOR2X9 U14988 ( .A(n15700), .B(n15660), .Z(n15661) );
  HS65_LH_NOR2X9 U14989 ( .A(n15700), .B(n15656), .Z(n15657) );
  HS65_LH_NOR2X9 U14990 ( .A(n15700), .B(n15644), .Z(n15645) );
  HS65_LH_NOR2X9 U14991 ( .A(n15700), .B(n15654), .Z(n15655) );
  HS65_LH_AOI222X2 U14992 ( .A(n8226), .B(n15209), .C(n15208), .D(
        \u_DataPath/data_read_ex_2_i [4]), .E(n15207), .F(
        \u_DataPath/dataOut_exe_i [4]), .Z(n14224) );
  HS65_LH_AOI222X2 U14993 ( .A(n9252), .B(n15209), .C(n15208), .D(n9202), .E(
        n15207), .F(n10704), .Z(n14217) );
  HS65_LH_AOI222X2 U14994 ( .A(n17311), .B(n17479), .C(n17478), .D(n17342), 
        .E(n17312), .F(\u_DataPath/dataOut_exe_i [31]), .Z(n15211) );
  HS65_LH_NOR2X9 U14995 ( .A(n15700), .B(n15652), .Z(n15653) );
  HS65_LH_NOR2X9 U14996 ( .A(n15700), .B(n15646), .Z(n15647) );
  HS65_LH_AOI222X2 U14997 ( .A(n6572), .B(n15209), .C(n15208), .D(
        \u_DataPath/data_read_ex_2_i [3]), .E(n15207), .F(
        \u_DataPath/dataOut_exe_i [3]), .Z(n14220) );
  HS65_LH_NOR2X9 U14998 ( .A(n15700), .B(n15658), .Z(n15659) );
  HS65_LH_NOR2X9 U14999 ( .A(n15700), .B(n15648), .Z(n15649) );
  HS65_LH_NOR3X1 U15000 ( .A(n12482), .B(n15643), .C(n15742), .Z(n178) );
  HS65_LH_CNIVX3 U15001 ( .A(n15474), .Z(n15475) );
  HS65_LH_CNIVX3 U15002 ( .A(n10158), .Z(n15477) );
  HS65_LL_OAI12X12 U15003 ( .A(n17306), .B(n101), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N136 ) );
  HS65_LL_OR2ABX27 U15005 ( .A(n15696), .B(n15694), .Z(write_op_snps_wire) );
  HS65_LH_NAND2X2 U15006 ( .A(n13578), .B(n12382), .Z(n16497) );
  HS65_LH_CNIVX3 U15007 ( .A(n9722), .Z(n14041) );
  HS65_LH_NAND2X2 U15008 ( .A(n9296), .B(n14076), .Z(n15702) );
  HS65_LH_IVX7 U15009 ( .A(n14065), .Z(n15696) );
  HS65_LL_OAI12X12 U15010 ( .A(n99), .B(n17306), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N128 ) );
  HS65_LL_OAI12X12 U15011 ( .A(n17306), .B(n104), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N144 ) );
  HS65_LL_OAI12X12 U15012 ( .A(n17306), .B(n113), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N152 ) );
  HS65_LH_NOR3X4 U15013 ( .A(n14291), .B(n15385), .C(n14244), .Z(n15151) );
  HS65_LH_NOR2X5 U15014 ( .A(\u_DataPath/cw_towb_i [1]), .B(
        \u_DataPath/regfile_addr_out_towb_i [1]), .Z(n15714) );
  HS65_LH_NOR3X7 U15015 ( .A(\u_DataPath/cw_to_ex_i [2]), .B(
        \u_DataPath/cw_to_ex_i [1]), .C(n15385), .Z(n15501) );
  HS65_LH_OR2X4 U15016 ( .A(\u_DataPath/cw_towb_i [1]), .B(
        \u_DataPath/regfile_addr_out_towb_i [4]), .Z(n14124) );
  HS65_LH_NOR2X5 U15017 ( .A(\u_DataPath/regfile_addr_out_towb_i [0]), .B(
        \u_DataPath/cw_towb_i [1]), .Z(n15711) );
  HS65_LH_MUXI21X2 U15018 ( .D0(n14039), .D1(n9568), .S0(
        \u_DataPath/rs_ex_i [0]), .Z(n14140) );
  HS65_LH_BFX4 U15019 ( .A(addr_to_iram_4), .Z(n14059) );
  HS65_LH_NAND2X2 U15020 ( .A(n11878), .B(n12291), .Z(n15781) );
  HS65_LH_NAND2X2 U15021 ( .A(n1912), .B(n1913), .Z(n15791) );
  HS65_LH_NAND2X2 U15022 ( .A(n15331), .B(n14930), .Z(n15417) );
  HS65_LH_NOR2X6 U15023 ( .A(n15245), .B(n6651), .Z(n15331) );
  HS65_LH_CNIVX3 U15024 ( .A(n14124), .Z(n17211) );
  HS65_LH_BFX4 U15026 ( .A(n14072), .Z(n15694) );
  HS65_LH_MUXI21X2 U15027 ( .D0(n12625), .D1(n10156), .S0(n14002), .Z(n14107)
         );
  HS65_LH_NAND2X2 U15028 ( .A(n2733), .B(n35704), .Z(n2048) );
  HS65_LH_NAND2X2 U15029 ( .A(n2733), .B(n31717), .Z(n2360) );
  HS65_LH_NAND2X2 U15030 ( .A(n2733), .B(n36304), .Z(n2336) );
  HS65_LH_NAND2X2 U15031 ( .A(n2733), .B(n36483), .Z(n2432) );
  HS65_LH_NAND2X2 U15032 ( .A(n2733), .B(n35844), .Z(n2240) );
  HS65_LH_NAND2X2 U15033 ( .A(n2733), .B(n38437), .Z(n2624) );
  HS65_LH_NAND2X2 U15034 ( .A(n2733), .B(n36770), .Z(n2456) );
  HS65_LH_NAND2X2 U15035 ( .A(n2733), .B(n38185), .Z(n2072) );
  HS65_LH_NAND2X2 U15036 ( .A(n2733), .B(n36008), .Z(n2144) );
  HS65_LH_NAND2X2 U15037 ( .A(n2733), .B(n38238), .Z(n1976) );
  HS65_LH_NAND2X2 U15038 ( .A(n2733), .B(n36430), .Z(n2408) );
  HS65_LH_NAND2X2 U15039 ( .A(n2733), .B(n36658), .Z(n2528) );
  HS65_LH_NAND2X2 U15040 ( .A(n2733), .B(n36569), .Z(n2384) );
  HS65_LH_NAND2X2 U15041 ( .A(n2733), .B(n38329), .Z(n2000) );
  HS65_LH_NAND2X2 U15042 ( .A(n2733), .B(n35942), .Z(n2192) );
  HS65_LH_NAND2X2 U15043 ( .A(n2733), .B(n36130), .Z(n2576) );
  HS65_LH_NAND2X2 U15044 ( .A(n2733), .B(n37340), .Z(n2096) );
  HS65_LH_NAND2X2 U15045 ( .A(n2733), .B(n36047), .Z(n2480) );
  HS65_LH_NAND2X2 U15046 ( .A(n2733), .B(n35907), .Z(n2120) );
  HS65_LH_NAND2X2 U15047 ( .A(n2733), .B(n37503), .Z(n2024) );
  HS65_LH_NAND2X2 U15048 ( .A(n2733), .B(n36394), .Z(n2168) );
  HS65_LH_NAND2X2 U15049 ( .A(n2733), .B(n38016), .Z(n2600) );
  HS65_LH_NAND2X2 U15050 ( .A(n2733), .B(n36714), .Z(n2504) );
  HS65_LH_NAND2X2 U15051 ( .A(n2733), .B(n38100), .Z(n2216) );
  HS65_LH_NAND2X2 U15052 ( .A(n2733), .B(n35810), .Z(n2312) );
  HS65_LH_NAND2X2 U15053 ( .A(n2733), .B(n36239), .Z(n2288) );
  HS65_LH_NAND2X2 U15054 ( .A(n2733), .B(n38385), .Z(n2648) );
  HS65_LH_NAND2X2 U15055 ( .A(n2733), .B(n36864), .Z(n2264) );
  HS65_LH_NAND2X2 U15056 ( .A(n2733), .B(n35736), .Z(n2552) );
  HS65_LH_NAND2X2 U15057 ( .A(n2733), .B(n37932), .Z(n2672) );
  HS65_LH_NAND2X2 U15058 ( .A(n2733), .B(n32443), .Z(n2729) );
  HS65_LH_NOR3AX4 U15059 ( .A(n15706), .B(n10732), .C(n10704), .Z(n15750) );
  HS65_LH_NOR2X3 U15060 ( .A(n15750), .B(\nibble[0]_snps_wire ), .Z(n17197) );
  HS65_LH_NAND2X2 U15061 ( .A(n2733), .B(n40882), .Z(n1952) );
  HS65_LH_NOR2X2 U15062 ( .A(rst), .B(n17830), .Z(n74) );
  HS65_LH_AOI211X1 U15063 ( .A(n29624), .B(n14537), .C(n14536), .D(n14535), 
        .Z(n14538) );
  HS65_LH_IVX44 U15064 ( .A(n15696), .Z(write_byte_snps_wire) );
  HS65_LH_NOR2X2 U15065 ( .A(rst), .B(n33770), .Z(
        \u_DataPath/from_alu_data_out_i [27]) );
  HS65_LH_NOR2X2 U15066 ( .A(rst), .B(n31771), .Z(
        \u_DataPath/from_alu_data_out_i [14]) );
  HS65_LH_NOR2X2 U15067 ( .A(rst), .B(n32578), .Z(
        \u_DataPath/from_alu_data_out_i [15]) );
  HS65_LH_NOR2X2 U15068 ( .A(rst), .B(n32964), .Z(
        \u_DataPath/from_alu_data_out_i [11]) );
  HS65_LH_NOR2X2 U15069 ( .A(rst), .B(n33760), .Z(
        \u_DataPath/from_alu_data_out_i [19]) );
  HS65_LH_NOR2X2 U15070 ( .A(rst), .B(n33935), .Z(
        \u_DataPath/from_alu_data_out_i [3]) );
  HS65_LH_NOR2X2 U15071 ( .A(rst), .B(n33179), .Z(
        \u_DataPath/from_alu_data_out_i [10]) );
  HS65_LH_NOR2X2 U15072 ( .A(rst), .B(n33775), .Z(
        \u_DataPath/from_alu_data_out_i [26]) );
  HS65_LH_NOR2X2 U15073 ( .A(rst), .B(n33750), .Z(
        \u_DataPath/from_alu_data_out_i [23]) );
  HS65_LH_NOR2X2 U15074 ( .A(rst), .B(n21749), .Z(
        \u_DataPath/from_alu_data_out_i [30]) );
  HS65_LH_NOR2X2 U15075 ( .A(rst), .B(n32889), .Z(
        \u_DataPath/from_alu_data_out_i [12]) );
  HS65_LH_NOR2X2 U15076 ( .A(rst), .B(n33438), .Z(
        \u_DataPath/from_alu_data_out_i [7]) );
  HS65_LH_NOR2X2 U15077 ( .A(rst), .B(n32813), .Z(
        \u_DataPath/from_alu_data_out_i [13]) );
  HS65_LH_NOR2X2 U15078 ( .A(rst), .B(n14653), .Z(
        \u_DataPath/from_alu_data_out_i [29]) );
  HS65_LH_NOR2X2 U15079 ( .A(rst), .B(n33752), .Z(
        \u_DataPath/from_alu_data_out_i [21]) );
  HS65_LH_NOR2X2 U15080 ( .A(rst), .B(n33896), .Z(
        \u_DataPath/from_alu_data_out_i [5]) );
  HS65_LH_NOR2X2 U15081 ( .A(rst), .B(n33772), .Z(
        \u_DataPath/from_alu_data_out_i [25]) );
  HS65_LH_NOR2X2 U15082 ( .A(rst), .B(n33366), .Z(
        \u_DataPath/from_alu_data_out_i [9]) );
  HS65_LH_NOR2X2 U15083 ( .A(rst), .B(n33757), .Z(
        \u_DataPath/from_alu_data_out_i [24]) );
  HS65_LH_NOR2X2 U15084 ( .A(rst), .B(n33783), .Z(
        \u_DataPath/from_alu_data_out_i [28]) );
  HS65_LH_NOR2X2 U15085 ( .A(rst), .B(n33765), .Z(
        \u_DataPath/from_alu_data_out_i [22]) );
  HS65_LH_NOR2X2 U15086 ( .A(rst), .B(n33904), .Z(
        \u_DataPath/from_alu_data_out_i [4]) );
  HS65_LH_NOR2X2 U15087 ( .A(rst), .B(n33402), .Z(
        \u_DataPath/from_alu_data_out_i [8]) );
  HS65_LH_NOR2X2 U15088 ( .A(rst), .B(n33777), .Z(
        \u_DataPath/from_alu_data_out_i [20]) );
  HS65_LH_NOR2X2 U15089 ( .A(rst), .B(n33649), .Z(
        \u_DataPath/from_alu_data_out_i [16]) );
  HS65_LH_NOR2X2 U15090 ( .A(rst), .B(n33738), .Z(
        \u_DataPath/from_alu_data_out_i [17]) );
  HS65_LH_NOR2X2 U15091 ( .A(rst), .B(n31972), .Z(
        \u_DataPath/mem_writedata_out_i [2]) );
  HS65_LH_NOR2X2 U15092 ( .A(rst), .B(n33950), .Z(
        \u_DataPath/from_alu_data_out_i [2]) );
  HS65_LH_NOR2X2 U15093 ( .A(rst), .B(n33743), .Z(
        \u_DataPath/from_alu_data_out_i [18]) );
  HS65_LH_NOR2X2 U15094 ( .A(rst), .B(n33824), .Z(
        \u_DataPath/from_alu_data_out_i [6]) );
  HS65_LH_NOR2X2 U15095 ( .A(rst), .B(n34063), .Z(
        \u_DataPath/from_alu_data_out_i [31]) );
  HS65_LH_NOR2X2 U15096 ( .A(rst), .B(n29744), .Z(\u_DataPath/u_idexreg/N25 )
         );
  HS65_LH_NOR2X2 U15097 ( .A(rst), .B(n38604), .Z(\u_DataPath/u_idexreg/N26 )
         );
  HS65_LH_NOR2X2 U15098 ( .A(rst), .B(n40524), .Z(\u_DataPath/u_idexreg/N27 )
         );
  HS65_LH_NOR2X2 U15099 ( .A(rst), .B(n29765), .Z(\u_DataPath/u_idexreg/N28 )
         );
  HS65_LH_NOR2X2 U15100 ( .A(rst), .B(n38583), .Z(\u_DataPath/u_idexreg/N30 )
         );
  HS65_LH_NOR2X2 U15101 ( .A(rst), .B(n38670), .Z(\u_DataPath/u_idexreg/N42 )
         );
  HS65_LH_NOR2X2 U15102 ( .A(rst), .B(n38626), .Z(\u_DataPath/idex_rt_i [2])
         );
  HS65_LH_NOR2X2 U15103 ( .A(rst), .B(n29705), .Z(\u_DataPath/u_idexreg/N44 )
         );
  HS65_LH_NOR2X2 U15104 ( .A(rst), .B(n39628), .Z(\u_DataPath/idex_rt_i [4])
         );
  HS65_LH_NOR2X2 U15105 ( .A(rst), .B(n40163), .Z(\u_DataPath/rs_ex_i [0]) );
  HS65_LH_NOR2X2 U15106 ( .A(rst), .B(n29767), .Z(\u_DataPath/rs_ex_i [1]) );
  HS65_LH_NOR2X2 U15107 ( .A(rst), .B(n40228), .Z(\u_DataPath/rs_ex_i [2]) );
  HS65_LH_NOR2X2 U15108 ( .A(rst), .B(n19087), .Z(\u_DataPath/rs_ex_i [3]) );
  HS65_LH_NOR2X2 U15109 ( .A(rst), .B(n34425), .Z(\u_DataPath/cw_tomem_i [3])
         );
  HS65_LH_NOR2X2 U15110 ( .A(rst), .B(n39629), .Z(\u_DataPath/idex_rt_i [0])
         );
  HS65_LH_NAND2X2 U15111 ( .A(n10710), .B(n14067), .Z(n14064) );
  HS65_LH_CNIVX3 U15115 ( .A(n11868), .Z(n1912) );
  HS65_LH_CNIVX3 U15116 ( .A(n12281), .Z(n1913) );
  HS65_LH_NOR4ABX4 U15117 ( .A(n10603), .B(n10721), .C(n10596), .D(n10678), 
        .Z(n14065) );
  HS65_LH_NOR2X2 U15118 ( .A(n10575), .B(n10573), .Z(n14076) );
  HS65_LH_NAND2X2 U15119 ( .A(n10721), .B(n14067), .Z(n14074) );
  HS65_LH_OA12X4 U15120 ( .A(n14067), .B(n10721), .C(n14074), .Z(n14068) );
  HS65_LH_CNIVX3 U15121 ( .A(n10704), .Z(n14070) );
  HS65_LH_NOR4ABX2 U15122 ( .A(n10575), .B(n10721), .C(n10573), .D(n10678), 
        .Z(n14077) );
  HS65_LL_AND2X18 U15123 ( .A(\u_DataPath/mem_writedata_out_i [0]), .B(
        write_op_snps_wire), .Z(Data_in_0) );
  HS65_LH_NOR4ABX2 U15124 ( .A(n10589), .B(n10721), .C(n10592), .D(n10585), 
        .Z(n14073) );
  HS65_LH_NAND3X2 U15125 ( .A(n15702), .B(n15696), .C(n9305), .Z(n15706) );
  HS65_LH_NAND2X2 U15126 ( .A(n14076), .B(n10676), .Z(n15704) );
  HS65_LH_NAND2AX4 U15127 ( .A(n14077), .B(n10565), .Z(n15185) );
  HS65_LL_AND2ABX18 U15128 ( .A(n14078), .B(n14877), .Z(Address_toRAM_20) );
  HS65_LL_AND2ABX18 U15129 ( .A(n17524), .B(n14802), .Z(Address_toRAM[22]) );
  HS65_LL_AND2ABX18 U15130 ( .A(n17524), .B(n26577), .Z(Address_toRAM[21]) );
  HS65_LL_AND2ABX18 U15131 ( .A(n17524), .B(n14747), .Z(Address_toRAM[23]) );
  HS65_LL_AND2ABX18 U15132 ( .A(n14078), .B(n14695), .Z(Address_toRAM_19) );
  HS65_LL_AND2ABX18 U15133 ( .A(n17524), .B(n14213), .Z(Address_toRAM[25]) );
  HS65_LL_AND2ABX18 U15134 ( .A(n17524), .B(n21749), .Z(Address_toRAM[28]) );
  HS65_LL_AND2ABX18 U15135 ( .A(n14078), .B(n14328), .Z(Address_toRAM_13) );
  HS65_LL_AND2ABX18 U15136 ( .A(n14078), .B(n15017), .Z(Address_toRAM_15) );
  HS65_LL_AND2ABX18 U15137 ( .A(n17524), .B(n26759), .Z(Address_toRAM[26]) );
  HS65_LL_AND2ABX18 U15138 ( .A(n17524), .B(n15387), .Z(Address_toRAM[29]) );
  HS65_LL_AND2ABX18 U15139 ( .A(n14078), .B(n15094), .Z(Address_toRAM_16) );
  HS65_LL_AND2ABX18 U15140 ( .A(n17524), .B(n14452), .Z(Address_toRAM[24]) );
  HS65_LL_AND2ABX18 U15141 ( .A(n14078), .B(n14990), .Z(Address_toRAM_14) );
  HS65_LL_AND2ABX18 U15142 ( .A(n14078), .B(n14379), .Z(Address_toRAM_17) );
  HS65_LL_AND2ABX18 U15143 ( .A(n17524), .B(n14653), .Z(Address_toRAM[27]) );
  HS65_LH_BFX4 U15144 ( .A(n14078), .Z(n15700) );
  HS65_LL_AND2ABX18 U15145 ( .A(n15700), .B(n14405), .Z(Address_toRAM_1) );
  HS65_LH_NAND3X2 U15146 ( .A(n14006), .B(n14004), .C(addr_to_iram_2), .Z(
        n15432) );
  HS65_LH_NOR2X2 U15147 ( .A(n14079), .B(n15432), .Z(n15431) );
  HS65_LH_NAND2X2 U15148 ( .A(n15431), .B(n14059), .Z(n15435) );
  HS65_LH_CB4I1X4 U15149 ( .A(n14004), .B(n12637), .C(addr_to_iram_2), .D(
        n15432), .Z(n14081) );
  HS65_LH_NOR2X2 U15150 ( .A(n14082), .B(n15435), .Z(n15434) );
  HS65_LH_NAND2X2 U15151 ( .A(n15434), .B(addr_to_iram_6), .Z(n15438) );
  HS65_LH_NOR2X2 U15152 ( .A(n14084), .B(n15438), .Z(n15437) );
  HS65_LH_NAND2X2 U15153 ( .A(n15437), .B(addr_to_iram_8), .Z(n15441) );
  HS65_LH_NOR2X2 U15154 ( .A(n14086), .B(n15441), .Z(n15440) );
  HS65_LH_NAND2X2 U15155 ( .A(n15440), .B(addr_to_iram_10), .Z(n15444) );
  HS65_LH_NOR2X2 U15156 ( .A(n14088), .B(n15444), .Z(n15443) );
  HS65_LH_NAND2X2 U15157 ( .A(n15443), .B(addr_to_iram_12), .Z(n15447) );
  HS65_LH_NOR2X2 U15158 ( .A(n14090), .B(n15447), .Z(n15446) );
  HS65_LH_NAND2X2 U15159 ( .A(n15446), .B(addr_to_iram_14), .Z(n15450) );
  HS65_LH_NOR2X2 U15160 ( .A(n14092), .B(n15450), .Z(n15449) );
  HS65_LH_NAND2X2 U15161 ( .A(n15449), .B(addr_to_iram_16), .Z(n15453) );
  HS65_LH_NOR2X2 U15162 ( .A(n14094), .B(n15453), .Z(n15452) );
  HS65_LH_NAND2X2 U15163 ( .A(n15452), .B(addr_to_iram_18), .Z(n15456) );
  HS65_LH_NOR2X2 U15164 ( .A(n14096), .B(n15456), .Z(n15455) );
  HS65_LH_NAND2X2 U15165 ( .A(n15455), .B(addr_to_iram_20), .Z(n15459) );
  HS65_LH_NOR2X2 U15166 ( .A(n14098), .B(n15459), .Z(n15458) );
  HS65_LH_NAND2X2 U15167 ( .A(n15458), .B(addr_to_iram_22), .Z(n15462) );
  HS65_LH_NOR2X2 U15168 ( .A(n17637), .B(n17481), .Z(n15461) );
  HS65_LH_NAND2X2 U15169 ( .A(n15461), .B(n18116), .Z(n15465) );
  HS65_LH_NAND2X2 U15171 ( .A(n15464), .B(n18118), .Z(n15468) );
  HS65_LH_NOR2X2 U15172 ( .A(n17635), .B(n15468), .Z(n15467) );
  HS65_LH_NAND2X2 U15173 ( .A(n15467), .B(n18119), .Z(n14108) );
  HS65_LH_OA12X4 U15174 ( .A(n15467), .B(n18119), .C(n14108), .Z(n14105) );
  HS65_LH_CNIVX3 U15175 ( .A(n9374), .Z(n14111) );
  HS65_LH_CNIVX3 U15176 ( .A(\u_DataPath/u_idexreg/N25 ), .Z(n15165) );
  HS65_LH_NOR2X2 U15177 ( .A(n14111), .B(n15165), .Z(n15164) );
  HS65_LH_MUX21X4 U15178 ( .D0(\u_DataPath/from_alu_data_out_i [18]), .D1(
        \u_DataPath/from_mem_data_out_i [18]), .S0(\u_DataPath/cw_towb_i [0]), 
        .Z(n14113) );
  HS65_LH_NAND4ABX3 U15179 ( .A(n9722), .B(n9652), .C(n14050), .D(n14039), .Z(
        n14114) );
  HS65_LH_OAI21X2 U15180 ( .A(n9803), .B(n14114), .C(n9996), .Z(n14139) );
  HS65_LH_CNIVX3 U15181 ( .A(\u_DataPath/idex_rt_i [0]), .Z(n14115) );
  HS65_LH_AOI22X1 U15182 ( .A(n14039), .B(n9597), .C(n14042), .D(n9832), .Z(
        n14116) );
  HS65_LH_OAI212X3 U15183 ( .A(n14039), .B(n9593), .C(n14042), .D(n9832), .E(
        n14116), .Z(n14122) );
  HS65_LH_CNIVX3 U15184 ( .A(n9744), .Z(n15485) );
  HS65_LH_CNIVX3 U15185 ( .A(n13537), .Z(n14117) );
  HS65_LH_CNIVX3 U15186 ( .A(\u_DataPath/idex_rt_i [4]), .Z(n14118) );
  HS65_LH_OAI22X1 U15187 ( .A(n14040), .B(n9682), .C(n14050), .D(n9890), .Z(
        n14119) );
  HS65_LH_AOI212X2 U15188 ( .A(n14040), .B(n9678), .C(n9884), .D(n14050), .E(
        n14119), .Z(n14120) );
  HS65_LH_OAI212X3 U15189 ( .A(n9722), .B(n15485), .C(n14041), .D(n9748), .E(
        n14120), .Z(n14121) );
  HS65_LH_NOR3X1 U15190 ( .A(n14139), .B(n14122), .C(n14121), .Z(n15207) );
  HS65_LH_CNIVX3 U15191 ( .A(n9834), .Z(n15488) );
  HS65_LH_CNIVX3 U15192 ( .A(n1907), .Z(n1106) );
  HS65_LH_CNIVX3 U15193 ( .A(\u_DataPath/regfile_addr_out_towb_i [2]), .Z(
        n15713) );
  HS65_LH_OAI31X1 U15194 ( .A(\u_DataPath/regfile_addr_out_towb_i [4]), .B(
        n105), .C(n1106), .D(n9538), .Z(n102) );
  HS65_LH_NOR2X2 U15195 ( .A(\u_DataPath/regfile_addr_out_towb_i [2]), .B(
        \u_DataPath/cw_towb_i [1]), .Z(n15670) );
  HS65_LH_AOI22X1 U15196 ( .A(n9587), .B(n15711), .C(n9754), .D(n15670), .Z(
        n14123) );
  HS65_LH_OAI212X3 U15197 ( .A(n9589), .B(n15711), .C(n9752), .D(n15670), .E(
        n14123), .Z(n14127) );
  HS65_LH_AOI22X1 U15198 ( .A(n9892), .B(n17211), .C(n9682), .D(n15714), .Z(
        n14125) );
  HS65_LH_OAI212X3 U15199 ( .A(n9890), .B(n17211), .C(n9682), .D(n15714), .E(
        n14125), .Z(n14126) );
  HS65_LH_NOR3X1 U15200 ( .A(n102), .B(n14127), .C(n14126), .Z(n14128) );
  HS65_LH_OAI212X3 U15201 ( .A(n9832), .B(n1907), .C(n15488), .D(n1106), .E(
        n14128), .Z(n14129) );
  HS65_LH_NOR2X2 U15202 ( .A(n15207), .B(n14129), .Z(n15209) );
  HS65_LH_CNIVX3 U15203 ( .A(n15209), .Z(n14257) );
  HS65_LH_BFX4 U15204 ( .A(n14257), .Z(n14274) );
  HS65_LH_CNIVX3 U15205 ( .A(n15207), .Z(n14256) );
  HS65_LH_BFX4 U15206 ( .A(n14256), .Z(n14272) );
  HS65_LH_AND2X4 U15207 ( .A(n14272), .B(n14129), .Z(n15208) );
  HS65_LH_CNIVX3 U15208 ( .A(n15208), .Z(n14206) );
  HS65_LH_OAI222X2 U15209 ( .A(n37125), .B(n17617), .C(n17614), .D(n17343), 
        .E(n17615), .F(n17262), .Z(n14276) );
  HS65_LH_AOI22X1 U15210 ( .A(n17211), .B(\u_DataPath/u_idexreg/N56 ), .C(
        n15711), .D(\u_DataPath/rs_ex_i [0]), .Z(n14130) );
  HS65_LH_OAI212X3 U15211 ( .A(n17211), .B(\u_DataPath/u_idexreg/N56 ), .C(
        n15711), .D(\u_DataPath/rs_ex_i [0]), .E(n14130), .Z(n14134) );
  HS65_LH_CNIVX3 U15212 ( .A(n15670), .Z(n15669) );
  HS65_LH_MUXI21X2 U15213 ( .D0(n15669), .D1(n15670), .S0(
        \u_DataPath/rs_ex_i [2]), .Z(n14133) );
  HS65_LH_OAI22X1 U15214 ( .A(n15714), .B(\u_DataPath/rs_ex_i [1]), .C(
        \u_DataPath/rs_ex_i [3]), .D(n1907), .Z(n14131) );
  HS65_LH_AOI212X2 U15215 ( .A(n15714), .B(\u_DataPath/rs_ex_i [1]), .C(n1907), 
        .D(\u_DataPath/rs_ex_i [3]), .E(n14131), .Z(n14132) );
  HS65_LH_NAND4ABX3 U15216 ( .A(n102), .B(n14134), .C(n14133), .D(n14132), .Z(
        n14142) );
  HS65_LH_OAI22X1 U15217 ( .A(n14042), .B(\u_DataPath/rs_ex_i [3]), .C(n14050), 
        .D(\u_DataPath/u_idexreg/N56 ), .Z(n14135) );
  HS65_LH_OAI22X1 U15218 ( .A(n14041), .B(\u_DataPath/rs_ex_i [2]), .C(n14040), 
        .D(\u_DataPath/rs_ex_i [1]), .Z(n14136) );
  HS65_LH_NAND4ABX3 U15219 ( .A(n14140), .B(n14139), .C(n14138), .D(n14137), 
        .Z(n14210) );
  HS65_LH_BFX4 U15220 ( .A(n14034), .Z(n14239) );
  HS65_LH_NAND2AX4 U15221 ( .A(n14142), .B(n14239), .Z(n14141) );
  HS65_LH_BFX4 U15222 ( .A(n14141), .Z(n14240) );
  HS65_LH_NAND2X5 U15223 ( .A(n14239), .B(n14142), .Z(n14238) );
  HS65_LH_BFX4 U15224 ( .A(n14238), .Z(n14242) );
  HS65_LH_OAI222X2 U15225 ( .A(n17611), .B(n17874), .C(n17631), .D(n17262), 
        .E(n17610), .F(n18014), .Z(n15099) );
  HS65_LH_FA1X4 U15226 ( .A0(n9020), .B0(n4411), .CI(n14143), .CO(n14185), 
        .S0(n14112) );
  HS65_LH_MUX21X4 U15227 ( .D0(\u_DataPath/from_alu_data_out_i [17]), .D1(
        \u_DataPath/from_mem_data_out_i [17]), .S0(\u_DataPath/cw_towb_i [0]), 
        .Z(n14145) );
  HS65_LH_CNIVX3 U15228 ( .A(n17478), .Z(n14273) );
  HS65_LH_OAI222X2 U15229 ( .A(n37075), .B(n17618), .C(n14273), .D(n17335), 
        .E(n17616), .F(n17261), .Z(n14261) );
  HS65_LH_OAI222X2 U15230 ( .A(n17611), .B(n17884), .C(n17612), .D(n17261), 
        .E(n17476), .F(n18013), .Z(n15032) );
  HS65_LH_FA1X4 U15231 ( .A0(n17536), .B0(n17500), .CI(n14146), .CO(n14152), 
        .S0(n14147) );
  HS65_LH_MUX21X4 U15232 ( .D0(\u_DataPath/from_alu_data_out_i [16]), .D1(
        \u_DataPath/from_mem_data_out_i [16]), .S0(\u_DataPath/cw_towb_i [0]), 
        .Z(n14148) );
  HS65_LH_OAI222X2 U15233 ( .A(n17611), .B(n17889), .C(n17612), .D(n17370), 
        .E(n17476), .F(n18012), .Z(n14550) );
  HS65_LH_FA1X4 U15234 ( .A0(n17535), .B0(n17492), .CI(n14149), .CO(n14146), 
        .S0(n14150) );
  HS65_LH_MUX21X4 U15235 ( .D0(\u_DataPath/from_alu_data_out_i [20]), .D1(
        \u_DataPath/from_mem_data_out_i [20]), .S0(\u_DataPath/cw_towb_i [0]), 
        .Z(n14151) );
  HS65_LH_FA1X4 U15236 ( .A0(n17872), .B0(n17499), .CI(n14152), .CO(n14203), 
        .S0(n14144) );
  HS65_LH_BFX4 U15237 ( .A(\u_DataPath/cw_towb_i [0]), .Z(n14232) );
  HS65_LH_MUX21X4 U15238 ( .D0(\u_DataPath/from_alu_data_out_i [8]), .D1(
        \u_DataPath/from_mem_data_out_i [8]), .S0(n14232), .Z(n14154) );
  HS65_LH_FA1X4 U15239 ( .A0(n8363), .B0(\u_DataPath/u_idexreg/N33 ), .CI(
        n14155), .CO(n14167), .S0(n14156) );
  HS65_LH_MUX21X4 U15240 ( .D0(\u_DataPath/from_alu_data_out_i [22]), .D1(
        \u_DataPath/from_mem_data_out_i [22]), .S0(\u_DataPath/cw_towb_i [0]), 
        .Z(n14157) );
  HS65_LH_OAI222X2 U15241 ( .A(n17611), .B(n17908), .C(n17631), .D(n17264), 
        .E(n17610), .F(n18010), .Z(n14880) );
  HS65_LH_FA1X4 U15242 ( .A0(n17892), .B0(n17497), .CI(n14158), .CO(n14176), 
        .S0(n14153) );
  HS65_LH_MUX21X4 U15243 ( .D0(\u_DataPath/from_alu_data_out_i [28]), .D1(
        \u_DataPath/from_mem_data_out_i [28]), .S0(n14232), .Z(n14160) );
  HS65_LH_OAI222X2 U15244 ( .A(n37503), .B(n17617), .C(n14273), .D(n32430), 
        .E(n17616), .F(n33785), .Z(n14514) );
  HS65_LH_OAI222X2 U15245 ( .A(n17611), .B(n17915), .C(n17631), .D(n33785), 
        .E(n17610), .F(n18009), .Z(n14852) );
  HS65_LH_FA1X4 U15246 ( .A0(n17906), .B0(n17495), .CI(n14161), .CO(n14194), 
        .S0(n14159) );
  HS65_LH_MUX21X4 U15247 ( .D0(\u_DataPath/from_alu_data_out_i [24]), .D1(
        \u_DataPath/from_mem_data_out_i [24]), .S0(\u_DataPath/cw_towb_i [0]), 
        .Z(n14163) );
  HS65_LH_OAI222X2 U15248 ( .A(n17611), .B(n17919), .C(n17631), .D(
        \u_DataPath/dataOut_exe_i [24]), .E(n17610), .F(n18008), .Z(n14817) );
  HS65_LH_FA1X4 U15249 ( .A0(n17543), .B0(n17493), .CI(n14164), .CO(n14170), 
        .S0(n14165) );
  HS65_LH_MUX21X4 U15250 ( .D0(\u_DataPath/from_alu_data_out_i [9]), .D1(
        \u_DataPath/from_mem_data_out_i [9]), .S0(\u_DataPath/cw_towb_i [0]), 
        .Z(n14166) );
  HS65_LH_OAI222X2 U15251 ( .A(n36058), .B(n17617), .C(n14273), .D(n17346), 
        .E(n17615), .F(n17291), .Z(n14267) );
  HS65_LH_OAI222X2 U15252 ( .A(n14141), .B(n7753), .C(n14239), .D(
        \u_DataPath/dataOut_exe_i [9]), .E(n14238), .F(n5001), .Z(n14785) );
  HS65_LH_FA1X4 U15253 ( .A0(\u_DataPath/pc_4_to_ex_i [9]), .B0(
        \u_DataPath/u_idexreg/N34 ), .CI(n14167), .CO(n14200), .S0(n14168) );
  HS65_LH_MUX21X4 U15254 ( .D0(\u_DataPath/from_alu_data_out_i [25]), .D1(
        \u_DataPath/from_mem_data_out_i [25]), .S0(n14232), .Z(n14169) );
  HS65_LH_OAI222X2 U15255 ( .A(n17611), .B(n17926), .C(n17631), .D(
        \u_DataPath/dataOut_exe_i [25]), .E(n17610), .F(n18006), .Z(n14755) );
  HS65_LH_IVX2 U15256 ( .A(n14755), .Z(n14752) );
  HS65_LH_FA1X4 U15257 ( .A0(n17544), .B0(n17526), .CI(n14170), .CO(n14197), 
        .S0(n14171) );
  HS65_LH_MUX21X4 U15258 ( .D0(\u_DataPath/from_alu_data_out_i [5]), .D1(
        \u_DataPath/from_mem_data_out_i [5]), .S0(n14232), .Z(n14172) );
  HS65_LH_OAI222X2 U15259 ( .A(n17477), .B(n17930), .C(n17612), .D(n17364), 
        .E(n17610), .F(n18004), .Z(n14730) );
  HS65_LH_FA1X4 U15260 ( .A0(\u_DataPath/pc_4_to_ex_i [5]), .B0(
        \u_DataPath/u_idexreg/N30 ), .CI(n14173), .CO(n14143), .S0(n14174) );
  HS65_LH_MUX21X4 U15261 ( .D0(\u_DataPath/from_alu_data_out_i [21]), .D1(
        \u_DataPath/from_mem_data_out_i [21]), .S0(\u_DataPath/cw_towb_i [0]), 
        .Z(n14175) );
  HS65_LH_OAI222X2 U15262 ( .A(n17611), .B(n17934), .C(n17631), .D(n17372), 
        .E(n17610), .F(n18003), .Z(n14709) );
  HS65_LH_FA1X4 U15263 ( .A0(n17540), .B0(n17496), .CI(n14176), .CO(n14161), 
        .S0(n14177) );
  HS65_LH_MUX21X4 U15264 ( .D0(\u_DataPath/from_alu_data_out_i [29]), .D1(
        \u_DataPath/from_mem_data_out_i [29]), .S0(n14232), .Z(n14178) );
  HS65_LH_OAI222X2 U15265 ( .A(n38331), .B(n17617), .C(n14273), .D(n32101), 
        .E(n17616), .F(n33654), .Z(n14513) );
  HS65_LH_FA1X4 U15266 ( .A0(n17914), .B0(n17526), .CI(n14179), .CO(n14191), 
        .S0(n14162) );
  HS65_LH_MUX21X4 U15267 ( .D0(\u_DataPath/from_alu_data_out_i [13]), .D1(
        \u_DataPath/from_mem_data_out_i [13]), .S0(\u_DataPath/cw_towb_i [0]), 
        .Z(n14181) );
  HS65_LH_OAI222X2 U15268 ( .A(n36582), .B(n17617), .C(n17614), .D(n17355), 
        .E(n17615), .F(n17368), .Z(n14263) );
  HS65_LH_OAI222X2 U15269 ( .A(n14141), .B(n7240), .C(n14239), .D(
        \u_DataPath/dataOut_exe_i [13]), .E(n14238), .F(n5308), .Z(n14631) );
  HS65_LH_FA1X4 U15270 ( .A0(n17532), .B0(n17559), .CI(n14182), .CO(n14305), 
        .S0(n14183) );
  HS65_LH_MUX21X4 U15271 ( .D0(\u_DataPath/from_alu_data_out_i [7]), .D1(
        \u_DataPath/from_mem_data_out_i [7]), .S0(n14232), .Z(n14184) );
  HS65_LH_OAI222X2 U15272 ( .A(n14141), .B(n7157), .C(n14239), .D(
        \u_DataPath/dataOut_exe_i [7]), .E(n14238), .F(n5374), .Z(n14613) );
  HS65_LH_FA1X4 U15273 ( .A0(\u_DataPath/pc_4_to_ex_i [7]), .B0(
        \u_DataPath/u_idexreg/N32 ), .CI(n14185), .CO(n14155), .S0(n14186) );
  HS65_LH_MUX21X4 U15274 ( .D0(\u_DataPath/from_alu_data_out_i [12]), .D1(
        \u_DataPath/from_mem_data_out_i [12]), .S0(\u_DataPath/cw_towb_i [0]), 
        .Z(n14187) );
  HS65_LH_FA1X4 U15275 ( .A0(n17531), .B0(n17558), .CI(n14188), .CO(n14182), 
        .S0(n14189) );
  HS65_LH_MUX21X4 U15276 ( .D0(\u_DataPath/from_alu_data_out_i [30]), .D1(
        \u_DataPath/from_mem_data_out_i [30]), .S0(n14232), .Z(n14190) );
  HS65_LH_OAI222X2 U15277 ( .A(n38254), .B(n17617), .C(n14273), .D(n32134), 
        .E(n17615), .F(n33653), .Z(n14511) );
  HS65_LH_OA222X4 U15278 ( .A(n17611), .B(n17954), .C(n17631), .D(n33653), .E(
        n17476), .F(n17362), .Z(n15396) );
  HS65_LH_FA1X4 U15279 ( .A0(n17548), .B0(n18002), .CI(n14191), .CO(n15471), 
        .S0(n14180) );
  HS65_LH_MUX21X4 U15280 ( .D0(\u_DataPath/from_alu_data_out_i [23]), .D1(
        \u_DataPath/from_mem_data_out_i [23]), .S0(\u_DataPath/cw_towb_i [0]), 
        .Z(n14193) );
  HS65_LH_OAI222X2 U15281 ( .A(n17611), .B(n17957), .C(n17631), .D(n33749), 
        .E(n17610), .F(n17999), .Z(n14494) );
  HS65_LH_FA1X4 U15282 ( .A0(n17542), .B0(n17494), .CI(n14194), .CO(n14164), 
        .S0(n14195) );
  HS65_LH_MUX21X4 U15283 ( .D0(\u_DataPath/from_alu_data_out_i [26]), .D1(
        \u_DataPath/from_mem_data_out_i [26]), .S0(n14232), .Z(n14196) );
  HS65_LH_OAI222X2 U15284 ( .A(n17611), .B(n17964), .C(n17631), .D(n33776), 
        .E(n17610), .F(n17360), .Z(n14470) );
  HS65_LH_IVX2 U15285 ( .A(n14470), .Z(n14553) );
  HS65_LH_FA1X4 U15286 ( .A0(n17963), .B0(n17526), .CI(n14197), .CO(n14211), 
        .S0(n14198) );
  HS65_LH_MUX21X4 U15287 ( .D0(\u_DataPath/from_alu_data_out_i [10]), .D1(
        \u_DataPath/from_mem_data_out_i [10]), .S0(\u_DataPath/cw_towb_i [0]), 
        .Z(n14199) );
  HS65_LH_OAI222X2 U15288 ( .A(n14141), .B(n6660), .C(n14239), .D(
        \u_DataPath/dataOut_exe_i [10]), .E(n14238), .F(n5703), .Z(n14409) );
  HS65_LH_FA1X4 U15289 ( .A0(n17967), .B0(n17556), .CI(n17277), .CO(n14207), 
        .S0(n14201) );
  HS65_LH_MUX21X4 U15290 ( .D0(\u_DataPath/from_alu_data_out_i [19]), .D1(
        \u_DataPath/from_mem_data_out_i [19]), .S0(\u_DataPath/cw_towb_i [0]), 
        .Z(n14202) );
  HS65_LH_OAI222X2 U15291 ( .A(n37804), .B(n17618), .C(n14273), .D(n17339), 
        .E(n17616), .F(n17371), .Z(n14260) );
  HS65_LH_OAI222X2 U15292 ( .A(n17611), .B(n17977), .C(n17631), .D(n17371), 
        .E(n17610), .F(n17998), .Z(n14633) );
  HS65_LH_IVX2 U15293 ( .A(n14633), .Z(n14388) );
  HS65_LH_FA1X4 U15294 ( .A0(n17538), .B0(n17498), .CI(n14203), .CO(n14158), 
        .S0(n14204) );
  HS65_LH_MUX21X4 U15295 ( .D0(\u_DataPath/from_alu_data_out_i [11]), .D1(
        \u_DataPath/from_mem_data_out_i [11]), .S0(\u_DataPath/cw_towb_i [0]), 
        .Z(n14205) );
  HS65_LH_OAI222X2 U15296 ( .A(n36495), .B(n17617), .C(n17614), .D(n17349), 
        .E(n17615), .F(n17293), .Z(n14265) );
  HS65_LH_OAI222X2 U15297 ( .A(n14141), .B(n6317), .C(n14239), .D(
        \u_DataPath/dataOut_exe_i [11]), .E(n14238), .F(n5835), .Z(n14616) );
  HS65_LH_FA1X4 U15298 ( .A0(n17530), .B0(n17557), .CI(n14207), .CO(n14188), 
        .S0(n14208) );
  HS65_LH_MUX21X4 U15299 ( .D0(\u_DataPath/from_alu_data_out_i [27]), .D1(
        \u_DataPath/from_mem_data_out_i [27]), .S0(\u_DataPath/cw_towb_i [0]), 
        .Z(n14209) );
  HS65_LH_OAI222X2 U15300 ( .A(n35704), .B(n17618), .C(n14273), .D(n32304), 
        .E(n17616), .F(n33771), .Z(n14243) );
  HS65_LH_OAI222X2 U15301 ( .A(n17611), .B(n17995), .C(n17278), .D(n33771), 
        .E(n17610), .F(n17997), .Z(n14843) );
  HS65_LH_FA1X4 U15302 ( .A0(n17546), .B0(n17526), .CI(n14211), .CO(n14179), 
        .S0(n14212) );
  HS65_LH_MUX21X4 U15303 ( .D0(\u_DataPath/from_alu_data_out_i [1]), .D1(
        \u_DataPath/from_mem_data_out_i [1]), .S0(n14232), .Z(n14214) );
  HS65_LH_MUX21I1X3 U15304 ( .D0(n31993), .D1(n17504), .S0(n17528), .Z(n15500)
         );
  HS65_LH_IVX2 U15305 ( .A(n15500), .Z(n15195) );
  HS65_LH_MUX21X4 U15306 ( .D0(\u_DataPath/from_alu_data_out_i [0]), .D1(
        \u_DataPath/from_mem_data_out_i [0]), .S0(n14232), .Z(n14216) );
  HS65_LH_CNIVX3 U15307 ( .A(\u_DataPath/u_idexreg/N25 ), .Z(n15641) );
  HS65_LH_AND2X4 U15308 ( .A(n15195), .B(n15341), .Z(n14622) );
  HS65_LH_IVX2 U15309 ( .A(n14622), .Z(n15328) );
  HS65_LH_NOR2X2 U15310 ( .A(n15328), .B(n15099), .Z(n14635) );
  HS65_LH_NOR2X2 U15312 ( .A(n14626), .B(n14550), .Z(n14640) );
  HS65_LH_NAND2X2 U15315 ( .A(n14218), .B(n14388), .Z(n14335) );
  HS65_LH_NOR2X2 U15316 ( .A(n15195), .B(n15341), .Z(n14643) );
  HS65_LH_NAND2X2 U15317 ( .A(n14643), .B(n15018), .Z(n14333) );
  HS65_LH_NAND4ABX3 U15318 ( .A(n14635), .B(n14640), .C(n14335), .D(n14333), 
        .Z(n15404) );
  HS65_LH_IVX2 U15319 ( .A(n15404), .Z(n14389) );
  HS65_LH_MUX21X4 U15320 ( .D0(\u_DataPath/from_alu_data_out_i [3]), .D1(
        \u_DataPath/from_mem_data_out_i [3]), .S0(n14232), .Z(n14219) );
  HS65_LH_MUX21I1X3 U15321 ( .D0(n32042), .D1(n17502), .S0(n17528), .Z(n14925)
         );
  HS65_LH_MUX21X4 U15323 ( .D0(\u_DataPath/from_alu_data_out_i [2]), .D1(
        \u_DataPath/from_mem_data_out_i [2]), .S0(n14232), .Z(n14221) );
  HS65_LH_MUX21I1X3 U15324 ( .D0(n31980), .D1(n17503), .S0(n17528), .Z(n15069)
         );
  HS65_LH_NOR2X5 U15325 ( .A(n14037), .B(n15069), .Z(n15329) );
  HS65_LH_MUX21X4 U15326 ( .D0(\u_DataPath/from_alu_data_out_i [4]), .D1(
        \u_DataPath/from_mem_data_out_i [4]), .S0(n14232), .Z(n14223) );
  HS65_LH_IVX4 U15327 ( .A(\u_DataPath/cw_to_ex_i [14]), .Z(n15212) );
  HS65_LH_MUX21I1X3 U15328 ( .D0(n17551), .D1(n32022), .S0(n17608), .Z(n14922)
         );
  HS65_LH_IVX2 U15329 ( .A(n14922), .Z(n14919) );
  HS65_LH_CNIVX3 U15330 ( .A(\u_DataPath/cw_to_ex_i [0]), .Z(n14225) );
  HS65_LH_CNIVX3 U15331 ( .A(n14225), .Z(n14244) );
  HS65_LH_CNIVX3 U15332 ( .A(\u_DataPath/cw_to_ex_i [2]), .Z(n15319) );
  HS65_LH_CNIVX3 U15333 ( .A(\u_DataPath/cw_to_ex_i [1]), .Z(n14278) );
  HS65_LH_NAND2X2 U15334 ( .A(n15319), .B(n14278), .Z(n15380) );
  HS65_LH_NOR3X1 U15335 ( .A(\u_DataPath/cw_to_ex_i [3]), .B(
        \u_DataPath/cw_to_ex_i [4]), .C(n15380), .Z(n14245) );
  HS65_LH_NAND2X2 U15336 ( .A(n14244), .B(n14245), .Z(n14230) );
  HS65_LH_NAND2X2 U15338 ( .A(n15329), .B(n14930), .Z(n15409) );
  HS65_LH_NAND2X2 U15339 ( .A(n14643), .B(n14752), .Z(n14331) );
  HS65_LH_IVX2 U15340 ( .A(n14226), .Z(n14231) );
  HS65_LH_NAND2X2 U15341 ( .A(n14231), .B(n14627), .Z(n14227) );
  HS65_LH_NOR2X2 U15342 ( .A(n15328), .B(n14470), .Z(n14628) );
  HS65_LH_NOR2X2 U15343 ( .A(n14626), .B(n14817), .Z(n14645) );
  HS65_LH_NOR4ABX2 U15344 ( .A(n14331), .B(n14227), .C(n14628), .D(n14645), 
        .Z(n15418) );
  HS65_LH_IVX2 U15346 ( .A(n15075), .Z(n14625) );
  HS65_LH_IVX2 U15347 ( .A(n14930), .Z(n14872) );
  HS65_LH_NOR2X5 U15348 ( .A(n14625), .B(n14872), .Z(n15499) );
  HS65_LH_IVX2 U15349 ( .A(n15499), .Z(n15026) );
  HS65_LH_OAI22X1 U15350 ( .A(n14389), .B(n15409), .C(n15418), .D(n15026), .Z(
        n14297) );
  HS65_LH_IVX2 U15351 ( .A(n14625), .Z(n15039) );
  HS65_LH_CNIVX3 U15352 ( .A(n14626), .Z(n15044) );
  HS65_LH_NOR2X2 U15353 ( .A(n15328), .B(n14852), .Z(n14678) );
  HS65_LH_AOI21X2 U15354 ( .A(n40560), .B(n15044), .C(n14678), .Z(n14228) );
  HS65_LH_NAND2X2 U15355 ( .A(n14643), .B(n14031), .Z(n15400) );
  HS65_LH_NAND3X2 U15356 ( .A(n14228), .B(n14227), .C(n15400), .Z(n14487) );
  HS65_LH_MUX21X4 U15357 ( .D0(\u_DataPath/from_alu_data_out_i [31]), .D1(
        \u_DataPath/from_mem_data_out_i [31]), .S0(n14232), .Z(n15210) );
  HS65_LH_NOR2X2 U15359 ( .A(n15039), .B(n10437), .Z(n14623) );
  HS65_LH_AOI21X2 U15360 ( .A(n15039), .B(n14487), .C(n14623), .Z(n14361) );
  HS65_LH_NOR2X2 U15361 ( .A(\u_DataPath/cw_to_ex_i [2]), .B(n14278), .Z(
        n15374) );
  HS65_LH_CNIVX3 U15362 ( .A(n15374), .Z(n14291) );
  HS65_LH_OR3X4 U15363 ( .A(\u_DataPath/cw_to_ex_i [3]), .B(
        \u_DataPath/cw_to_ex_i [4]), .C(n14291), .Z(n15407) );
  HS65_LH_NOR2X2 U15364 ( .A(n14919), .B(n35213), .Z(n15042) );
  HS65_LH_NAND2X2 U15365 ( .A(n33045), .B(n15042), .Z(n15120) );
  HS65_LH_NAND2X2 U15366 ( .A(n29624), .B(n15331), .Z(n14710) );
  HS65_LH_IVX2 U15367 ( .A(n14710), .Z(n14879) );
  HS65_LH_NOR2X2 U15368 ( .A(n14226), .B(n17254), .Z(n14410) );
  HS65_LH_IVX2 U15369 ( .A(n14643), .Z(n15508) );
  HS65_LH_NOR2X2 U15370 ( .A(n15508), .B(n14730), .Z(n14412) );
  HS65_LH_OAI222X2 U15371 ( .A(n17901), .B(n17611), .C(n17610), .D(n17903), 
        .E(n17612), .F(n17289), .Z(n14921) );
  HS65_LH_NAND2X2 U15372 ( .A(n15044), .B(n14918), .Z(n15510) );
  HS65_LH_MUX21X4 U15373 ( .D0(\u_DataPath/from_alu_data_out_i [6]), .D1(
        \u_DataPath/from_mem_data_out_i [6]), .S0(n14232), .Z(n14233) );
  HS65_LH_OAI222X2 U15374 ( .A(n14141), .B(n9079), .C(n14239), .D(
        \u_DataPath/dataOut_exe_i [6]), .E(n14238), .F(
        \u_DataPath/data_read_ex_1_i [6]), .Z(n15136) );
  HS65_LH_NAND2X2 U15375 ( .A(n14622), .B(n14029), .Z(n14722) );
  HS65_LH_NAND4ABX3 U15376 ( .A(n14410), .B(n14412), .C(n15510), .D(n14722), 
        .Z(n14491) );
  HS65_LH_NOR2X3 U15377 ( .A(n14037), .B(n15245), .Z(n15333) );
  HS65_LH_NAND2X2 U15378 ( .A(n15333), .B(n14930), .Z(n14827) );
  HS65_LH_IVX2 U15379 ( .A(n14827), .Z(n15405) );
  HS65_LH_OAI222X2 U15380 ( .A(n14141), .B(n7075), .C(n14239), .D(
        \u_DataPath/dataOut_exe_i [12]), .E(n14238), .F(
        \u_DataPath/data_read_ex_1_i [12]), .Z(n15238) );
  HS65_LH_NOR2X2 U15381 ( .A(n14626), .B(n17250), .Z(n14728) );
  HS65_LH_MUX21X4 U15382 ( .D0(\u_DataPath/from_alu_data_out_i [14]), .D1(
        \u_DataPath/from_mem_data_out_i [14]), .S0(\u_DataPath/cw_towb_i [0]), 
        .Z(n14234) );
  HS65_LH_OAI222X2 U15383 ( .A(n14141), .B(n6148), .C(n14239), .D(n6170), .E(
        n14238), .F(n6131), .Z(n14365) );
  HS65_LH_NOR2X2 U15384 ( .A(n15328), .B(n17249), .Z(n14641) );
  HS65_LH_MUX21X4 U15385 ( .D0(\u_DataPath/from_alu_data_out_i [15]), .D1(
        \u_DataPath/from_mem_data_out_i [15]), .S0(\u_DataPath/cw_towb_i [0]), 
        .Z(n14235) );
  HS65_LH_OAI222X2 U15386 ( .A(n14141), .B(n6233), .C(n14239), .D(
        \u_DataPath/dataOut_exe_i [15]), .E(n14238), .F(
        \u_DataPath/data_read_ex_1_i [15]), .Z(n14338) );
  HS65_LH_NAND2X2 U15387 ( .A(n14218), .B(n14035), .Z(n14334) );
  HS65_LH_IVX2 U15388 ( .A(n15508), .Z(n15325) );
  HS65_LH_NAND2X2 U15389 ( .A(n15325), .B(n14032), .Z(n14366) );
  HS65_LH_NAND4ABX3 U15390 ( .A(n14728), .B(n14641), .C(n14334), .D(n14366), 
        .Z(n14490) );
  HS65_LH_AOI22X1 U15391 ( .A(n14879), .B(n14491), .C(n15405), .D(n14490), .Z(
        n14236) );
  HS65_LH_OAI21X2 U15392 ( .A(n14361), .B(n15120), .C(n14236), .Z(n14296) );
  HS65_LH_NAND2X2 U15394 ( .A(n14218), .B(n38579), .Z(n15398) );
  HS65_LH_IVX2 U15395 ( .A(n15398), .Z(n15403) );
  HS65_LH_MUXI21X2 U15396 ( .D0(n15403), .D1(n14487), .S0(n15245), .Z(n14382)
         );
  HS65_LH_NOR2X2 U15397 ( .A(n6651), .B(n14382), .Z(n14362) );
  HS65_LH_IVX2 U15398 ( .A(n15042), .Z(n15344) );
  HS65_LH_NOR2X2 U15399 ( .A(n33045), .B(n15344), .Z(n14900) );
  HS65_LH_NAND2X2 U15400 ( .A(n29624), .B(n15039), .Z(n14999) );
  HS65_LH_IVX2 U15401 ( .A(n14999), .Z(n15100) );
  HS65_LH_NOR2X2 U15402 ( .A(n15328), .B(n17253), .Z(n14729) );
  HS65_LH_NOR2X2 U15403 ( .A(n14226), .B(n17252), .Z(n14367) );
  HS65_LH_NAND2X2 U15404 ( .A(n15325), .B(n14545), .Z(n14411) );
  HS65_LH_NAND2X2 U15405 ( .A(n15044), .B(n14030), .Z(n14723) );
  HS65_LH_NAND4ABX3 U15406 ( .A(n14729), .B(n14367), .C(n14411), .D(n14723), 
        .Z(n14489) );
  HS65_LH_AOI22X1 U15407 ( .A(n14362), .B(n14900), .C(n15100), .D(n14489), .Z(
        n14249) );
  HS65_LH_NOR2X2 U15408 ( .A(n35213), .B(n14922), .Z(n15529) );
  HS65_LH_NAND2X2 U15409 ( .A(n32353), .B(n15529), .Z(n15080) );
  HS65_LH_IVX2 U15410 ( .A(n15080), .Z(n15128) );
  HS65_LH_NAND2X4 U15411 ( .A(n38579), .B(n15128), .Z(n15098) );
  HS65_LH_OAI222X2 U15412 ( .A(n17477), .B(n17864), .C(n17612), .D(n17859), 
        .E(n17610), .F(n17356), .Z(n15505) );
  HS65_LH_IVX2 U15413 ( .A(n15505), .Z(n15502) );
  HS65_LH_OAI222X2 U15414 ( .A(n17972), .B(n17611), .C(n17610), .D(n17358), 
        .E(n17612), .F(n17288), .Z(n15507) );
  HS65_LH_AOI22X1 U15415 ( .A(n15502), .B(n14643), .C(n15246), .D(n14231), .Z(
        n14241) );
  HS65_LH_OAI222X2 U15416 ( .A(n17860), .B(n17611), .C(n17612), .D(n17761), 
        .E(n17476), .F(n17862), .Z(n15337) );
  HS65_LH_NAND2X2 U15417 ( .A(n15163), .B(n15044), .Z(n14271) );
  HS65_LH_OAI222X2 U15418 ( .A(n17879), .B(n17611), .C(n17610), .D(n17357), 
        .E(n17612), .F(n17287), .Z(n15062) );
  HS65_LH_NAND2X2 U15419 ( .A(n15324), .B(n14622), .Z(n15511) );
  HS65_LH_NAND3X2 U15420 ( .A(n14241), .B(n14271), .C(n15511), .Z(n14587) );
  HS65_LH_IVX2 U15421 ( .A(n14587), .Z(n14495) );
  HS65_LH_NAND2X2 U15422 ( .A(n29624), .B(n15329), .Z(n14824) );
  HS65_LH_NAND2X2 U15423 ( .A(n14643), .B(n15268), .Z(n14336) );
  HS65_LH_OAI222X2 U15424 ( .A(n17611), .B(n17894), .C(n17631), .D(n17263), 
        .E(n17610), .F(n17359), .Z(n15272) );
  HS65_LH_IVX2 U15425 ( .A(n15272), .Z(\u_DataPath/u_execute/A_inALU_i [20])
         );
  HS65_LH_NAND2X2 U15426 ( .A(n15044), .B(\u_DataPath/u_execute/A_inALU_i [20]), .Z(n14634) );
  HS65_LH_NOR2X2 U15427 ( .A(n15328), .B(n14880), .Z(n14644) );
  HS65_LH_NOR2X2 U15428 ( .A(n14226), .B(n14494), .Z(n14332) );
  HS65_LH_NOR4ABX2 U15429 ( .A(n14336), .B(n14634), .C(n14644), .D(n14332), 
        .Z(n15410) );
  HS65_LH_OAI22X1 U15430 ( .A(n14495), .B(n14824), .C(n15410), .D(n15417), .Z(
        n14248) );
  HS65_LH_MUX21I1X3 U15431 ( .D0(n17991), .D1(n32307), .S0(n17608), .Z(n14520)
         );
  HS65_LH_NAND2AX4 U15432 ( .A(\u_DataPath/cw_to_ex_i [4]), .B(
        \u_DataPath/cw_to_ex_i [3]), .Z(n15385) );
  HS65_LH_NAND2X4 U15433 ( .A(n15501), .B(n14225), .Z(n15408) );
  HS65_LH_CNIVX3 U15434 ( .A(n15408), .Z(n14821) );
  HS65_LH_IVX2 U15435 ( .A(n14520), .Z(n14517) );
  HS65_LH_NAND2X2 U15436 ( .A(n14245), .B(n14225), .Z(n14966) );
  HS65_LH_CBI4I1X3 U15437 ( .A(n35562), .B(n14517), .C(n17515), .D(n14627), 
        .Z(n14246) );
  HS65_LH_OAI21X2 U15438 ( .A(n14520), .B(n17523), .C(n14246), .Z(n14247) );
  HS65_LH_MUX21I1X3 U15439 ( .D0(n32218), .D1(n29693), .S0(n17528), .Z(n14468)
         );
  HS65_LH_MUX21I1X3 U15440 ( .D0(n29692), .D1(n32243), .S0(n17608), .Z(n14756)
         );
  HS65_LH_MUX21I1X3 U15441 ( .D0(n32262), .D1(n29693), .S0(n17528), .Z(n14820)
         );
  HS65_LH_MUX21I1X3 U15442 ( .D0(n17527), .D1(n32287), .S0(n17608), .Z(n14288)
         );
  HS65_LH_MUX21I1X3 U15443 ( .D0(n31580), .D1(n17527), .S0(n17528), .Z(n14287)
         );
  HS65_LH_MUX21I1X3 U15444 ( .D0(n17527), .D1(n31602), .S0(n17608), .Z(n15269)
         );
  HS65_LH_MUX21I1X3 U15445 ( .D0(n31627), .D1(n29692), .S0(n17528), .Z(n15271)
         );
  HS65_LH_MUX21I1X3 U15446 ( .D0(n17527), .D1(n31648), .S0(n17608), .Z(n14386)
         );
  HS65_LH_MUX21I1X3 U15447 ( .D0(n17527), .D1(n31694), .S0(n17608), .Z(n15033)
         );
  HS65_LH_MUX21I1X3 U15448 ( .D0(n31715), .D1(n17527), .S0(n17528), .Z(n14998)
         );
  HS65_LH_OAI222X2 U15449 ( .A(n36314), .B(n17617), .C(n14273), .D(n17353), 
        .E(n17615), .F(n17369), .Z(n14301) );
  HS65_LH_MUX21I1X3 U15450 ( .D0(n18158), .D1(n14301), .S0(n17608), .Z(n14349)
         );
  HS65_LH_AOI222X2 U15451 ( .A(n6145), .B(n15209), .C(n15208), .D(n6099), .E(
        n15207), .F(n6170), .Z(n14304) );
  HS65_LH_MUX21I1X3 U15452 ( .D0(n17247), .D1(n17560), .S0(n17528), .Z(n14309)
         );
  HS65_LH_MUX21I1X3 U15453 ( .D0(n17559), .D1(n14263), .S0(n17608), .Z(n14632)
         );
  HS65_LH_IVX2 U15454 ( .A(n17250), .Z(\u_DataPath/u_execute/A_inALU_i [12])
         );
  HS65_LH_MUX21I1X3 U15455 ( .D0(n14264), .D1(n17558), .S0(n17528), .Z(n15237)
         );
  HS65_LH_MUX21I1X3 U15456 ( .D0(n17557), .D1(n14265), .S0(n17608), .Z(n14285)
         );
  HS65_LH_MUX21I1X3 U15457 ( .D0(n14266), .D1(n17556), .S0(n17528), .Z(n14433)
         );
  HS65_LH_MUX21I1X3 U15458 ( .D0(n17555), .D1(n14267), .S0(n17608), .Z(n14784)
         );
  HS65_LH_MUX21I1X3 U15459 ( .D0(n14268), .D1(n17554), .S0(n17528), .Z(n15239)
         );
  HS65_LH_MUX21I1X3 U15460 ( .D0(n17553), .D1(n14269), .S0(n17608), .Z(n14586)
         );
  HS65_LH_MUX21I1X3 U15461 ( .D0(n17501), .D1(n14270), .S0(n17608), .Z(n14731)
         );
  HS65_LH_NAND2X2 U15462 ( .A(n15163), .B(n15341), .Z(n15512) );
  HS65_LH_AOI22X1 U15463 ( .A(n15195), .B(n15512), .C(n14271), .D(n15505), .Z(
        n15087) );
  HS65_LH_PAOI2X1 U15464 ( .A(n15324), .B(n15087), .P(n15069), .Z(n14419) );
  HS65_LH_PAOI2X1 U15465 ( .A(n14037), .B(n14419), .P(n15507), .Z(n14912) );
  HS65_LH_PAOI2X1 U15466 ( .A(n14918), .B(n14919), .P(n14912), .Z(n14738) );
  HS65_LH_PAOI2X1 U15467 ( .A(n14731), .B(n14738), .P(n14730), .Z(n15150) );
  HS65_LH_OAI222X2 U15468 ( .A(n35736), .B(n17617), .C(n14273), .D(n17347), 
        .E(n17615), .F(n17365), .Z(n14275) );
  HS65_LH_MUX21I1X3 U15469 ( .D0(n14275), .D1(n17552), .S0(n17528), .Z(n15134)
         );
  HS65_LH_PAOI2X1 U15470 ( .A(n14029), .B(n15150), .P(n15134), .Z(n14600) );
  HS65_LH_PAOI2X1 U15471 ( .A(n14586), .B(n14600), .P(n17254), .Z(n14946) );
  HS65_LH_PAOI2X1 U15472 ( .A(n14030), .B(n15239), .P(n14946), .Z(n14791) );
  HS65_LH_PAOI2X1 U15473 ( .A(n14784), .B(n14791), .P(n17256), .Z(n14439) );
  HS65_LH_PAOI2X1 U15474 ( .A(n14033), .B(n14433), .P(n14439), .Z(n14372) );
  HS65_LH_PAOI2X1 U15475 ( .A(n14285), .B(n14372), .P(n17252), .Z(n14570) );
  HS65_LH_PAOI2X1 U15476 ( .A(\u_DataPath/u_execute/A_inALU_i [12]), .B(n15237), .P(n14570), .Z(n14610) );
  HS65_LH_PAOI2X1 U15477 ( .A(n14632), .B(n14610), .P(n32851), .Z(n14321) );
  HS65_LH_PAOI2X1 U15478 ( .A(n14036), .B(n14309), .P(n14321), .Z(n14348) );
  HS65_LH_PAOI2X1 U15479 ( .A(n14349), .B(n14348), .P(n32625), .Z(n15009) );
  HS65_LH_PAOI2X1 U15480 ( .A(n14997), .B(n14998), .P(n15009), .Z(n15023) );
  HS65_LH_PAOI2X1 U15481 ( .A(n15033), .B(n15032), .P(n15023), .Z(n15113) );
  HS65_LH_MUX21I1X3 U15482 ( .D0(n31671), .D1(n17527), .S0(n17528), .Z(n15095)
         );
  HS65_LH_PAOI2X1 U15483 ( .A(n15096), .B(n15113), .P(n15095), .Z(n14398) );
  HS65_LH_PAOI2X1 U15484 ( .A(n14386), .B(n14398), .P(n14633), .Z(n14973) );
  HS65_LH_PAOI2X1 U15485 ( .A(\u_DataPath/u_execute/A_inALU_i [20]), .B(n15271), .P(n14973), .Z(n14704) );
  HS65_LH_PAOI2X1 U15486 ( .A(n15269), .B(n14704), .P(n14709), .Z(n14890) );
  HS65_LH_PAOI2X1 U15487 ( .A(n14559), .B(n14287), .P(n14890), .Z(n14502) );
  HS65_LH_PAOI2X1 U15488 ( .A(n14288), .B(n14494), .P(n14502), .Z(n14830) );
  HS65_LH_PAOI2X1 U15489 ( .A(n14822), .B(n14820), .P(n14830), .Z(n14762) );
  HS65_LH_PAOI2X1 U15490 ( .A(n14756), .B(n14762), .P(n14755), .Z(n14458) );
  HS65_LH_PAOI2X1 U15491 ( .A(n14553), .B(n14468), .P(n14458), .Z(n14519) );
  HS65_LH_NOR2X2 U15492 ( .A(\u_DataPath/cw_to_ex_i [3]), .B(
        \u_DataPath/cw_to_ex_i [4]), .Z(n14277) );
  HS65_LH_NAND2X2 U15493 ( .A(n14277), .B(\u_DataPath/cw_to_ex_i [2]), .Z(
        n15709) );
  HS65_LH_OR2X4 U15494 ( .A(\u_DataPath/cw_to_ex_i [1]), .B(n15709), .Z(n15149) );
  HS65_LH_BFX4 U15495 ( .A(n15149), .Z(n15495) );
  HS65_LH_OR2X4 U15496 ( .A(n14278), .B(n15709), .Z(n15720) );
  HS65_LH_BFX4 U15497 ( .A(n15720), .Z(n15393) );
  HS65_LH_IVX2 U15498 ( .A(n14820), .Z(n14818) );
  HS65_LH_NOR2X2 U15499 ( .A(n14818), .B(n14822), .Z(n15234) );
  HS65_LH_IVX2 U15500 ( .A(n15269), .Z(n14707) );
  HS65_LH_NOR2X2 U15501 ( .A(n14707), .B(n14709), .Z(n14286) );
  HS65_LH_IVX2 U15502 ( .A(n15271), .Z(n14976) );
  HS65_LH_NOR2X2 U15503 ( .A(n15095), .B(n15099), .Z(n15116) );
  HS65_LH_AOI21X2 U15504 ( .A(n14388), .B(n14386), .C(n15116), .Z(n15273) );
  HS65_LH_NOR2X2 U15505 ( .A(n14550), .B(n14998), .Z(n15019) );
  HS65_LH_AOI21X2 U15506 ( .A(n15033), .B(n15018), .C(n15019), .Z(n15276) );
  HS65_LH_NOR2X2 U15507 ( .A(n17249), .B(n14309), .Z(n14343) );
  HS65_LH_AOI21X2 U15508 ( .A(n14349), .B(n14035), .C(n14343), .Z(n15255) );
  HS65_LH_IVX2 U15509 ( .A(n14309), .Z(n14311) );
  HS65_LH_NOR2X2 U15510 ( .A(n14036), .B(n14311), .Z(n14323) );
  HS65_LH_NOR2X2 U15511 ( .A(n14032), .B(n14632), .Z(n14608) );
  HS65_LH_NOR2X2 U15512 ( .A(n14323), .B(n14608), .Z(n15258) );
  HS65_LH_NAND2X2 U15513 ( .A(n14032), .B(n14632), .Z(n15236) );
  HS65_LH_IVX2 U15514 ( .A(n15237), .Z(n15252) );
  HS65_LH_IVX2 U15515 ( .A(n14285), .Z(n14279) );
  HS65_LH_NOR2X2 U15516 ( .A(n17252), .B(n14279), .Z(n15262) );
  HS65_LH_NOR2X2 U15517 ( .A(n17253), .B(n14433), .Z(n14441) );
  HS65_LH_NOR2X2 U15518 ( .A(n15262), .B(n14441), .Z(n15300) );
  HS65_LH_NAND2X2 U15519 ( .A(n17253), .B(n14433), .Z(n15298) );
  HS65_LH_IVX2 U15520 ( .A(n15239), .Z(n14943) );
  HS65_LH_NOR2X2 U15521 ( .A(n15245), .B(n15324), .Z(n14406) );
  HS65_LH_AOI21X2 U15522 ( .A(n6651), .B(n15507), .C(n14406), .Z(n15244) );
  HS65_LH_NAND2X2 U15523 ( .A(n15337), .B(n15341), .Z(n15513) );
  HS65_LH_PAOI2X1 U15524 ( .A(n15502), .B(n15195), .P(n15513), .Z(n15086) );
  HS65_LH_OAI21X2 U15525 ( .A(n15062), .B(n15069), .C(n15086), .Z(n14407) );
  HS65_LH_NOR2X2 U15526 ( .A(n6651), .B(n15507), .Z(n15242) );
  HS65_LH_AOI21X2 U15527 ( .A(n15244), .B(n14407), .C(n15242), .Z(n14913) );
  HS65_LH_IVX2 U15528 ( .A(n15134), .Z(n15147) );
  HS65_LH_NAND2X2 U15529 ( .A(n14029), .B(n15147), .Z(n15146) );
  HS65_LH_IVX2 U15530 ( .A(n15146), .Z(n14280) );
  HS65_LH_AOI21X2 U15531 ( .A(n14586), .B(n14583), .C(n14280), .Z(n14282) );
  HS65_LH_IVX2 U15532 ( .A(n14731), .Z(n14733) );
  HS65_LH_NAND2X2 U15533 ( .A(n14730), .B(n14733), .Z(n15143) );
  HS65_LH_OAI21X2 U15534 ( .A(n14029), .B(n15147), .C(n15143), .Z(n14578) );
  HS65_LH_NOR2X2 U15535 ( .A(n14583), .B(n14586), .Z(n14281) );
  HS65_LH_AOI21X2 U15536 ( .A(n14282), .B(n14578), .C(n14281), .Z(n14283) );
  HS65_LH_NAND2X2 U15537 ( .A(n14919), .B(n14921), .Z(n14910) );
  HS65_LH_NOR2X2 U15538 ( .A(n14919), .B(n14921), .Z(n14911) );
  HS65_LH_NOR2X2 U15539 ( .A(n14730), .B(n14733), .Z(n15145) );
  HS65_LH_IVX2 U15540 ( .A(n14282), .Z(n14284) );
  HS65_LH_OAI31X1 U15541 ( .A(n14911), .B(n15145), .C(n14284), .D(n14283), .Z(
        n15247) );
  HS65_LH_OAI21X2 U15542 ( .A(n14913), .B(n15248), .C(n15247), .Z(n14944) );
  HS65_LH_AOI21X2 U15543 ( .A(n14030), .B(n14943), .C(n14944), .Z(n14790) );
  HS65_LH_NOR2X2 U15544 ( .A(n14545), .B(n14784), .Z(n15301) );
  HS65_LH_AOI21X2 U15545 ( .A(n17260), .B(n15239), .C(n15301), .Z(n15299) );
  HS65_LH_IVX2 U15546 ( .A(n15299), .Z(n15253) );
  HS65_LH_NAND2X2 U15547 ( .A(n14545), .B(n14784), .Z(n15254) );
  HS65_LH_OAI21X2 U15548 ( .A(n14790), .B(n15253), .C(n15254), .Z(n14438) );
  HS65_LH_NAND2X2 U15549 ( .A(n15298), .B(n14438), .Z(n14368) );
  HS65_LH_NOR2X2 U15550 ( .A(n14358), .B(n14285), .Z(n15306) );
  HS65_LH_AOI21X2 U15551 ( .A(n15300), .B(n14368), .C(n15306), .Z(n14569) );
  HS65_LH_PAOI2X1 U15552 ( .A(\u_DataPath/u_execute/A_inALU_i [12]), .B(n15252), .P(n14569), .Z(n14612) );
  HS65_LH_NAND2X2 U15553 ( .A(n15236), .B(n14612), .Z(n14318) );
  HS65_LH_NAND2X2 U15554 ( .A(n15258), .B(n14318), .Z(n14344) );
  HS65_LH_NOR2X2 U15555 ( .A(n14035), .B(n14349), .Z(n15251) );
  HS65_LH_AOI21X2 U15556 ( .A(n15255), .B(n14344), .C(n15251), .Z(n15008) );
  HS65_LH_NAND2X2 U15557 ( .A(n14550), .B(n14998), .Z(n15284) );
  HS65_LH_NAND2X2 U15558 ( .A(n15008), .B(n15284), .Z(n15020) );
  HS65_LH_NOR2X2 U15559 ( .A(n15018), .B(n15033), .Z(n15265) );
  HS65_LH_AOI21X2 U15560 ( .A(n15276), .B(n15020), .C(n15265), .Z(n15115) );
  HS65_LH_NAND2X2 U15561 ( .A(n15095), .B(n15099), .Z(n15266) );
  HS65_LH_NAND2X2 U15562 ( .A(n15115), .B(n15266), .Z(n14383) );
  HS65_LH_NOR2X2 U15563 ( .A(n14386), .B(n14388), .Z(n15274) );
  HS65_LH_AOI21X2 U15564 ( .A(n15273), .B(n14383), .C(n15274), .Z(n14975) );
  HS65_LH_PAOI2X1 U15565 ( .A(n14976), .B(\u_DataPath/u_execute/A_inALU_i [20]), .P(n14975), .Z(n14701) );
  HS65_LH_IVX2 U15566 ( .A(n14286), .Z(n15264) );
  HS65_LH_OAI21X2 U15567 ( .A(n15269), .B(n15268), .C(n15264), .Z(n14713) );
  HS65_LH_NOR2X2 U15568 ( .A(n14701), .B(n14713), .Z(n14700) );
  HS65_LH_NOR2X2 U15569 ( .A(n14286), .B(n14700), .Z(n14891) );
  HS65_LH_IVX2 U15570 ( .A(n14287), .Z(n14881) );
  HS65_LH_NOR2X2 U15571 ( .A(n14559), .B(n14881), .Z(n14888) );
  HS65_LH_NOR2X2 U15572 ( .A(n14891), .B(n14888), .Z(n14289) );
  HS65_LH_NAND2X2 U15573 ( .A(n14288), .B(n14642), .Z(n14501) );
  HS65_LH_NAND2X2 U15574 ( .A(n14559), .B(n14881), .Z(n14889) );
  HS65_LH_NAND2X2 U15575 ( .A(n14501), .B(n14889), .Z(n15263) );
  HS65_LH_IVX2 U15576 ( .A(n14288), .Z(n14492) );
  HS65_LH_NAND2X2 U15577 ( .A(n14492), .B(n14494), .Z(n15277) );
  HS65_LH_OAI21X2 U15578 ( .A(n14289), .B(n15263), .C(n15277), .Z(n14831) );
  HS65_LH_NOR2X2 U15579 ( .A(n15234), .B(n14831), .Z(n14456) );
  HS65_LH_NAND2X2 U15580 ( .A(n14756), .B(n14752), .Z(n14761) );
  HS65_LH_NAND2X2 U15581 ( .A(n14818), .B(n14822), .Z(n14829) );
  HS65_LH_NAND2X2 U15582 ( .A(n14761), .B(n14829), .Z(n15291) );
  HS65_LH_NOR2X2 U15583 ( .A(n14456), .B(n15291), .Z(n14515) );
  HS65_LH_IVX2 U15584 ( .A(n14468), .Z(n14461) );
  HS65_LH_IVX2 U15585 ( .A(n14756), .Z(n14751) );
  HS65_LH_NAND2X2 U15586 ( .A(n14751), .B(n14755), .Z(n14760) );
  HS65_LH_OAI21X2 U15587 ( .A(n14461), .B(n14553), .C(n14760), .Z(n15233) );
  HS65_LH_NAND2X2 U15588 ( .A(n14461), .B(n14553), .Z(n14516) );
  HS65_LH_OAI21X2 U15589 ( .A(n14515), .B(n15233), .C(n14516), .Z(n14290) );
  HS65_LH_OAI22X1 U15590 ( .A(n14519), .B(n32759), .C(n33067), .D(n14290), .Z(
        n14294) );
  HS65_LH_NAND2X2 U15591 ( .A(n14517), .B(n14843), .Z(n15235) );
  HS65_LH_OAI21X2 U15592 ( .A(n14843), .B(n14517), .C(n15235), .Z(n15219) );
  HS65_LH_CNIVX3 U15593 ( .A(n15393), .Z(n15514) );
  HS65_LH_CNIVX3 U15594 ( .A(n15495), .Z(n15397) );
  HS65_LH_AOI22X1 U15595 ( .A(n32629), .B(n14290), .C(n32748), .D(n14519), .Z(
        n14292) );
  HS65_LH_NAND3X2 U15596 ( .A(n14292), .B(n17638), .C(n15219), .Z(n14293) );
  HS65_LH_OAI21X2 U15597 ( .A(n14294), .B(n15219), .C(n14293), .Z(n14295) );
  HS65_LH_NAND4ABX3 U15598 ( .A(n14297), .B(n14296), .C(n32096), .D(n14295), 
        .Z(n15574) );
  HS65_LH_NAND3X2 U15599 ( .A(n8860), .B(n6650), .C(
        \u_DataPath/pc_4_to_ex_i [4]), .Z(n14941) );
  HS65_LH_CNIVX3 U15600 ( .A(\u_DataPath/pc_4_to_ex_i [5]), .Z(n14720) );
  HS65_LH_NOR2X2 U15601 ( .A(n14941), .B(n14720), .Z(n15160) );
  HS65_LH_NAND2X2 U15602 ( .A(n15160), .B(n9020), .Z(n15159) );
  HS65_LH_CNIVX3 U15603 ( .A(\u_DataPath/pc_4_to_ex_i [7]), .Z(n14576) );
  HS65_LH_NOR2X2 U15604 ( .A(n15159), .B(n14576), .Z(n14963) );
  HS65_LH_NAND2X2 U15605 ( .A(n14963), .B(n8363), .Z(n14962) );
  HS65_LH_CNIVX3 U15606 ( .A(\u_DataPath/pc_4_to_ex_i [9]), .Z(n14800) );
  HS65_LH_NOR2X2 U15607 ( .A(n14962), .B(n14800), .Z(n14799) );
  HS65_LH_NAND2X2 U15608 ( .A(n14799), .B(n6703), .Z(n14450) );
  HS65_LH_CNIVX3 U15609 ( .A(\u_DataPath/pc_4_to_ex_i [11]), .Z(n14356) );
  HS65_LH_NOR2X2 U15610 ( .A(n14450), .B(n14356), .Z(n14542) );
  HS65_LH_NAND2X2 U15611 ( .A(n14542), .B(\u_DataPath/pc_4_to_ex_i [12]), .Z(
        n14606) );
  HS65_LH_NOR2X2 U15612 ( .A(n14606), .B(n14605), .Z(n14604) );
  HS65_LH_NAND2X2 U15613 ( .A(n14604), .B(n6189), .Z(n14329) );
  HS65_LH_CNIVX3 U15614 ( .A(\u_DataPath/pc_4_to_ex_i [15]), .Z(n14298) );
  HS65_LH_NOR2X2 U15615 ( .A(n14329), .B(n6311), .Z(n15015) );
  HS65_LH_NAND2X2 U15616 ( .A(n15015), .B(\u_DataPath/pc_4_to_ex_i [16]), .Z(
        n15053) );
  HS65_LH_CNIVX3 U15617 ( .A(\u_DataPath/pc_4_to_ex_i [17]), .Z(n15052) );
  HS65_LH_NOR2X2 U15618 ( .A(n15053), .B(n15052), .Z(n15123) );
  HS65_LH_NAND2X2 U15619 ( .A(n17465), .B(n17872), .Z(n15122) );
  HS65_LH_CNIVX3 U15620 ( .A(\u_DataPath/pc_4_to_ex_i [19]), .Z(n14380) );
  HS65_LH_NOR2X2 U15621 ( .A(n15122), .B(n17597), .Z(n14988) );
  HS65_LH_NAND2X2 U15622 ( .A(n14988), .B(n17892), .Z(n14987) );
  HS65_LH_CNIVX3 U15623 ( .A(\u_DataPath/pc_4_to_ex_i [21]), .Z(n14696) );
  HS65_LH_NOR2X2 U15624 ( .A(n14987), .B(n17596), .Z(n14906) );
  HS65_LH_NAND2X2 U15625 ( .A(n14906), .B(n17906), .Z(n14905) );
  HS65_LH_CNIVX3 U15626 ( .A(\u_DataPath/pc_4_to_ex_i [23]), .Z(n14484) );
  HS65_LH_NOR2X2 U15627 ( .A(n14905), .B(n17595), .Z(n14839) );
  HS65_LH_NAND2X2 U15628 ( .A(n14839), .B(n17543), .Z(n14838) );
  HS65_LH_CNIVX3 U15629 ( .A(\u_DataPath/pc_4_to_ex_i [25]), .Z(n14749) );
  HS65_LH_NOR2X2 U15630 ( .A(n14838), .B(n17594), .Z(n14748) );
  HS65_LH_NAND2X2 U15631 ( .A(n14748), .B(n17963), .Z(n14481) );
  HS65_LH_CNIVX3 U15632 ( .A(\u_DataPath/pc_4_to_ex_i [27]), .Z(n14299) );
  HS65_LH_NOR2X2 U15633 ( .A(n14481), .B(n40472), .Z(n14875) );
  HS65_LH_FA1X4 U15634 ( .A0(n17534), .B0(n18158), .CI(n14302), .CO(n14149), 
        .S0(n14303) );
  HS65_LH_FA1X4 U15635 ( .A0(n17986), .B0(n17560), .CI(n14305), .CO(n14302), 
        .S0(n14306) );
  HS65_LH_NAND2X2 U15636 ( .A(n14218), .B(n40560), .Z(n14527) );
  HS65_LH_OAI21X2 U15637 ( .A(n14218), .B(n10437), .C(n14527), .Z(n15076) );
  HS65_LH_AOI21X2 U15638 ( .A(n15039), .B(n15076), .C(n14623), .Z(n14534) );
  HS65_LH_NOR2X5 U15639 ( .A(n14625), .B(n15344), .Z(n15525) );
  HS65_LH_NAND2X2 U15640 ( .A(n14218), .B(n14036), .Z(n14317) );
  HS65_LH_NAND2X2 U15641 ( .A(n15044), .B(n15018), .Z(n14808) );
  HS65_LH_NOR2X2 U15642 ( .A(n15508), .B(n14550), .Z(n14467) );
  HS65_LH_NOR2X2 U15643 ( .A(n15328), .B(n32625), .Z(n14805) );
  HS65_LH_NOR4ABX2 U15644 ( .A(n14317), .B(n14808), .C(n14467), .D(n14805), 
        .Z(n14431) );
  HS65_LH_IVX2 U15645 ( .A(n14431), .Z(n15138) );
  HS65_LH_IVX2 U15646 ( .A(n15329), .Z(n14897) );
  HS65_LH_NOR2X2 U15648 ( .A(n14226), .B(n14880), .Z(n14471) );
  HS65_LH_NOR2X2 U15649 ( .A(n15508), .B(n14817), .Z(n14454) );
  HS65_LH_NAND2X2 U15650 ( .A(n14622), .B(n14642), .Z(n14813) );
  HS65_LH_NAND2X2 U15651 ( .A(n15044), .B(n14752), .Z(n14844) );
  HS65_LH_NAND4ABX3 U15652 ( .A(n14471), .B(n14454), .C(n14813), .D(n14844), 
        .Z(n15073) );
  HS65_LH_AOI22X1 U15653 ( .A(n15525), .B(n15138), .C(n15517), .D(n15073), .Z(
        n14315) );
  HS65_LH_IVX2 U15654 ( .A(n15331), .Z(n14547) );
  HS65_LH_NOR2X2 U15655 ( .A(n15508), .B(n15272), .Z(n14472) );
  HS65_LH_NOR2X2 U15656 ( .A(n14626), .B(n14709), .Z(n14815) );
  HS65_LH_NAND2X2 U15657 ( .A(n14218), .B(n15096), .Z(n14466) );
  HS65_LH_NAND2X2 U15658 ( .A(n14622), .B(n14388), .Z(n14807) );
  HS65_LH_NAND4ABX3 U15659 ( .A(n14472), .B(n14815), .C(n14466), .D(n14807), 
        .Z(n15129) );
  HS65_LH_AND2X4 U15660 ( .A(n15333), .B(n15042), .Z(n15497) );
  HS65_LH_IVX2 U15661 ( .A(n14622), .Z(n14621) );
  HS65_LH_NOR2X2 U15662 ( .A(n14226), .B(n14470), .Z(n14453) );
  HS65_LH_NOR2X2 U15663 ( .A(n15508), .B(n14852), .Z(n14526) );
  HS65_LH_AOI211X1 U15664 ( .A(n14031), .B(n15044), .C(n14453), .D(n14526), 
        .Z(n14308) );
  HS65_LH_OAI21X2 U15665 ( .A(n14621), .B(n14843), .C(n14308), .Z(n15074) );
  HS65_LH_AOI22X1 U15666 ( .A(n13892), .B(n15129), .C(n15497), .D(n15074), .Z(
        n14314) );
  HS65_LH_NAND2X2 U15667 ( .A(n14036), .B(n14309), .Z(n14310) );
  HS65_LH_OAI21X2 U15668 ( .A(n10437), .B(n14621), .C(n14527), .Z(n15078) );
  HS65_LH_IVX2 U15669 ( .A(n15078), .Z(n14895) );
  HS65_LH_NAND2X2 U15670 ( .A(n17607), .B(n15529), .Z(n15079) );
  HS65_LH_IVX2 U15671 ( .A(n15079), .Z(n15126) );
  HS65_LH_NAND2X2 U15672 ( .A(n15039), .B(n15126), .Z(n14636) );
  HS65_LH_OAI22X1 U15673 ( .A(n14310), .B(n17471), .C(n14895), .D(n14636), .Z(
        n14313) );
  HS65_LH_CNIVX3 U15674 ( .A(n15414), .Z(n15506) );
  HS65_LH_CBI4I6X2 U15675 ( .A(n14311), .B(n17523), .C(n17249), .D(n33880), 
        .Z(n14312) );
  HS65_LH_NOR4ABX2 U15676 ( .A(n14315), .B(n14314), .C(n14313), .D(n14312), 
        .Z(n14316) );
  HS65_LH_NOR2X2 U15677 ( .A(n14621), .B(n17256), .Z(n14928) );
  HS65_LH_NOR2X2 U15678 ( .A(n14226), .B(n17253), .Z(n14446) );
  HS65_LH_NAND2X2 U15679 ( .A(n15325), .B(n14030), .Z(n15061) );
  HS65_LH_NAND2X2 U15680 ( .A(n15044), .B(n14583), .Z(n14915) );
  HS65_LH_NAND4ABX3 U15681 ( .A(n14928), .B(n14446), .C(n15061), .D(n14915), 
        .Z(n15101) );
  HS65_LH_NOR2X2 U15682 ( .A(n14626), .B(n17252), .Z(n14929) );
  HS65_LH_NOR2X2 U15683 ( .A(n15328), .B(n32851), .Z(n14558) );
  HS65_LH_NAND2X2 U15684 ( .A(n15325), .B(\u_DataPath/u_execute/A_inALU_i [12]), .Z(n14445) );
  HS65_LH_NAND4ABX3 U15685 ( .A(n14929), .B(n14558), .C(n14317), .D(n14445), 
        .Z(n15103) );
  HS65_LH_NOR2X2 U15686 ( .A(n14626), .B(n15507), .Z(n15348) );
  HS65_LH_NOR2X2 U15687 ( .A(n14621), .B(n14730), .Z(n14917) );
  HS65_LH_NAND2X2 U15688 ( .A(n14218), .B(n14029), .Z(n15057) );
  HS65_LH_NAND2X2 U15689 ( .A(n15325), .B(n14918), .Z(n15082) );
  HS65_LH_NAND4ABX3 U15690 ( .A(n15348), .B(n14917), .C(n15057), .D(n15082), 
        .Z(n15131) );
  HS65_LH_NOR2X2 U15691 ( .A(n15337), .B(n15341), .Z(n15335) );
  HS65_LH_AOI21X2 U15692 ( .A(n15502), .B(n15195), .C(n15335), .Z(n15241) );
  HS65_LH_MUXI21X2 U15693 ( .D0(n15241), .D1(n15062), .S0(n14218), .Z(n15132)
         );
  HS65_LH_MX41X4 U15694 ( .D0(n15101), .S0(n15331), .D1(n15103), .S1(n15039), 
        .D2(n15131), .S2(n15329), .D3(n15132), .S3(n15333), .Z(n14537) );
  HS65_LH_CNIVX3 U15695 ( .A(n15393), .Z(n15493) );
  HS65_LH_NOR2AX3 U15696 ( .A(n14318), .B(n14608), .Z(n14320) );
  HS65_LH_OAI21X2 U15697 ( .A(n14321), .B(n17468), .C(n17638), .Z(n14319) );
  HS65_LH_AOI21X2 U15698 ( .A(n17591), .B(n14320), .C(n14319), .Z(n14325) );
  HS65_LH_IVX2 U15699 ( .A(n14320), .Z(n14322) );
  HS65_LH_AOI22X1 U15700 ( .A(n32629), .B(n14322), .C(n32748), .D(n14321), .Z(
        n14324) );
  HS65_LH_NOR2X2 U15701 ( .A(n14323), .B(n14343), .Z(n15216) );
  HS65_LH_MUXI21X2 U15702 ( .D0(n14325), .D1(n14324), .S0(n15216), .Z(n14326)
         );
  HS65_LH_AOI21X2 U15703 ( .A(n14930), .B(n14537), .C(n14326), .Z(n14327) );
  HS65_LH_MX41X4 U15704 ( .D0(n14490), .S0(n15039), .D1(n14489), .S1(n15331), 
        .D2(n14491), .S2(n15329), .D3(n14587), .S3(n15333), .Z(n15421) );
  HS65_LH_NOR2X2 U15705 ( .A(n14621), .B(n14817), .Z(n14667) );
  HS65_LH_NAND2X2 U15706 ( .A(n15044), .B(n14553), .Z(n14677) );
  HS65_LH_NAND4ABX3 U15707 ( .A(n14332), .B(n14667), .C(n14331), .D(n14677), 
        .Z(n14486) );
  HS65_LH_AOI22X1 U15708 ( .A(n15517), .B(n14486), .C(n15497), .D(n14487), .Z(
        n14354) );
  HS65_LH_NOR2X2 U15709 ( .A(n14626), .B(n15099), .Z(n14671) );
  HS65_LH_NOR2X2 U15710 ( .A(n14621), .B(n14550), .Z(n14664) );
  HS65_LH_NAND4ABX3 U15711 ( .A(n14671), .B(n14664), .C(n14334), .D(n14333), 
        .Z(n14589) );
  HS65_LH_NOR2X2 U15712 ( .A(n14626), .B(n14880), .Z(n14668) );
  HS65_LH_IVX2 U15713 ( .A(n14335), .Z(n14337) );
  HS65_LH_NAND2X2 U15714 ( .A(n14622), .B(\u_DataPath/u_execute/A_inALU_i [20]), .Z(n14673) );
  HS65_LH_NAND4ABX3 U15715 ( .A(n14668), .B(n14337), .C(n14336), .D(n14673), 
        .Z(n14588) );
  HS65_LH_AOI22X1 U15716 ( .A(n15525), .B(n14589), .C(n13892), .D(n14588), .Z(
        n14342) );
  HS65_LH_CBI4I6X2 U15717 ( .A(n14349), .B(n17523), .C(n17248), .D(n33880), 
        .Z(n14341) );
  HS65_LH_NAND2AX4 U15718 ( .A(n14349), .B(n14035), .Z(n14339) );
  HS65_LH_OAI22X1 U15719 ( .A(n14339), .B(n17471), .C(n15398), .D(n14636), .Z(
        n14340) );
  HS65_LH_NOR4ABX2 U15720 ( .A(n14342), .B(n15098), .C(n14341), .D(n14340), 
        .Z(n14353) );
  HS65_LH_NOR2AX3 U15721 ( .A(n14344), .B(n14343), .Z(n14346) );
  HS65_LH_AOI21X2 U15722 ( .A(n14348), .B(n17600), .C(n33882), .Z(n14345) );
  HS65_LH_OAI21X2 U15723 ( .A(n14346), .B(n17467), .C(n14345), .Z(n14351) );
  HS65_LH_IVX2 U15724 ( .A(n14346), .Z(n14347) );
  HS65_LH_OAI22X1 U15725 ( .A(n14348), .B(n17468), .C(n17467), .D(n14347), .Z(
        n14350) );
  HS65_LH_AOI21X2 U15726 ( .A(n14349), .B(n14035), .C(n15251), .Z(n15213) );
  HS65_LH_MUXI21X2 U15727 ( .D0(n14351), .D1(n14350), .S0(n15213), .Z(n14352)
         );
  HS65_LH_NAND3X2 U15728 ( .A(n14354), .B(n14353), .C(n14352), .Z(n14355) );
  HS65_LH_AOI22X1 U15729 ( .A(n14358), .B(n17515), .C(n13892), .D(n14589), .Z(
        n14360) );
  HS65_LH_OAI211X1 U15730 ( .A(n14361), .B(n15080), .C(n14360), .D(n14359), 
        .Z(n14378) );
  HS65_LH_IVX2 U15731 ( .A(n14491), .Z(n14584) );
  HS65_LH_IVX2 U15732 ( .A(n15409), .Z(n15102) );
  HS65_LH_AOI22X1 U15733 ( .A(n15497), .B(n14486), .C(n15102), .D(n14587), .Z(
        n14364) );
  HS65_LH_AOI22X1 U15734 ( .A(n15126), .B(n14362), .C(n15499), .D(n14489), .Z(
        n14363) );
  HS65_LH_OAI211X1 U15735 ( .A(n14584), .B(n15417), .C(n14364), .D(n14363), 
        .Z(n14377) );
  HS65_LH_NOR2X2 U15736 ( .A(n14626), .B(n17249), .Z(n14663) );
  HS65_LH_NAND2X2 U15737 ( .A(n14622), .B(\u_DataPath/u_execute/A_inALU_i [12]), .Z(n14617) );
  HS65_LH_NAND4ABX3 U15738 ( .A(n14367), .B(n14663), .C(n14366), .D(n14617), 
        .Z(n14590) );
  HS65_LH_AOI22X1 U15739 ( .A(n15525), .B(n14590), .C(n15517), .D(n14588), .Z(
        n14376) );
  HS65_LH_NOR2AX3 U15740 ( .A(n14368), .B(n14441), .Z(n14370) );
  HS65_LH_AOI21X2 U15741 ( .A(n14372), .B(n17600), .C(n33882), .Z(n14369) );
  HS65_LH_OAI21X2 U15742 ( .A(n14370), .B(n17467), .C(n14369), .Z(n14374) );
  HS65_LH_IVX2 U15743 ( .A(n14370), .Z(n14371) );
  HS65_LH_OAI22X1 U15744 ( .A(n14372), .B(n17468), .C(n17467), .D(n14371), .Z(
        n14373) );
  HS65_LH_NOR2X2 U15745 ( .A(n15306), .B(n15262), .Z(n15193) );
  HS65_LH_MUXI21X2 U15746 ( .D0(n14374), .D1(n14373), .S0(n15193), .Z(n14375)
         );
  HS65_LH_NAND4ABX3 U15747 ( .A(n14378), .B(n14377), .C(n14376), .D(n14375), 
        .Z(n15554) );
  HS65_LH_AOI22X1 U15748 ( .A(n15331), .B(n14486), .C(n15075), .D(n14588), .Z(
        n14384) );
  HS65_LH_OAI21X2 U15749 ( .A(n14037), .B(n14382), .C(n14384), .Z(n14426) );
  HS65_LH_NOR2AX3 U15750 ( .A(n14383), .B(n15116), .Z(n14401) );
  HS65_LH_AOI21X2 U15751 ( .A(n14388), .B(n14386), .C(n15274), .Z(n14397) );
  HS65_LH_IVX2 U15752 ( .A(n14397), .Z(n15205) );
  HS65_LH_OAI21X2 U15753 ( .A(n15205), .B(n14401), .C(n17591), .Z(n14400) );
  HS65_LH_AOI21X2 U15754 ( .A(n14398), .B(n14397), .C(n17468), .Z(n14396) );
  HS65_LH_NAND2X2 U15755 ( .A(n6651), .B(n38579), .Z(n14952) );
  HS65_LH_NOR2X2 U15756 ( .A(n14952), .B(n15245), .Z(n14698) );
  HS65_LH_IVX2 U15757 ( .A(n14384), .Z(n14385) );
  HS65_LH_AOI211X1 U15758 ( .A(n15329), .B(n14487), .C(n14698), .D(n14385), 
        .Z(n14424) );
  HS65_LH_AOI22X1 U15759 ( .A(n15102), .B(n14489), .C(n15100), .D(n14587), .Z(
        n14394) );
  HS65_LH_IVX2 U15760 ( .A(n15417), .Z(n15133) );
  HS65_LH_AOI22X1 U15761 ( .A(n15405), .B(n14491), .C(n15133), .D(n14490), .Z(
        n14392) );
  HS65_LH_AOI21X2 U15762 ( .A(n17607), .B(n14633), .C(n14386), .Z(n14387) );
  HS65_LH_AOI22X1 U15763 ( .A(n14388), .B(n17515), .C(n17314), .D(n14387), .Z(
        n14391) );
  HS65_LH_IVX2 U15764 ( .A(n15098), .Z(n15030) );
  HS65_LH_OAI22X1 U15765 ( .A(n14397), .B(n17638), .C(n14389), .D(n15026), .Z(
        n14390) );
  HS65_LH_NOR4ABX2 U15766 ( .A(n14392), .B(n14391), .C(n15030), .D(n14390), 
        .Z(n14393) );
  HS65_LH_OAI211X1 U15767 ( .A(n14424), .B(n15120), .C(n14394), .D(n14393), 
        .Z(n14395) );
  HS65_LH_CBI4I6X2 U15768 ( .A(n14398), .B(n14397), .C(n14396), .D(n14395), 
        .Z(n14399) );
  HS65_LH_CBI4I1X3 U15769 ( .A(n14401), .B(n15205), .C(n14400), .D(n14399), 
        .Z(n14402) );
  HS65_LH_FA1X4 U15770 ( .A0(n6650), .B0(\u_DataPath/u_idexreg/N28 ), .CI(
        n14403), .CO(n14908), .S0(n14404) );
  HS65_LH_NOR2AX3 U15771 ( .A(n14407), .B(n14406), .Z(n14420) );
  HS65_LH_CNIVX3 U15772 ( .A(n15495), .Z(n15715) );
  HS65_LH_AOI22X1 U15773 ( .A(n17591), .B(n14420), .C(n17590), .D(n14419), .Z(
        n14428) );
  HS65_LH_MUXI21X2 U15774 ( .D0(n6651), .D1(n14037), .S0(n15246), .Z(n15196)
         );
  HS65_LH_AOI22X1 U15775 ( .A(n15497), .B(n14589), .C(n15517), .D(n14590), .Z(
        n14418) );
  HS65_LH_OAI211X1 U15776 ( .A(n17606), .B(n15246), .C(n17314), .D(n6651), .Z(
        n14417) );
  HS65_LH_NAND2X2 U15777 ( .A(n14622), .B(n14030), .Z(n14614) );
  HS65_LH_NOR2X2 U15778 ( .A(n14626), .B(n17253), .Z(n14618) );
  HS65_LH_NOR4ABX2 U15779 ( .A(n14411), .B(n14614), .C(n14410), .D(n14618), 
        .Z(n14593) );
  HS65_LH_NAND2X2 U15781 ( .A(n15246), .B(n14218), .Z(n14413) );
  HS65_LH_NAND2X2 U15782 ( .A(n15044), .B(n14029), .Z(n14615) );
  HS65_LH_NOR2X2 U15783 ( .A(n14621), .B(n14921), .Z(n14619) );
  HS65_LH_NOR4ABX2 U15784 ( .A(n14413), .B(n14615), .C(n14412), .D(n14619), 
        .Z(n14414) );
  HS65_LH_IVX2 U15785 ( .A(n15525), .Z(n15141) );
  HS65_LH_OAI22X1 U15786 ( .A(n14593), .B(n29699), .C(n14414), .D(n15141), .Z(
        n14416) );
  HS65_LH_OAI22X1 U15787 ( .A(n14495), .B(n15026), .C(n33880), .D(n15507), .Z(
        n14415) );
  HS65_LH_NOR4ABX2 U15788 ( .A(n14418), .B(n14417), .C(n14416), .D(n14415), 
        .Z(n14423) );
  HS65_LH_IVX2 U15789 ( .A(n14419), .Z(n14421) );
  HS65_LH_NOR2X2 U15790 ( .A(n14420), .B(n17467), .Z(n15070) );
  HS65_LH_CBI4I1X3 U15791 ( .A(n17590), .B(n14421), .C(n15070), .D(n15196), 
        .Z(n14422) );
  HS65_LH_OAI211X1 U15792 ( .A(n14424), .B(n15080), .C(n14423), .D(n14422), 
        .Z(n14425) );
  HS65_LH_AOI21X2 U15793 ( .A(n15126), .B(n14426), .C(n14425), .Z(n14427) );
  HS65_LH_MUXI21X2 U15794 ( .D0(n8855), .D1(n8860), .S0(n6650), .Z(n14429) );
  HS65_LH_IVX2 U15795 ( .A(n15076), .Z(n14898) );
  HS65_LH_NAND2X2 U15796 ( .A(n15039), .B(n15074), .Z(n14444) );
  HS65_LH_OA112X4 U15797 ( .A(n14547), .B(n14898), .C(n14444), .D(n14952), .Z(
        n14474) );
  HS65_LH_AOI22X1 U15798 ( .A(n15499), .B(n15101), .C(n15497), .D(n15073), .Z(
        n14435) );
  HS65_LH_CBI4I1X3 U15799 ( .A(n17606), .B(n14433), .C(n14033), .D(n17515), 
        .Z(n14430) );
  HS65_LH_OAI21X2 U15800 ( .A(n14431), .B(n29699), .C(n14430), .Z(n14432) );
  HS65_LH_AOI31X2 U15801 ( .A(n14033), .B(n17314), .C(n14433), .D(n14432), .Z(
        n14434) );
  HS65_LH_OAI21X2 U15802 ( .A(n14439), .B(n17468), .C(n17638), .Z(n14437) );
  HS65_LH_AOI21X2 U15803 ( .A(n17591), .B(n14438), .C(n14437), .Z(n14443) );
  HS65_LH_IVX2 U15804 ( .A(n14438), .Z(n14440) );
  HS65_LH_AOI22X1 U15805 ( .A(n17601), .B(n14440), .C(n17590), .D(n14439), .Z(
        n14442) );
  HS65_LH_IVX2 U15806 ( .A(n15298), .Z(n15302) );
  HS65_LH_NOR2X2 U15807 ( .A(n15302), .B(n14441), .Z(n15192) );
  HS65_LH_MUXI21X2 U15808 ( .D0(n14443), .D1(n14442), .S0(n15192), .Z(n14449)
         );
  HS65_LH_AO22X4 U15809 ( .A(n15331), .B(n15131), .C(n15329), .D(n15132), .Z(
        n14465) );
  HS65_LH_OAI21X2 U15810 ( .A(n14895), .B(n14547), .C(n14444), .Z(n14464) );
  HS65_LH_AOI22X1 U15811 ( .A(n14930), .B(n14465), .C(n15126), .D(n14464), .Z(
        n14448) );
  HS65_LH_NOR2X2 U15812 ( .A(n15328), .B(n17252), .Z(n14546) );
  HS65_LH_NAND2X2 U15813 ( .A(n15044), .B(n14032), .Z(n14803) );
  HS65_LH_NAND4ABX3 U15814 ( .A(n14446), .B(n14546), .C(n14445), .D(n14803), 
        .Z(n15130) );
  HS65_LH_AOI22X1 U15815 ( .A(n15525), .B(n15130), .C(n15517), .D(n15129), .Z(
        n14447) );
  HS65_LH_NAND4ABX3 U15816 ( .A(n14436), .B(n14449), .C(n33254), .D(n14447), 
        .Z(n15544) );
  HS65_LH_IVX2 U15817 ( .A(n15103), .Z(n14455) );
  HS65_LH_NAND2X2 U15818 ( .A(n15044), .B(n14642), .Z(n14561) );
  HS65_LH_NAND2X2 U15819 ( .A(n14622), .B(n14752), .Z(n14554) );
  HS65_LH_NOR4ABX2 U15820 ( .A(n14561), .B(n14554), .C(n14454), .D(n14453), 
        .Z(n14529) );
  HS65_LH_OAI22X1 U15821 ( .A(n14455), .B(n14827), .C(n14529), .D(n15026), .Z(
        n14480) );
  HS65_LH_OAI21X2 U15822 ( .A(n14456), .B(n15291), .C(n14760), .Z(n14457) );
  HS65_LH_AOI22X1 U15823 ( .A(n32629), .B(n14457), .C(n32748), .D(n14458), .Z(
        n14463) );
  HS65_LH_IVX2 U15824 ( .A(n14457), .Z(n14460) );
  HS65_LH_OAI21X2 U15825 ( .A(n14458), .B(n17468), .C(n17638), .Z(n14459) );
  HS65_LH_AOI21X2 U15826 ( .A(n17591), .B(n14460), .C(n14459), .Z(n14462) );
  HS65_LH_OAI21X2 U15827 ( .A(n14461), .B(n14553), .C(n14516), .Z(n15227) );
  HS65_LH_MUXI21X2 U15828 ( .D0(n14463), .D1(n14462), .S0(n15227), .Z(n14479)
         );
  HS65_LH_AOI22X1 U15829 ( .A(n29624), .B(n14465), .C(n14900), .D(n14464), .Z(
        n14478) );
  HS65_LH_NOR2X2 U15830 ( .A(n14621), .B(n15032), .Z(n14551) );
  HS65_LH_NAND2X2 U15831 ( .A(n15044), .B(n14035), .Z(n14556) );
  HS65_LH_NAND4ABX3 U15832 ( .A(n14551), .B(n14467), .C(n14556), .D(n14466), 
        .Z(n15110) );
  HS65_LH_OAI211X1 U15833 ( .A(n33045), .B(n14553), .C(n17314), .D(n14468), 
        .Z(n14469) );
  HS65_LH_OAI211X1 U15834 ( .A(n33880), .B(n14470), .C(n15098), .D(n14469), 
        .Z(n14476) );
  HS65_LH_NOR2X2 U15835 ( .A(n14621), .B(n14709), .Z(n14560) );
  HS65_LH_NOR2X2 U15836 ( .A(n14626), .B(n14633), .Z(n14552) );
  HS65_LH_OR4X4 U15837 ( .A(n14560), .B(n14552), .C(n14472), .D(n14471), .Z(
        n14878) );
  HS65_LH_AOI22X1 U15838 ( .A(n15133), .B(n14878), .C(n15100), .D(n15101), .Z(
        n14473) );
  HS65_LH_OAI21X2 U15839 ( .A(n14474), .B(n15120), .C(n14473), .Z(n14475) );
  HS65_LH_AOI211X1 U15840 ( .A(n15102), .B(n15110), .C(n14476), .D(n14475), 
        .Z(n14477) );
  HS65_LH_NAND4ABX3 U15841 ( .A(n14480), .B(n14479), .C(n14478), .D(n32152), 
        .Z(n15573) );
  HS65_LH_AOI22X1 U15842 ( .A(n15331), .B(n14487), .C(n15075), .D(n14486), .Z(
        n14488) );
  HS65_LH_OAI21X2 U15843 ( .A(n14897), .B(n15398), .C(n14488), .Z(n14580) );
  HS65_LH_IVX2 U15844 ( .A(n15120), .Z(n14899) );
  HS65_LH_NAND2X2 U15845 ( .A(n14488), .B(n14952), .Z(n14581) );
  HS65_LH_AOI22X1 U15846 ( .A(n14900), .B(n14580), .C(n14899), .D(n14581), .Z(
        n14508) );
  HS65_LH_AOI22X1 U15847 ( .A(n15102), .B(n14490), .C(n15405), .D(n14489), .Z(
        n14499) );
  HS65_LH_AOI22X1 U15848 ( .A(n15133), .B(n15404), .C(n15100), .D(n14491), .Z(
        n14498) );
  HS65_LH_AOI22X1 U15849 ( .A(n17314), .B(n14492), .C(n14642), .D(n17515), .Z(
        n14493) );
  HS65_LH_CBI4I1X3 U15850 ( .A(n14494), .B(n17523), .C(n14493), .D(n15098), 
        .Z(n14497) );
  HS65_LH_OAI22X1 U15851 ( .A(n14495), .B(n14710), .C(n15410), .D(n15026), .Z(
        n14496) );
  HS65_LH_OAI21X2 U15852 ( .A(n14891), .B(n14888), .C(n14889), .Z(n14503) );
  HS65_LH_OAI22X1 U15853 ( .A(n17467), .B(n14503), .C(n32759), .D(n14502), .Z(
        n14506) );
  HS65_LH_NAND2X2 U15854 ( .A(n15277), .B(n14501), .Z(n15215) );
  HS65_LH_AOI22X1 U15855 ( .A(n32629), .B(n14503), .C(n17590), .D(n14502), .Z(
        n14504) );
  HS65_LH_NAND3X2 U15856 ( .A(n14504), .B(n17638), .C(n15215), .Z(n14505) );
  HS65_LH_OAI21X2 U15857 ( .A(n14506), .B(n15215), .C(n14505), .Z(n14507) );
  HS65_LH_NAND2X2 U15858 ( .A(n14875), .B(n17914), .Z(n14874) );
  HS65_LH_CNIVX3 U15859 ( .A(\u_DataPath/pc_4_to_ex_i [29]), .Z(n14655) );
  HS65_LH_NOR2X2 U15860 ( .A(n14874), .B(n40650), .Z(n14654) );
  HS65_LH_NAND2X2 U15861 ( .A(n14654), .B(n17549), .Z(n15388) );
  HS65_LH_MUX21I1X3 U15862 ( .D0(n32121), .D1(n29692), .S0(n17528), .Z(n15394)
         );
  HS65_LH_IVX2 U15865 ( .A(n33227), .Z(n15349) );
  HS65_LH_NOR2X2 U15866 ( .A(n29635), .B(n40560), .Z(n15311) );
  HS65_LH_NOR2X2 U15867 ( .A(n15349), .B(n15311), .Z(n15200) );
  HS65_LH_MUX21I1X3 U15868 ( .D0(n29692), .D1(n32104), .S0(n17608), .Z(n14522)
         );
  HS65_LH_IVX2 U15869 ( .A(n14522), .Z(n14685) );
  HS65_LH_NOR2X2 U15870 ( .A(n14521), .B(n14685), .Z(n14658) );
  HS65_LH_MUX21I1X3 U15871 ( .D0(n32381), .D1(n29693), .S0(n17528), .Z(n14849)
         );
  HS65_LH_NOR2X2 U15872 ( .A(n14852), .B(n14849), .Z(n14864) );
  HS65_LH_NOR2X2 U15873 ( .A(n14658), .B(n14864), .Z(n15351) );
  HS65_LH_NOR2X2 U15874 ( .A(n14515), .B(n15233), .Z(n14518) );
  HS65_LH_OAI21X2 U15875 ( .A(n14843), .B(n14517), .C(n14516), .Z(n15290) );
  HS65_LH_OAI21X2 U15876 ( .A(n14518), .B(n15290), .C(n15235), .Z(n14862) );
  HS65_LH_NAND2X2 U15877 ( .A(n15351), .B(n14862), .Z(n15390) );
  HS65_LH_NOR2X2 U15878 ( .A(n14031), .B(n14522), .Z(n14657) );
  HS65_LH_IVX2 U15879 ( .A(n14849), .Z(n14853) );
  HS65_LH_NOR2X2 U15880 ( .A(n14850), .B(n14853), .Z(n14863) );
  HS65_LH_NOR2X2 U15881 ( .A(n14657), .B(n14863), .Z(n15370) );
  HS65_LH_NOR2X2 U15882 ( .A(n14658), .B(n15370), .Z(n15296) );
  HS65_LH_NOR2AX3 U15883 ( .A(n15390), .B(n15296), .Z(n14524) );
  HS65_LH_PAOI2X1 U15884 ( .A(n14520), .B(n14519), .P(n14843), .Z(n14861) );
  HS65_LH_PAOI2X1 U15885 ( .A(n14850), .B(n14849), .P(n14861), .Z(n14661) );
  HS65_LH_PAOI2X1 U15886 ( .A(n14522), .B(n14521), .P(n14661), .Z(n15395) );
  HS65_LH_IVX2 U15889 ( .A(n40544), .Z(n14540) );
  HS65_LH_IVX2 U15890 ( .A(n14524), .Z(n14525) );
  HS65_LH_AOI22X1 U15891 ( .A(n32629), .B(n14525), .C(n32748), .D(n15395), .Z(
        n14539) );
  HS65_LH_NAND2X2 U15892 ( .A(n14622), .B(n14031), .Z(n14548) );
  HS65_LH_NOR2X2 U15893 ( .A(n14626), .B(n14843), .Z(n14555) );
  HS65_LH_NOR4ABX2 U15894 ( .A(n14527), .B(n14548), .C(n14555), .D(n14526), 
        .Z(n14528) );
  HS65_LH_OAI22X1 U15895 ( .A(n14529), .B(n15417), .C(n14528), .D(n15026), .Z(
        n14536) );
  HS65_LH_AOI22X1 U15896 ( .A(n15405), .B(n15110), .C(n15102), .D(n14878), .Z(
        n14533) );
  HS65_LH_NAND2X2 U15897 ( .A(n15039), .B(n14900), .Z(n15399) );
  HS65_LH_CNIVX3 U15898 ( .A(n15411), .Z(n15342) );
  HS65_LH_CBI4I1X3 U15899 ( .A(n17587), .B(n15394), .C(n40560), .D(n17515), 
        .Z(n14530) );
  HS65_LH_OAI211X1 U15900 ( .A(n14895), .B(n15399), .C(n15098), .D(n14530), 
        .Z(n14531) );
  HS65_LH_AOI31X2 U15901 ( .A(n40560), .B(n35562), .C(n15394), .D(n14531), .Z(
        n14532) );
  HS65_LH_OAI211X1 U15902 ( .A(n14534), .B(n15120), .C(n14533), .D(n14532), 
        .Z(n14535) );
  HS65_LH_NAND2X2 U15903 ( .A(n14218), .B(n14030), .Z(n14927) );
  HS65_LH_NAND2X2 U15904 ( .A(n15325), .B(n14029), .Z(n14914) );
  HS65_LH_NOR2X2 U15905 ( .A(n15328), .B(n17254), .Z(n15058) );
  HS65_LH_NOR2X2 U15906 ( .A(n14626), .B(n14730), .Z(n15083) );
  HS65_LH_NOR4ABX2 U15907 ( .A(n14927), .B(n14914), .C(n15058), .D(n15083), 
        .Z(n15006) );
  HS65_LH_NAND2X2 U15908 ( .A(n15195), .B(n15335), .Z(n15327) );
  HS65_LH_IVX2 U15909 ( .A(n15327), .Z(n14947) );
  HS65_LH_NOR2X2 U15910 ( .A(n14226), .B(n14921), .Z(n14916) );
  HS65_LH_NOR2X2 U15911 ( .A(n15328), .B(n15507), .Z(n15084) );
  HS65_LH_AOI211X1 U15912 ( .A(n15502), .B(n15044), .C(n14916), .D(n15084), 
        .Z(n14544) );
  HS65_LH_OAI21X2 U15913 ( .A(n15508), .B(n15062), .C(n14544), .Z(n15003) );
  HS65_LH_MUXI21X2 U15914 ( .D0(n14947), .D1(n15003), .S0(n15245), .Z(n14924)
         );
  HS65_LH_NOR2X2 U15915 ( .A(n14226), .B(n17250), .Z(n14557) );
  HS65_LH_NAND2X2 U15916 ( .A(n15325), .B(n14033), .Z(n14926) );
  HS65_LH_NAND2X2 U15917 ( .A(n15044), .B(n14545), .Z(n15060) );
  HS65_LH_NAND4ABX3 U15918 ( .A(n14557), .B(n14546), .C(n14926), .D(n15060), 
        .Z(n14996) );
  HS65_LH_IVX2 U15919 ( .A(n14996), .Z(n14828) );
  HS65_LH_OAI222X2 U15920 ( .A(n14547), .B(n15006), .C(n14924), .D(n14037), 
        .E(n14625), .F(n14828), .Z(n14869) );
  HS65_LH_NOR2X2 U15921 ( .A(n14626), .B(n10437), .Z(n14769) );
  HS65_LH_OAI21X2 U15922 ( .A(n14852), .B(n14226), .C(n14548), .Z(n14549) );
  HS65_LH_AOI211X1 U15923 ( .A(n40560), .B(n15325), .C(n14769), .D(n14549), 
        .Z(n14855) );
  HS65_LH_IVX2 U15924 ( .A(n14855), .Z(n14991) );
  HS65_LH_AOI21X2 U15925 ( .A(n15039), .B(n14991), .C(n14623), .Z(n14854) );
  HS65_LH_NOR2X2 U15926 ( .A(n14226), .B(n14550), .Z(n14806) );
  HS65_LH_NOR2X2 U15927 ( .A(n15508), .B(n15099), .Z(n14810) );
  HS65_LH_OR4X4 U15928 ( .A(n14552), .B(n14551), .C(n14806), .D(n14810), .Z(
        n14993) );
  HS65_LH_NOR2X2 U15929 ( .A(n14226), .B(n14817), .Z(n14816) );
  HS65_LH_NAND2X2 U15930 ( .A(n15325), .B(n14553), .Z(n14845) );
  HS65_LH_NAND4ABX3 U15931 ( .A(n14555), .B(n14816), .C(n14554), .D(n14845), 
        .Z(n14992) );
  HS65_LH_AOI22X1 U15932 ( .A(n13892), .B(n14993), .C(n15497), .D(n14992), .Z(
        n14567) );
  HS65_LH_NAND2X2 U15933 ( .A(n15325), .B(n14036), .Z(n14804) );
  HS65_LH_NAND4ABX3 U15934 ( .A(n14558), .B(n14557), .C(n14556), .D(n14804), 
        .Z(n15334) );
  HS65_LH_NAND2X2 U15935 ( .A(n15325), .B(n14559), .Z(n14814) );
  HS65_LH_NOR2X2 U15936 ( .A(n14226), .B(n15272), .Z(n14809) );
  HS65_LH_NOR4ABX2 U15937 ( .A(n14561), .B(n14814), .C(n14560), .D(n14809), 
        .Z(n14937) );
  HS65_LH_IVX2 U15938 ( .A(n15517), .Z(n15063) );
  HS65_LH_OAI22X1 U15939 ( .A(n14937), .B(n15063), .C(n14855), .D(n14636), .Z(
        n14565) );
  HS65_LH_OAI21X2 U15940 ( .A(n33505), .B(n17250), .C(n17523), .Z(n14562) );
  HS65_LH_OAI21X2 U15941 ( .A(\u_DataPath/u_execute/A_inALU_i [12]), .B(n15237), .C(n14562), .Z(n14563) );
  HS65_LH_OAI31X1 U15942 ( .A(n17471), .B(n15252), .C(n17250), .D(n14563), .Z(
        n14564) );
  HS65_LH_AOI211X1 U15943 ( .A(n15525), .B(n15334), .C(n14565), .D(n14564), 
        .Z(n14566) );
  HS65_LH_OAI211X1 U15944 ( .A(n14854), .B(n15080), .C(n14567), .D(n14566), 
        .Z(n14575) );
  HS65_LH_OAI21X2 U15945 ( .A(n14570), .B(n17468), .C(n17638), .Z(n14568) );
  HS65_LH_AOI21X2 U15946 ( .A(n17591), .B(n14569), .C(n14568), .Z(n14573) );
  HS65_LH_IVX2 U15947 ( .A(n14569), .Z(n14571) );
  HS65_LH_AOI22X1 U15948 ( .A(n17591), .B(n14571), .C(n17600), .D(n14570), .Z(
        n14572) );
  HS65_LH_MUXI21X2 U15949 ( .D0(n17250), .D1(
        \u_DataPath/u_execute/A_inALU_i [12]), .S0(n15252), .Z(n15189) );
  HS65_LH_MUXI21X2 U15950 ( .D0(n14573), .D1(n14572), .S0(n15189), .Z(n14574)
         );
  HS65_LH_MUXI21X2 U15951 ( .D0(n17254), .D1(n14583), .S0(n14586), .Z(n15206)
         );
  HS65_LH_PAOI2X1 U15952 ( .A(n14913), .B(n14921), .P(n14919), .Z(n15144) );
  HS65_LH_NOR2X2 U15953 ( .A(n15145), .B(n15144), .Z(n14579) );
  HS65_LH_OAI21X2 U15954 ( .A(n14579), .B(n14578), .C(n15146), .Z(n14603) );
  HS65_LH_AOI21X2 U15955 ( .A(n15206), .B(n14603), .C(n33640), .Z(n14602) );
  HS65_LH_OAI21X2 U15956 ( .A(n14600), .B(n15206), .C(n17600), .Z(n14599) );
  HS65_LH_AOI22X1 U15957 ( .A(n15128), .B(n14581), .C(n15126), .D(n14580), .Z(
        n14597) );
  HS65_LH_IVX2 U15958 ( .A(n15206), .Z(n14582) );
  HS65_LH_AOI22X1 U15959 ( .A(n14583), .B(n17515), .C(n33882), .D(n14582), .Z(
        n14596) );
  HS65_LH_OAI21X2 U15960 ( .A(n17606), .B(n14583), .C(n17314), .Z(n14585) );
  HS65_LH_OAI22X1 U15961 ( .A(n14586), .B(n14585), .C(n14584), .D(n15026), .Z(
        n14595) );
  HS65_LH_AOI22X1 U15962 ( .A(n15497), .B(n14588), .C(n15133), .D(n14587), .Z(
        n14592) );
  HS65_LH_AOI22X1 U15963 ( .A(n13892), .B(n14590), .C(n15517), .D(n14589), .Z(
        n14591) );
  HS65_LH_OAI211X1 U15964 ( .A(n14593), .B(n15141), .C(n14592), .D(n14591), 
        .Z(n14594) );
  HS65_LH_NOR4ABX2 U15965 ( .A(n14597), .B(n14596), .C(n14595), .D(n14594), 
        .Z(n14598) );
  HS65_LH_CBI4I1X3 U15966 ( .A(n15206), .B(n14600), .C(n14599), .D(n14598), 
        .Z(n14601) );
  HS65_LH_NOR2AX3 U15967 ( .A(n15236), .B(n14608), .Z(n14652) );
  HS65_LH_IVX2 U15968 ( .A(n14612), .Z(n14609) );
  HS65_LH_OAI22X1 U15969 ( .A(n14609), .B(n17467), .C(n14610), .D(n17468), .Z(
        n14651) );
  HS65_LH_IVX2 U15970 ( .A(n14652), .Z(n15187) );
  HS65_LH_AOI21X2 U15971 ( .A(n14610), .B(n17600), .C(n33882), .Z(n14611) );
  HS65_LH_OAI21X2 U15972 ( .A(n17467), .B(n14612), .C(n14611), .Z(n14650) );
  HS65_LH_NOR2X2 U15973 ( .A(n14226), .B(n17256), .Z(n14727) );
  HS65_LH_NOR2X2 U15974 ( .A(n15508), .B(n17254), .Z(n14725) );
  HS65_LH_NAND4ABX3 U15975 ( .A(n14727), .B(n14725), .C(n14615), .D(n14614), 
        .Z(n14779) );
  HS65_LH_NOR2X2 U15976 ( .A(n15508), .B(n17252), .Z(n14726) );
  HS65_LH_NAND2X2 U15977 ( .A(n14231), .B(n14032), .Z(n14639) );
  HS65_LH_NAND4ABX3 U15978 ( .A(n14726), .B(n14618), .C(n14617), .D(n14639), 
        .Z(n15025) );
  HS65_LH_NOR2X2 U15979 ( .A(n14226), .B(n14730), .Z(n14724) );
  HS65_LH_AOI211X1 U15980 ( .A(n15324), .B(n15044), .C(n14724), .D(n14619), 
        .Z(n14620) );
  HS65_LH_OAI21X2 U15981 ( .A(n15508), .B(n15507), .C(n14620), .Z(n15036) );
  HS65_LH_NAND3AX3 U15982 ( .A(n15341), .B(n15195), .C(n15502), .Z(n15509) );
  HS65_LH_OAI21X2 U15983 ( .A(n14621), .B(n15337), .C(n15509), .Z(n15498) );
  HS65_LH_MX41X4 U15984 ( .D0(n14779), .S0(n15331), .D1(n15025), .S1(n15039), 
        .D2(n15036), .S2(n15329), .D3(n15498), .S3(n15333), .Z(n14676) );
  HS65_LH_NAND2X2 U15985 ( .A(n14622), .B(n40560), .Z(n15401) );
  HS65_LH_NAND2X2 U15986 ( .A(n14231), .B(n14031), .Z(n14681) );
  HS65_LH_OAI211X1 U15987 ( .A(n10437), .B(n15508), .C(n15401), .D(n14681), 
        .Z(n15037) );
  HS65_LH_AOI21X2 U15988 ( .A(n15044), .B(n38579), .C(n15037), .Z(n14699) );
  HS65_LH_IVX2 U15989 ( .A(n14623), .Z(n14624) );
  HS65_LH_OAI21X2 U15990 ( .A(n14699), .B(n14625), .C(n14624), .Z(n14675) );
  HS65_LH_AOI22X1 U15991 ( .A(n14930), .B(n14676), .C(n15128), .D(n14675), .Z(
        n14648) );
  HS65_LH_NOR2X2 U15992 ( .A(n14626), .B(n14852), .Z(n15402) );
  HS65_LH_NAND2X2 U15993 ( .A(n14643), .B(n14627), .Z(n14680) );
  HS65_LH_NAND2X2 U15994 ( .A(n14231), .B(n14752), .Z(n14670) );
  HS65_LH_NAND4ABX3 U15995 ( .A(n14628), .B(n15402), .C(n14680), .D(n14670), 
        .Z(n15038) );
  HS65_LH_NOR3X1 U15996 ( .A(n14632), .B(n17255), .C(n17471), .Z(n14629) );
  HS65_LH_CBI4I6X2 U15997 ( .A(n14032), .B(n17587), .C(n17515), .D(n14629), 
        .Z(n14630) );
  HS65_LH_AOI21X2 U15998 ( .A(n14632), .B(n32851), .C(n14630), .Z(n14638) );
  HS65_LH_NOR2X2 U15999 ( .A(n15508), .B(n14633), .Z(n14672) );
  HS65_LH_NAND2X2 U16000 ( .A(n14218), .B(n15018), .Z(n14666) );
  HS65_LH_NAND4ABX3 U16001 ( .A(n14635), .B(n14672), .C(n14634), .D(n14666), 
        .Z(n15040) );
  HS65_LH_IVX2 U16002 ( .A(n15040), .Z(n14783) );
  HS65_LH_IVX2 U16003 ( .A(n15037), .Z(n14706) );
  HS65_LH_OAI22X1 U16004 ( .A(n14783), .B(n29699), .C(n14706), .D(n14636), .Z(
        n14637) );
  HS65_LH_AOI211X1 U16005 ( .A(n15497), .B(n15038), .C(n14638), .D(n14637), 
        .Z(n14647) );
  HS65_LH_NAND2X2 U16006 ( .A(n15325), .B(n14035), .Z(n14665) );
  HS65_LH_NAND4ABX3 U16007 ( .A(n14641), .B(n14640), .C(n14639), .D(n14665), 
        .Z(n15496) );
  HS65_LH_NAND2X2 U16008 ( .A(n14643), .B(n14642), .Z(n14669) );
  HS65_LH_NAND2X2 U16009 ( .A(n14218), .B(n15268), .Z(n14674) );
  HS65_LH_NAND4ABX3 U16010 ( .A(n14645), .B(n14644), .C(n14669), .D(n14674), 
        .Z(n15041) );
  HS65_LH_AOI22X1 U16011 ( .A(n15525), .B(n15496), .C(n15517), .D(n15041), .Z(
        n14646) );
  HS65_LH_NAND3X2 U16012 ( .A(n14648), .B(n14647), .C(n14646), .Z(n14649) );
  HS65_LH_NOR2X2 U16013 ( .A(n14658), .B(n14657), .Z(n14694) );
  HS65_LH_IVX2 U16014 ( .A(n14864), .Z(n14659) );
  HS65_LH_AOI21X2 U16015 ( .A(n14862), .B(n14659), .C(n14863), .Z(n14662) );
  HS65_LH_AO12X4 U16016 ( .A(n17591), .B(n14662), .C(n33882), .Z(n14660) );
  HS65_LH_OAI22X1 U16018 ( .A(n14662), .B(n33067), .C(n32759), .D(n14661), .Z(
        n14691) );
  HS65_LH_NOR4ABX2 U16019 ( .A(n14666), .B(n14665), .C(n14664), .D(n14663), 
        .Z(n15027) );
  HS65_LH_OAI22X1 U16020 ( .A(n14706), .B(n15399), .C(n15027), .D(n14827), .Z(
        n14689) );
  HS65_LH_NOR4ABX2 U16021 ( .A(n14670), .B(n14669), .C(n14668), .D(n14667), 
        .Z(n14768) );
  HS65_LH_NOR4ABX2 U16022 ( .A(n14674), .B(n14673), .C(n14672), .D(n14671), 
        .Z(n14767) );
  HS65_LH_OAI22X1 U16023 ( .A(n14768), .B(n15417), .C(n14767), .D(n15409), .Z(
        n14688) );
  HS65_LH_AOI22X1 U16024 ( .A(n29624), .B(n14676), .C(n14899), .D(n14675), .Z(
        n14687) );
  HS65_LH_IVX2 U16025 ( .A(n14677), .Z(n14679) );
  HS65_LH_NOR4ABX2 U16026 ( .A(n14681), .B(n14680), .C(n14679), .D(n14678), 
        .Z(n14683) );
  HS65_LH_CBI4I1X3 U16027 ( .A(n17587), .B(n14685), .C(n14031), .D(n17515), 
        .Z(n14682) );
  HS65_LH_OAI211X1 U16028 ( .A(n14683), .B(n15026), .C(n15098), .D(n14682), 
        .Z(n14684) );
  HS65_LH_AOI31X2 U16029 ( .A(n14031), .B(n35562), .C(n14685), .D(n14684), .Z(
        n14686) );
  HS65_LH_NAND4ABX3 U16030 ( .A(n14689), .B(n14688), .C(n14687), .D(n14686), 
        .Z(n14690) );
  HS65_LH_AOI21X2 U16031 ( .A(n14691), .B(n14694), .C(n14690), .Z(n14692) );
  HS65_LH_AOI22X1 U16032 ( .A(n15331), .B(n15038), .C(n15075), .D(n15041), .Z(
        n14705) );
  HS65_LH_IVX2 U16033 ( .A(n14698), .Z(n14936) );
  HS65_LH_OAI211X1 U16034 ( .A(n14699), .B(n14897), .C(n14705), .D(n14936), 
        .Z(n14740) );
  HS65_LH_NOR2X2 U16035 ( .A(n14700), .B(n17467), .Z(n14887) );
  HS65_LH_NAND2X2 U16036 ( .A(n14701), .B(n14713), .Z(n14702) );
  HS65_LH_AOI22X1 U16037 ( .A(n14899), .B(n14740), .C(n14887), .D(n14702), .Z(
        n14719) );
  HS65_LH_IVX2 U16038 ( .A(n14713), .Z(n15203) );
  HS65_LH_IVX2 U16039 ( .A(n14704), .Z(n14703) );
  HS65_LH_OAI212X3 U16040 ( .A(n15203), .B(n14704), .C(n14713), .D(n14703), 
        .E(n17590), .Z(n14718) );
  HS65_LH_IVX2 U16041 ( .A(n14779), .Z(n15047) );
  HS65_LH_OAI22X1 U16042 ( .A(n15047), .B(n14827), .C(n14767), .D(n15026), .Z(
        n14717) );
  HS65_LH_OA12X4 U16043 ( .A(n14897), .B(n14706), .C(n14705), .Z(n14737) );
  HS65_LH_IVX2 U16044 ( .A(n14900), .Z(n15106) );
  HS65_LH_AOI22X1 U16045 ( .A(n15102), .B(n15025), .C(n15100), .D(n15036), .Z(
        n14715) );
  HS65_LH_OAI211X1 U16046 ( .A(n33045), .B(n15268), .C(n17314), .D(n14707), 
        .Z(n14708) );
  HS65_LH_OAI211X1 U16047 ( .A(n33880), .B(n14709), .C(n15098), .D(n14708), 
        .Z(n14712) );
  HS65_LH_IVX2 U16048 ( .A(n15498), .Z(n14786) );
  HS65_LH_OAI22X1 U16049 ( .A(n14786), .B(n14710), .C(n15027), .D(n15417), .Z(
        n14711) );
  HS65_LH_AOI211X1 U16050 ( .A(n33882), .B(n14713), .C(n14712), .D(n14711), 
        .Z(n14714) );
  HS65_LH_OAI211X1 U16051 ( .A(n14737), .B(n15106), .C(n14715), .D(n14714), 
        .Z(n14716) );
  HS65_LH_NOR4ABX2 U16052 ( .A(n14719), .B(n14718), .C(n14717), .D(n14716), 
        .Z(n15562) );
  HS65_LH_NAND4ABX3 U16053 ( .A(n14725), .B(n14724), .C(n14723), .D(n14722), 
        .Z(n15518) );
  HS65_LH_AOI22X1 U16054 ( .A(n15525), .B(n15518), .C(n15497), .D(n15040), .Z(
        n14746) );
  HS65_LH_NOR4X4 U16055 ( .A(n14729), .B(n14728), .C(n14727), .D(n14726), .Z(
        n14778) );
  HS65_LH_IVX2 U16056 ( .A(n14778), .Z(n15516) );
  HS65_LH_AOI22X1 U16057 ( .A(n15499), .B(n15036), .C(n13892), .D(n15516), .Z(
        n14745) );
  HS65_LH_CBI4I6X2 U16058 ( .A(n14731), .B(n17523), .C(n14730), .D(n33880), 
        .Z(n14732) );
  HS65_LH_AOI31X2 U16059 ( .A(n14734), .B(n35562), .C(n14733), .D(n14732), .Z(
        n14736) );
  HS65_LH_AOI22X1 U16060 ( .A(n15133), .B(n15498), .C(n15517), .D(n15496), .Z(
        n14735) );
  HS65_LH_OAI211X1 U16061 ( .A(n14737), .B(n15079), .C(n14736), .D(n14735), 
        .Z(n14744) );
  HS65_LH_AOI22X1 U16062 ( .A(n17591), .B(n15144), .C(n17590), .D(n14738), .Z(
        n14742) );
  HS65_LH_NOR2AX3 U16063 ( .A(n15143), .B(n15145), .Z(n15230) );
  HS65_LH_OAI22X1 U16064 ( .A(n14738), .B(n17468), .C(n15144), .D(n17467), .Z(
        n14739) );
  HS65_LH_AOI22X1 U16065 ( .A(n15128), .B(n14740), .C(n15230), .D(n14739), .Z(
        n14741) );
  HS65_LH_CBI4I1X3 U16066 ( .A(n14742), .B(n17638), .C(n15230), .D(n14741), 
        .Z(n14743) );
  HS65_LH_NOR4ABX2 U16067 ( .A(n14746), .B(n14745), .C(n14744), .D(n14743), 
        .Z(n15540) );
  HS65_LH_OAI21X2 U16068 ( .A(n14752), .B(n17587), .C(n17515), .Z(n14754) );
  HS65_LH_NAND3X2 U16069 ( .A(n14752), .B(n35562), .C(n14751), .Z(n14753) );
  HS65_LH_CBI4I1X3 U16070 ( .A(n14756), .B(n14755), .C(n14754), .D(n14753), 
        .Z(n14759) );
  HS65_LH_AOI22X1 U16071 ( .A(n15037), .B(n15331), .C(n15038), .D(n15075), .Z(
        n14770) );
  HS65_LH_IVX2 U16072 ( .A(n14770), .Z(n14776) );
  HS65_LH_AOI22X1 U16073 ( .A(n14900), .B(n14776), .C(n14879), .D(n15036), .Z(
        n14757) );
  HS65_LH_OAI21X2 U16074 ( .A(n15027), .B(n15409), .C(n14757), .Z(n14758) );
  HS65_LH_AOI211X1 U16075 ( .A(n15100), .B(n14779), .C(n14759), .D(n14758), 
        .Z(n14775) );
  HS65_LH_OAI21X2 U16076 ( .A(n15234), .B(n14831), .C(n14829), .Z(n14763) );
  HS65_LH_OAI22X1 U16077 ( .A(n14762), .B(n32759), .C(n17467), .D(n14763), .Z(
        n14766) );
  HS65_LH_NAND2X2 U16078 ( .A(n14761), .B(n14760), .Z(n15226) );
  HS65_LH_AOI22X1 U16079 ( .A(n32629), .B(n14763), .C(n32748), .D(n14762), .Z(
        n14764) );
  HS65_LH_NAND3X2 U16080 ( .A(n14764), .B(n17638), .C(n15226), .Z(n14765) );
  HS65_LH_OAI21X2 U16081 ( .A(n14766), .B(n15226), .C(n14765), .Z(n14774) );
  HS65_LH_OAI22X1 U16082 ( .A(n14768), .B(n15026), .C(n14767), .D(n15417), .Z(
        n14773) );
  HS65_LH_NAND2X2 U16083 ( .A(n14769), .B(n15069), .Z(n15528) );
  HS65_LH_NAND3X2 U16084 ( .A(n14770), .B(n14952), .C(n15528), .Z(n14780) );
  HS65_LH_AOI22X1 U16085 ( .A(n15405), .B(n15025), .C(n14899), .D(n14780), .Z(
        n14771) );
  HS65_LH_OAI211X1 U16086 ( .A(n14786), .B(n14824), .C(n14771), .D(n15098), 
        .Z(n14772) );
  HS65_LH_NOR4ABX2 U16087 ( .A(n14775), .B(n14774), .C(n14773), .D(n14772), 
        .Z(n15570) );
  HS65_LH_AOI22X1 U16088 ( .A(n15497), .B(n15041), .C(n15126), .D(n14776), .Z(
        n14777) );
  HS65_LH_OAI21X2 U16089 ( .A(n14778), .B(n15141), .C(n14777), .Z(n14798) );
  HS65_LH_AOI22X1 U16090 ( .A(n15133), .B(n15036), .C(n15499), .D(n14779), .Z(
        n14782) );
  HS65_LH_AOI22X1 U16091 ( .A(n15128), .B(n14780), .C(n13892), .D(n15496), .Z(
        n14781) );
  HS65_LH_OAI211X1 U16092 ( .A(n14783), .B(n15063), .C(n14782), .D(n14781), 
        .Z(n14797) );
  HS65_LH_PAOI2X1 U16093 ( .A(n14784), .B(n17256), .P(n17607), .Z(n14788) );
  HS65_LH_OAI22X1 U16094 ( .A(n14786), .B(n15409), .C(n17256), .D(n33505), .Z(
        n14787) );
  HS65_LH_AOI21X2 U16095 ( .A(n17260), .B(n15239), .C(n14790), .Z(n14792) );
  HS65_LH_OAI22X1 U16096 ( .A(n14791), .B(n17468), .C(n14792), .D(n17467), .Z(
        n14795) );
  HS65_LH_NAND2AX4 U16097 ( .A(n15301), .B(n15254), .Z(n15204) );
  HS65_LH_AOI22X1 U16098 ( .A(n17591), .B(n14792), .C(n17600), .D(n14791), .Z(
        n14793) );
  HS65_LH_NAND3X2 U16099 ( .A(n14793), .B(n17638), .C(n15204), .Z(n14794) );
  HS65_LH_OAI21X2 U16100 ( .A(n14795), .B(n15204), .C(n14794), .Z(n14796) );
  HS65_LH_NAND4ABX3 U16101 ( .A(n14798), .B(n14797), .C(n33501), .D(n14796), 
        .Z(n15550) );
  HS65_LH_NAND4ABX3 U16102 ( .A(n14806), .B(n14805), .C(n14804), .D(n14803), 
        .Z(n14995) );
  HS65_LH_NAND4ABX3 U16103 ( .A(n14810), .B(n14809), .C(n14808), .D(n14807), 
        .Z(n14982) );
  HS65_LH_AOI22X1 U16104 ( .A(n15133), .B(n14982), .C(n14879), .D(n15003), .Z(
        n14811) );
  HS65_LH_OAI21X2 U16105 ( .A(n15006), .B(n14999), .C(n14811), .Z(n14812) );
  HS65_LH_AOI21X2 U16106 ( .A(n15102), .B(n14995), .C(n14812), .Z(n14837) );
  HS65_LH_NAND4ABX3 U16107 ( .A(n14816), .B(n14815), .C(n14814), .D(n14813), 
        .Z(n14842) );
  HS65_LH_CBI4I6X2 U16108 ( .A(n14818), .B(n17607), .C(n14817), .D(n33880), 
        .Z(n14819) );
  HS65_LH_AOI31X2 U16109 ( .A(n14822), .B(n35562), .C(n14820), .D(n14819), .Z(
        n14823) );
  HS65_LH_OR2X4 U16110 ( .A(n14952), .B(n15120), .Z(n14968) );
  HS65_LH_OAI211X1 U16111 ( .A(n15327), .B(n14824), .C(n14823), .D(n14968), 
        .Z(n14825) );
  HS65_LH_AOI211X1 U16112 ( .A(n15499), .B(n14842), .C(n15030), .D(n14825), 
        .Z(n14826) );
  HS65_LH_AOI22X1 U16113 ( .A(n15331), .B(n14991), .C(n15075), .D(n14992), .Z(
        n14953) );
  HS65_LH_OAI22X1 U16114 ( .A(n14828), .B(n14827), .C(n14953), .D(n15344), .Z(
        n14836) );
  HS65_LH_AOI22X1 U16115 ( .A(n32629), .B(n14831), .C(n32748), .D(n14830), .Z(
        n14834) );
  HS65_LH_NAND2AX4 U16116 ( .A(n15234), .B(n14829), .Z(n15198) );
  HS65_LH_OAI22X1 U16117 ( .A(n33067), .B(n14831), .C(n17468), .D(n14830), .Z(
        n14832) );
  HS65_LH_OAI21X2 U16118 ( .A(n14832), .B(n33882), .C(n15198), .Z(n14833) );
  HS65_LH_OAI21X2 U16119 ( .A(n14834), .B(n15198), .C(n14833), .Z(n14835) );
  HS65_LH_NOR4ABX2 U16120 ( .A(n14837), .B(n14826), .C(n14836), .D(n14835), 
        .Z(n15566) );
  HS65_LH_AOI222X2 U16121 ( .A(n14995), .B(n15333), .C(n14842), .D(n15331), 
        .E(n14982), .F(n15329), .Z(n14873) );
  HS65_LH_NOR2X2 U16122 ( .A(n15328), .B(n14843), .Z(n14847) );
  HS65_LH_NOR2X2 U16123 ( .A(n14226), .B(n14852), .Z(n14846) );
  HS65_LH_NAND4ABX3 U16124 ( .A(n14847), .B(n14846), .C(n14845), .D(n14844), 
        .Z(n14858) );
  HS65_LH_OAI21X2 U16125 ( .A(n14852), .B(n33505), .C(n17523), .Z(n14848) );
  HS65_LH_CBI4I6X2 U16126 ( .A(n14850), .B(n14849), .C(n14848), .D(n15030), 
        .Z(n14851) );
  HS65_LH_OAI31X1 U16127 ( .A(n14853), .B(n14852), .C(n17471), .D(n14851), .Z(
        n14857) );
  HS65_LH_OAI22X1 U16128 ( .A(n14855), .B(n15399), .C(n14854), .D(n15120), .Z(
        n14856) );
  HS65_LH_AOI211X1 U16129 ( .A(n15499), .B(n14858), .C(n14857), .D(n14856), 
        .Z(n14871) );
  HS65_LH_IVX2 U16130 ( .A(n14862), .Z(n14860) );
  HS65_LH_OAI21X2 U16131 ( .A(n14861), .B(n32759), .C(n17638), .Z(n14859) );
  HS65_LH_AOI21X2 U16132 ( .A(n17591), .B(n14860), .C(n14859), .Z(n14867) );
  HS65_LH_AOI22X1 U16133 ( .A(n32629), .B(n14862), .C(n17590), .D(n14861), .Z(
        n14866) );
  HS65_LH_NOR2X2 U16134 ( .A(n14864), .B(n14863), .Z(n14865) );
  HS65_LH_MUXI21X2 U16135 ( .D0(n14867), .D1(n14866), .S0(n14865), .Z(n14868)
         );
  HS65_LH_AOI21X2 U16136 ( .A(n29624), .B(n14869), .C(n14868), .Z(n14870) );
  HS65_LH_IVX2 U16137 ( .A(n14878), .Z(n14886) );
  HS65_LH_AOI22X1 U16138 ( .A(n15102), .B(n15103), .C(n14879), .D(n15132), .Z(
        n14885) );
  HS65_LH_AOI222X2 U16139 ( .A(n14880), .B(n17523), .C(n14880), .D(n14881), 
        .E(n17523), .F(n33505), .Z(n14883) );
  HS65_LH_OAI31X1 U16140 ( .A(n14881), .B(n14880), .C(n17471), .D(n15098), .Z(
        n14882) );
  HS65_LH_AOI211X1 U16141 ( .A(n15100), .B(n15131), .C(n14883), .D(n14882), 
        .Z(n14884) );
  HS65_LH_OAI211X1 U16142 ( .A(n14886), .B(n15026), .C(n14885), .D(n14884), 
        .Z(n14904) );
  HS65_LH_AOI22X1 U16143 ( .A(n17590), .B(n14890), .C(n14887), .D(n15264), .Z(
        n14894) );
  HS65_LH_IVX2 U16144 ( .A(n14888), .Z(n15267) );
  HS65_LH_NAND2X2 U16145 ( .A(n15267), .B(n14889), .Z(n15218) );
  HS65_LH_OAI22X1 U16146 ( .A(n14891), .B(n17467), .C(n32759), .D(n14890), .Z(
        n14892) );
  HS65_LH_OAI21X2 U16147 ( .A(n14892), .B(n33882), .C(n15218), .Z(n14893) );
  HS65_LH_AOI22X1 U16149 ( .A(n15331), .B(n15074), .C(n15075), .D(n15073), .Z(
        n14896) );
  HS65_LH_OAI21X2 U16150 ( .A(n14895), .B(n14897), .C(n14896), .Z(n15125) );
  HS65_LH_OAI211X1 U16151 ( .A(n14898), .B(n14897), .C(n14896), .D(n14936), 
        .Z(n15127) );
  HS65_LH_AOI22X1 U16152 ( .A(n14900), .B(n15125), .C(n14899), .D(n15127), .Z(
        n14902) );
  HS65_LH_AOI22X1 U16153 ( .A(n15133), .B(n15110), .C(n15405), .D(n15101), .Z(
        n14901) );
  HS65_LH_NAND4ABX3 U16154 ( .A(n14904), .B(n14903), .C(n14902), .D(n14901), 
        .Z(n15563) );
  HS65_LH_FA1X4 U16155 ( .A0(\u_DataPath/pc_4_to_ex_i [4]), .B0(
        \u_DataPath/u_idexreg/N29 ), .CI(n14908), .CO(n14173), .S0(n14909) );
  HS65_LH_AOI22X1 U16156 ( .A(n17591), .B(n14913), .C(n17590), .D(n14912), .Z(
        n14940) );
  HS65_LH_NAND2AX4 U16157 ( .A(n14911), .B(n14910), .Z(n15214) );
  HS65_LH_OAI22X1 U16158 ( .A(n14913), .B(n17467), .C(n17468), .D(n14912), .Z(
        n14935) );
  HS65_LH_NAND4ABX3 U16159 ( .A(n14917), .B(n14916), .C(n14915), .D(n14914), 
        .Z(n15332) );
  HS65_LH_AOI22X1 U16160 ( .A(n15525), .B(n15332), .C(n15497), .D(n14993), .Z(
        n14933) );
  HS65_LH_CBI4I1X3 U16161 ( .A(n17587), .B(n14919), .C(n14918), .D(n17515), 
        .Z(n14920) );
  HS65_LH_OAI31X1 U16162 ( .A(n14922), .B(n14921), .C(n17471), .D(n14920), .Z(
        n14923) );
  HS65_LH_AOI21X2 U16163 ( .A(n15517), .B(n15334), .C(n14923), .Z(n14932) );
  HS65_LH_NOR2X2 U16164 ( .A(n14925), .B(n14924), .Z(n14980) );
  HS65_LH_NAND4ABX3 U16165 ( .A(n14929), .B(n14928), .C(n14927), .D(n14926), 
        .Z(n15330) );
  HS65_LH_AOI22X1 U16166 ( .A(n14930), .B(n14980), .C(n13892), .D(n15330), .Z(
        n14931) );
  HS65_LH_NAND3X2 U16167 ( .A(n14933), .B(n14932), .C(n14931), .Z(n14934) );
  HS65_LH_CBI4I6X2 U16168 ( .A(n33882), .B(n14935), .C(n15214), .D(n14934), 
        .Z(n14939) );
  HS65_LH_NOR2X2 U16169 ( .A(n17607), .B(n14936), .Z(n15043) );
  HS65_LH_IVX2 U16170 ( .A(n14937), .Z(n14994) );
  HS65_LH_AO222X4 U16171 ( .A(n15075), .B(n14994), .C(n15329), .D(n14991), .E(
        n15331), .F(n14992), .Z(n14979) );
  HS65_LH_OAI21X2 U16172 ( .A(n15043), .B(n14979), .C(n15529), .Z(n14938) );
  HS65_LH_NOR2X2 U16173 ( .A(n14943), .B(n17260), .Z(n14948) );
  HS65_LH_AOI21X2 U16174 ( .A(n14943), .B(n17260), .C(n14948), .Z(n15202) );
  HS65_LH_IVX2 U16175 ( .A(n14944), .Z(n15359) );
  HS65_LH_AOI22X1 U16176 ( .A(n17591), .B(n15359), .C(n17600), .D(n14946), .Z(
        n14961) );
  HS65_LH_AOI21X2 U16177 ( .A(n17591), .B(n14944), .C(n33882), .Z(n14945) );
  HS65_LH_OAI21X2 U16178 ( .A(n17468), .B(n14946), .C(n14945), .Z(n14959) );
  HS65_LH_AOI22X1 U16179 ( .A(n14948), .B(n17314), .C(n15102), .D(n14947), .Z(
        n14950) );
  HS65_LH_CBI4I1X3 U16180 ( .A(n17587), .B(n15239), .C(n14030), .D(n17515), 
        .Z(n14949) );
  HS65_LH_OAI211X1 U16181 ( .A(n14953), .B(n15079), .C(n14950), .D(n14949), 
        .Z(n14957) );
  HS65_LH_AOI22X1 U16182 ( .A(n13892), .B(n15334), .C(n15517), .D(n14993), .Z(
        n14951) );
  HS65_LH_CBI4I1X3 U16183 ( .A(n14953), .B(n14952), .C(n15080), .D(n14951), 
        .Z(n14956) );
  HS65_LH_IVX2 U16184 ( .A(n15006), .Z(n14981) );
  HS65_LH_AOI22X1 U16185 ( .A(n15499), .B(n14981), .C(n15497), .D(n14994), .Z(
        n14955) );
  HS65_LH_AOI22X1 U16186 ( .A(n15133), .B(n15003), .C(n15525), .D(n15330), .Z(
        n14954) );
  HS65_LH_NAND4ABX3 U16187 ( .A(n14957), .B(n14956), .C(n14955), .D(n14954), 
        .Z(n14958) );
  HS65_LH_AOI21X2 U16188 ( .A(n14959), .B(n33693), .C(n14958), .Z(n14960) );
  HS65_LH_NOR2X2 U16189 ( .A(\u_DataPath/u_execute/A_inALU_i [20]), .B(n15271), 
        .Z(n14965) );
  HS65_LH_CBI4I6X2 U16190 ( .A(n15272), .B(n33505), .C(n17523), .D(n14965), 
        .Z(n14971) );
  HS65_LH_NAND2X2 U16191 ( .A(\u_DataPath/u_execute/A_inALU_i [20]), .B(n15271), .Z(n14967) );
  HS65_LH_OAI22X1 U16192 ( .A(n15245), .B(n14968), .C(n17471), .D(n14967), .Z(
        n14970) );
  HS65_LH_AOI22X1 U16193 ( .A(n15133), .B(n14995), .C(n15102), .D(n14996), .Z(
        n14969) );
  HS65_LH_NAND4ABX3 U16194 ( .A(n14971), .B(n14970), .C(n14969), .D(n15098), 
        .Z(n14986) );
  HS65_LH_IVX2 U16195 ( .A(n14975), .Z(n14972) );
  HS65_LH_AOI22X1 U16196 ( .A(n32629), .B(n14972), .C(n17590), .D(n14973), .Z(
        n14978) );
  HS65_LH_OAI21X2 U16197 ( .A(n14973), .B(n17468), .C(n17638), .Z(n14974) );
  HS65_LH_AOI21X2 U16198 ( .A(n17591), .B(n14975), .C(n14974), .Z(n14977) );
  HS65_LH_MUXI21X2 U16199 ( .D0(n14976), .D1(n15271), .S0(
        \u_DataPath/u_execute/A_inALU_i [20]), .Z(n15188) );
  HS65_LH_MUXI21X2 U16200 ( .D0(n14978), .D1(n14977), .S0(n15188), .Z(n14985)
         );
  HS65_LH_AOI22X1 U16201 ( .A(n29624), .B(n14980), .C(n15042), .D(n14979), .Z(
        n14984) );
  HS65_LH_AOI22X1 U16202 ( .A(n15499), .B(n14982), .C(n15405), .D(n14981), .Z(
        n14983) );
  HS65_LH_NAND4ABX3 U16203 ( .A(n14986), .B(n14985), .C(n14984), .D(n14983), 
        .Z(n15564) );
  HS65_LH_MX41X4 U16204 ( .D0(n14994), .S0(n15331), .D1(n14993), .S1(n15039), 
        .D2(n14992), .S2(n15329), .D3(n14991), .S3(n15333), .Z(n15381) );
  HS65_LH_AOI22X1 U16205 ( .A(n15133), .B(n14996), .C(n15499), .D(n14995), .Z(
        n15005) );
  HS65_LH_AOI21X2 U16206 ( .A(n17314), .B(n14998), .C(n17515), .Z(n15001) );
  HS65_LH_AOI21X2 U16207 ( .A(n17587), .B(n14998), .C(n14997), .Z(n15000) );
  HS65_LH_OAI22X1 U16208 ( .A(n15001), .B(n15000), .C(n14999), .D(n15327), .Z(
        n15002) );
  HS65_LH_AOI211X1 U16209 ( .A(n15405), .B(n15003), .C(n15030), .D(n15002), 
        .Z(n15004) );
  HS65_LH_OAI211X1 U16210 ( .A(n15006), .B(n15409), .C(n15005), .D(n15004), 
        .Z(n15014) );
  HS65_LH_OAI21X2 U16211 ( .A(n15009), .B(n17468), .C(n17638), .Z(n15007) );
  HS65_LH_AOI21X2 U16212 ( .A(n17591), .B(n15008), .C(n15007), .Z(n15012) );
  HS65_LH_IVX2 U16213 ( .A(n15008), .Z(n15010) );
  HS65_LH_AOI22X1 U16214 ( .A(n32629), .B(n15010), .C(n32748), .D(n15009), .Z(
        n15011) );
  HS65_LH_NOR2AX3 U16215 ( .A(n15284), .B(n15019), .Z(n15190) );
  HS65_LH_MUXI21X2 U16216 ( .D0(n15012), .D1(n15011), .S0(n15190), .Z(n15013)
         );
  HS65_LH_AOI21X2 U16217 ( .A(n15033), .B(n15018), .C(n15265), .Z(n15217) );
  HS65_LH_NOR2AX3 U16218 ( .A(n15020), .B(n15019), .Z(n15022) );
  HS65_LH_OAI21X2 U16219 ( .A(n15022), .B(n17467), .C(n17638), .Z(n15021) );
  HS65_LH_AOI21X2 U16220 ( .A(n32748), .B(n15023), .C(n15021), .Z(n15051) );
  HS65_LH_IVX2 U16221 ( .A(n15022), .Z(n15024) );
  HS65_LH_OAI22X1 U16222 ( .A(n33067), .B(n15024), .C(n32759), .D(n15023), .Z(
        n15049) );
  HS65_LH_IVX2 U16223 ( .A(n15025), .Z(n15028) );
  HS65_LH_OAI22X1 U16224 ( .A(n15028), .B(n15417), .C(n15027), .D(n15026), .Z(
        n15035) );
  HS65_LH_CBI4I6X2 U16225 ( .A(n15033), .B(n17523), .C(n15032), .D(n33880), 
        .Z(n15029) );
  HS65_LH_AOI211X1 U16226 ( .A(n15100), .B(n15498), .C(n15030), .D(n15029), 
        .Z(n15031) );
  HS65_LH_OAI31X1 U16227 ( .A(n15033), .B(n15032), .C(n17471), .D(n15031), .Z(
        n15034) );
  HS65_LH_AOI211X1 U16228 ( .A(n15405), .B(n15036), .C(n15035), .D(n15034), 
        .Z(n15046) );
  HS65_LH_MX41X4 U16229 ( .D0(n15041), .S0(n15331), .D1(n15040), .S1(n15039), 
        .D2(n15038), .S2(n15329), .D3(n15037), .S3(n15333), .Z(n15530) );
  HS65_LH_CBI4I1X3 U16230 ( .A(n15044), .B(n15043), .C(n15530), .D(n15042), 
        .Z(n15045) );
  HS65_LH_OAI211X1 U16231 ( .A(n15047), .B(n15409), .C(n15046), .D(n15045), 
        .Z(n15048) );
  HS65_LH_FA1X4 U16232 ( .A0(n8860), .B0(\u_DataPath/u_idexreg/N27 ), .CI(
        n15055), .CO(n14403), .S0(n15056) );
  HS65_LH_IVX2 U16233 ( .A(n15057), .Z(n15059) );
  HS65_LH_NOR4ABX2 U16234 ( .A(n15061), .B(n15060), .C(n15059), .D(n15058), 
        .Z(n15142) );
  HS65_LH_CBI4I6X2 U16235 ( .A(n15245), .B(n17523), .C(n15062), .D(n33880), 
        .Z(n15066) );
  HS65_LH_IVX2 U16236 ( .A(n15130), .Z(n15064) );
  HS65_LH_NAND2X2 U16237 ( .A(n15324), .B(n15069), .Z(n15068) );
  HS65_LH_OAI22X1 U16238 ( .A(n15064), .B(n15063), .C(n15068), .D(n17471), .Z(
        n15065) );
  HS65_LH_AOI211X1 U16239 ( .A(n15499), .B(n15132), .C(n15066), .D(n15065), 
        .Z(n15067) );
  HS65_LH_OAI21X2 U16240 ( .A(n15324), .B(n15069), .C(n15068), .Z(n15197) );
  HS65_LH_CBI4I1X3 U16241 ( .A(n15087), .B(n17590), .C(n15070), .D(n15197), 
        .Z(n15071) );
  HS65_LH_OAI211X1 U16242 ( .A(n15142), .B(n29699), .C(n15067), .D(n15071), 
        .Z(n15093) );
  HS65_LH_AO222X4 U16243 ( .A(n15129), .B(n15075), .C(n15074), .D(n15329), .E(
        n15073), .F(n15331), .Z(n15077) );
  HS65_LH_AOI21X2 U16244 ( .A(n15333), .B(n15076), .C(n15077), .Z(n15121) );
  HS65_LH_AOI21X2 U16245 ( .A(n15333), .B(n15078), .C(n15077), .Z(n15107) );
  HS65_LH_OAI22X1 U16246 ( .A(n15121), .B(n15080), .C(n15107), .D(n15079), .Z(
        n15092) );
  HS65_LH_NAND2X2 U16247 ( .A(n15324), .B(n14218), .Z(n15081) );
  HS65_LH_NAND4ABX3 U16248 ( .A(n15084), .B(n15083), .C(n15082), .D(n15081), 
        .Z(n15085) );
  HS65_LH_AOI22X1 U16249 ( .A(n15497), .B(n15138), .C(n15525), .D(n15085), .Z(
        n15091) );
  HS65_LH_OAI22X1 U16250 ( .A(n15087), .B(n17468), .C(n17467), .D(n15086), .Z(
        n15089) );
  HS65_LH_IVX2 U16251 ( .A(n15197), .Z(n15088) );
  HS65_LH_OAI21X2 U16252 ( .A(n33882), .B(n15089), .C(n15088), .Z(n15090) );
  HS65_LH_NAND4ABX3 U16253 ( .A(n15093), .B(n15092), .C(n15091), .D(n15090), 
        .Z(n15538) );
  HS65_LH_OAI211X1 U16254 ( .A(n33045), .B(n15096), .C(n17314), .D(n15095), 
        .Z(n15097) );
  HS65_LH_OAI211X1 U16255 ( .A(n33880), .B(n15099), .C(n15098), .D(n15097), 
        .Z(n15109) );
  HS65_LH_AOI22X1 U16256 ( .A(n15405), .B(n15131), .C(n15100), .D(n15132), .Z(
        n15105) );
  HS65_LH_AOI22X1 U16257 ( .A(n15133), .B(n15103), .C(n15102), .D(n15101), .Z(
        n15104) );
  HS65_LH_OAI211X1 U16258 ( .A(n15107), .B(n15106), .C(n15105), .D(n15104), 
        .Z(n15108) );
  HS65_LH_AOI211X1 U16259 ( .A(n15499), .B(n15110), .C(n15109), .D(n15108), 
        .Z(n15111) );
  HS65_LH_AOI21X2 U16260 ( .A(n15115), .B(n17591), .C(n33882), .Z(n15112) );
  HS65_LH_OAI21X2 U16261 ( .A(n15113), .B(n17468), .C(n15112), .Z(n15118) );
  HS65_LH_IVX2 U16262 ( .A(n15113), .Z(n15114) );
  HS65_LH_OAI22X1 U16263 ( .A(n15115), .B(n17467), .C(n17468), .D(n15114), .Z(
        n15117) );
  HS65_LH_NOR2AX3 U16264 ( .A(n15266), .B(n15116), .Z(n15231) );
  HS65_LH_MUXI21X2 U16265 ( .D0(n15118), .D1(n15117), .S0(n15231), .Z(n15119)
         );
  HS65_LH_AOI22X1 U16266 ( .A(n15128), .B(n15127), .C(n15126), .D(n15125), .Z(
        n15158) );
  HS65_LH_AOI22X1 U16267 ( .A(n13892), .B(n15130), .C(n15497), .D(n15129), .Z(
        n15157) );
  HS65_LH_AOI22X1 U16268 ( .A(n15133), .B(n15132), .C(n15499), .D(n15131), .Z(
        n15140) );
  HS65_LH_CBI4I1X3 U16269 ( .A(n17587), .B(n15134), .C(n14029), .D(n17515), 
        .Z(n15135) );
  HS65_LH_OAI31X1 U16270 ( .A(n15147), .B(n33513), .C(n17471), .D(n15135), .Z(
        n15137) );
  HS65_LH_AOI21X2 U16271 ( .A(n15517), .B(n15138), .C(n15137), .Z(n15139) );
  HS65_LH_OAI211X1 U16272 ( .A(n15142), .B(n15141), .C(n15140), .D(n15139), 
        .Z(n15156) );
  HS65_LH_OAI21X2 U16273 ( .A(n15145), .B(n15144), .C(n15143), .Z(n15148) );
  HS65_LH_AOI22X1 U16274 ( .A(n17591), .B(n15148), .C(n17600), .D(n15150), .Z(
        n15154) );
  HS65_LH_OAI21X2 U16275 ( .A(n14029), .B(n15147), .C(n15146), .Z(n15201) );
  HS65_LH_OAI22X1 U16276 ( .A(n15150), .B(n17468), .C(n17467), .D(n15148), .Z(
        n15152) );
  HS65_LH_OAI21X2 U16277 ( .A(n15152), .B(n33882), .C(n15201), .Z(n15153) );
  HS65_LH_OAI21X2 U16278 ( .A(n15154), .B(n15201), .C(n15153), .Z(n15155) );
  HS65_LH_NOR4ABX2 U16279 ( .A(n15158), .B(n15157), .C(n15156), .D(n15155), 
        .Z(n15545) );
  HS65_LH_FA1X4 U16280 ( .A0(n10766), .B0(\u_DataPath/u_idexreg/N26 ), .CI(
        n15164), .CO(n15055), .S0(n15162) );
  HS65_LH_CNIVX3 U16281 ( .A(n12416), .Z(n15167) );
  HS65_LH_CNIVX3 U16282 ( .A(n12395), .Z(n15168) );
  HS65_LH_CNIVX3 U16283 ( .A(n12438), .Z(n15169) );
  HS65_LH_OAI212X3 U16284 ( .A(n17518), .B(n17696), .C(n17619), .D(n17584), 
        .E(n17844), .Z(n15174) );
  HS65_LH_CNIVX3 U16285 ( .A(n12471), .Z(n15170) );
  HS65_LH_OAI22X1 U16286 ( .A(n17506), .B(n17701), .C(n17628), .D(n17694), .Z(
        n15171) );
  HS65_LH_AOI212X2 U16287 ( .A(n17506), .B(n17701), .C(n17694), .D(n17628), 
        .E(n15171), .Z(n15172) );
  HS65_LH_OAI21X2 U16288 ( .A(n17648), .B(n17508), .C(n15172), .Z(n15173) );
  HS65_LH_CNIVX3 U16289 ( .A(n12327), .Z(n1928) );
  HS65_LH_OAI22X1 U16290 ( .A(n17506), .B(n17728), .C(n17508), .D(n17709), .Z(
        n15178) );
  HS65_LH_CNIVX3 U16291 ( .A(n12370), .Z(n15179) );
  HS65_LH_OAI22X1 U16292 ( .A(n17480), .B(n17707), .C(n17702), .D(n17628), .Z(
        n15180) );
  HS65_LH_NAND4ABX3 U16293 ( .A(n9508), .B(n15177), .C(n15182), .D(n15181), 
        .Z(n15183) );
  HS65_LH_CNIVX3 U16294 ( .A(n15702), .Z(n15186) );
  HS65_LH_NAND2X2 U16295 ( .A(n14070), .B(n10729), .Z(n15703) );
  HS65_LH_NOR4ABX2 U16296 ( .A(n15190), .B(n15189), .C(n15188), .D(n15187), 
        .Z(n15191) );
  HS65_LH_NAND3X2 U16297 ( .A(n15193), .B(n15192), .C(n15191), .Z(n15229) );
  HS65_LH_NAND2X2 U16298 ( .A(n15195), .B(n15502), .Z(n15194) );
  HS65_LH_OAI21X2 U16299 ( .A(n15195), .B(n15502), .C(n15194), .Z(n15515) );
  HS65_LH_NAND4ABX3 U16300 ( .A(n15198), .B(n15515), .C(n15197), .D(n15196), 
        .Z(n15199) );
  HS65_LH_NOR4ABX2 U16301 ( .A(n15200), .B(n15513), .C(n15335), .D(n15199), 
        .Z(n15225) );
  HS65_LH_NOR4ABX2 U16302 ( .A(n15351), .B(n15203), .C(n33693), .D(n15201), 
        .Z(n15223) );
  HS65_LH_NOR4ABX2 U16303 ( .A(n15370), .B(n15206), .C(n15205), .D(n15204), 
        .Z(n15222) );
  HS65_LH_MUX21I1X3 U16304 ( .D0(n29693), .D1(n38578), .S0(n17608), .Z(n15717)
         );
  HS65_LH_NAND2X2 U16305 ( .A(n15717), .B(n38579), .Z(n15352) );
  HS65_LH_IVX2 U16306 ( .A(n15352), .Z(n15728) );
  HS65_LH_NOR2X2 U16307 ( .A(n15717), .B(n38579), .Z(n15724) );
  HS65_LH_NOR2X2 U16308 ( .A(n15728), .B(n38565), .Z(n15427) );
  HS65_LH_NAND4ABX3 U16309 ( .A(n15215), .B(n15214), .C(n15427), .D(n15213), 
        .Z(n15221) );
  HS65_LH_NAND4ABX3 U16310 ( .A(n15219), .B(n15218), .C(n15217), .D(n15216), 
        .Z(n15220) );
  HS65_LH_NOR4ABX2 U16311 ( .A(n15223), .B(n15222), .C(n15221), .D(n15220), 
        .Z(n15224) );
  HS65_LH_NAND4ABX3 U16312 ( .A(n15227), .B(n15226), .C(n15225), .D(n15224), 
        .Z(n15228) );
  HS65_LH_NOR4ABX2 U16313 ( .A(n15231), .B(n15230), .C(n15229), .D(n15228), 
        .Z(n15323) );
  HS65_LH_IVX2 U16314 ( .A(n15233), .Z(n15232) );
  HS65_LH_CBI4I1X3 U16315 ( .A(n15232), .B(n15291), .C(n15290), .D(n15235), 
        .Z(n15367) );
  HS65_LH_NOR3AX2 U16316 ( .A(n15235), .B(n15234), .C(n15233), .Z(n15312) );
  HS65_LH_NOR2AX3 U16317 ( .A(n15367), .B(n15312), .Z(n15364) );
  HS65_LH_OAI211X1 U16318 ( .A(n17250), .B(n15237), .C(n15255), .D(n15236), 
        .Z(n15256) );
  HS65_LH_OAI211X1 U16319 ( .A(n17260), .B(n15239), .C(n15300), .D(n15254), 
        .Z(n15304) );
  HS65_LH_NOR2X2 U16320 ( .A(n15256), .B(n15304), .Z(n15288) );
  HS65_LH_AOI21X2 U16321 ( .A(n15500), .B(n15505), .C(n15241), .Z(n15243) );
  HS65_LH_AOI21X2 U16322 ( .A(n15244), .B(n15243), .C(n15242), .Z(n15250) );
  HS65_LH_OAI211X1 U16323 ( .A(n14037), .B(n15246), .C(n15245), .D(n15324), 
        .Z(n15249) );
  HS65_LH_CB4I1X4 U16324 ( .A(n15250), .B(n15249), .C(n15248), .D(n15247), .Z(
        n15310) );
  HS65_LH_NOR2X2 U16325 ( .A(n15306), .B(n15302), .Z(n15261) );
  HS65_LH_IVX2 U16326 ( .A(n15251), .Z(n15257) );
  HS65_LH_OAI211X1 U16327 ( .A(\u_DataPath/u_execute/A_inALU_i [12]), .B(
        n15252), .C(n15258), .D(n15257), .Z(n15305) );
  HS65_LH_AOI31X2 U16328 ( .A(n15300), .B(n15254), .C(n15253), .D(n15305), .Z(
        n15260) );
  HS65_LH_IVX2 U16329 ( .A(n15255), .Z(n15259) );
  HS65_LH_OA112X4 U16330 ( .A(n15259), .B(n15258), .C(n15257), .D(n15256), .Z(
        n15307) );
  HS65_LH_CBI4I6X2 U16331 ( .A(n15262), .B(n15261), .C(n15260), .D(n15307), 
        .Z(n15287) );
  HS65_LH_AOI21X2 U16332 ( .A(n15288), .B(n15310), .C(n15287), .Z(n15295) );
  HS65_LH_IVX2 U16333 ( .A(n15263), .Z(n15283) );
  HS65_LH_OAI211X1 U16334 ( .A(n15271), .B(n15272), .C(n15264), .D(n15283), 
        .Z(n15278) );
  HS65_LH_NAND3AX3 U16335 ( .A(n15278), .B(n15276), .C(n15273), .Z(n15294) );
  HS65_LH_NOR3AX2 U16336 ( .A(n15266), .B(n15274), .C(n15265), .Z(n15286) );
  HS65_LH_IVX2 U16337 ( .A(n15277), .Z(n15270) );
  HS65_LH_OAI21X2 U16338 ( .A(n15269), .B(n15268), .C(n15267), .Z(n15282) );
  HS65_LH_AOI211X1 U16339 ( .A(n15271), .B(n15272), .C(n15270), .D(n15282), 
        .Z(n15285) );
  HS65_LH_NAND2X2 U16340 ( .A(n15272), .B(n15271), .Z(n15280) );
  HS65_LH_IVX2 U16341 ( .A(n15286), .Z(n15275) );
  HS65_LH_OAI22X1 U16342 ( .A(n15276), .B(n15275), .C(n15274), .D(n15273), .Z(
        n15279) );
  HS65_LH_CBI4I1X3 U16343 ( .A(n15280), .B(n15279), .C(n15278), .D(n15277), 
        .Z(n15281) );
  HS65_LH_AOI21X2 U16344 ( .A(n15283), .B(n15282), .C(n15281), .Z(n15308) );
  HS65_LH_AOI31X2 U16345 ( .A(n15286), .B(n15285), .C(n15284), .D(n15308), .Z(
        n15356) );
  HS65_LH_IVX2 U16346 ( .A(n15356), .Z(n15293) );
  HS65_LH_AOI21X2 U16347 ( .A(n15288), .B(n15359), .C(n15287), .Z(n15289) );
  HS65_LH_OAI21X2 U16348 ( .A(n15289), .B(n15294), .C(n15293), .Z(n15354) );
  HS65_LH_NOR2X2 U16349 ( .A(n15291), .B(n15290), .Z(n15355) );
  HS65_LH_OAI21X2 U16350 ( .A(n17283), .B(n15354), .C(n15355), .Z(n15292) );
  HS65_LH_CBI4I6X2 U16351 ( .A(n15295), .B(n15294), .C(n15293), .D(n15292), 
        .Z(n15297) );
  HS65_LH_NOR3AX2 U16352 ( .A(n15351), .B(n15349), .C(n38565), .Z(n15316) );
  HS65_LH_NOR2X2 U16353 ( .A(n15311), .B(n15296), .Z(n15391) );
  HS65_LH_OAI31X1 U16354 ( .A(n15349), .B(n15391), .C(n38565), .D(n15352), .Z(
        n15315) );
  HS65_LH_CBI4I6X2 U16355 ( .A(n15364), .B(n15297), .C(n15316), .D(n15315), 
        .Z(n15321) );
  HS65_LH_NAND4ABX3 U16356 ( .A(n15306), .B(n15305), .C(n15299), .D(n15298), 
        .Z(n15358) );
  HS65_LH_OAI21X2 U16357 ( .A(n15302), .B(n15301), .C(n15300), .Z(n15303) );
  HS65_LH_NAND4ABX3 U16358 ( .A(n15306), .B(n15305), .C(n15304), .D(n15303), 
        .Z(n15309) );
  HS65_LH_NOR3AX2 U16359 ( .A(n15309), .B(n15308), .C(n15307), .Z(n15357) );
  HS65_LH_CB4I6X4 U16360 ( .A(n15358), .B(n15310), .C(n15357), .D(n15356), .Z(
        n15366) );
  HS65_LH_IVX2 U16361 ( .A(n15311), .Z(n15369) );
  HS65_LH_NAND3X2 U16362 ( .A(n15370), .B(n15369), .C(n15352), .Z(n15314) );
  HS65_LH_NOR2AX3 U16363 ( .A(n15312), .B(n15314), .Z(n15361) );
  HS65_LH_IVX2 U16364 ( .A(n15361), .Z(n15313) );
  HS65_LH_OAI21X2 U16365 ( .A(n15366), .B(n15313), .C(n17283), .Z(n15318) );
  HS65_LH_OAI22X1 U16366 ( .A(n15316), .B(n15315), .C(n15367), .D(n15314), .Z(
        n15360) );
  HS65_LH_IVX2 U16367 ( .A(n15323), .Z(n15317) );
  HS65_LH_OAI21X2 U16368 ( .A(n15318), .B(n15360), .C(n15317), .Z(n15320) );
  HS65_LH_AOI212X2 U16369 ( .A(n15321), .B(n17606), .C(n15320), .D(n17607), 
        .E(n17605), .Z(n15322) );
  HS65_LH_AOI31X2 U16370 ( .A(n17473), .B(n33045), .C(n15323), .D(n15322), .Z(
        n15386) );
  HS65_LH_NAND2X2 U16371 ( .A(n15325), .B(n15324), .Z(n15326) );
  HS65_LH_OAI211X1 U16372 ( .A(n15328), .B(n15505), .C(n15327), .D(n15326), 
        .Z(n15347) );
  HS65_LH_AOI222X2 U16373 ( .A(n15334), .B(n15333), .C(n15332), .D(n15331), 
        .E(n15330), .F(n15329), .Z(n15345) );
  HS65_LH_IVX2 U16374 ( .A(n15513), .Z(n15492) );
  HS65_LH_NOR2X2 U16375 ( .A(n15492), .B(n15335), .Z(n15336) );
  HS65_LH_AOI21X2 U16376 ( .A(n17469), .B(n17638), .C(n15336), .Z(n15340) );
  HS65_LH_AOI22X1 U16377 ( .A(n15499), .B(n14218), .C(n17314), .D(n15341), .Z(
        n15338) );
  HS65_LH_AOI21X2 U16378 ( .A(n33880), .B(n15338), .C(n15337), .Z(n15339) );
  HS65_LH_AOI211X1 U16379 ( .A(n17587), .B(n15341), .C(n15340), .D(n15339), 
        .Z(n15343) );
  HS65_LH_OAI21X2 U16380 ( .A(n15345), .B(n15344), .C(n15343), .Z(n15346) );
  HS65_LH_CBI4I6X2 U16381 ( .A(n15348), .B(n15347), .C(n15525), .D(n15346), 
        .Z(n15384) );
  HS65_LH_NOR2X2 U16382 ( .A(n15349), .B(n15728), .Z(n15722) );
  HS65_LH_IVX2 U16383 ( .A(n15391), .Z(n15350) );
  HS65_LH_AOI21X2 U16384 ( .A(n15722), .B(n15350), .C(n38565), .Z(n15377) );
  HS65_LH_NAND3X2 U16385 ( .A(n33227), .B(n15352), .C(n15351), .Z(n15376) );
  HS65_LH_IVX2 U16386 ( .A(n15376), .Z(n15353) );
  HS65_LH_CBI4I1X3 U16387 ( .A(n15355), .B(n15354), .C(n15364), .D(n15353), 
        .Z(n15363) );
  HS65_LH_CBI4I6X2 U16388 ( .A(n15359), .B(n15358), .C(n15357), .D(n15356), 
        .Z(n15365) );
  HS65_LH_AOI21X2 U16389 ( .A(n15365), .B(n15361), .C(n15360), .Z(n15362) );
  HS65_LH_AO32X4 U16390 ( .A(n15377), .B(n17606), .C(n15363), .D(n17607), .E(
        n15362), .Z(n15379) );
  HS65_LH_IVX2 U16391 ( .A(n15364), .Z(n15373) );
  HS65_LH_IVX2 U16392 ( .A(n15365), .Z(n15368) );
  HS65_LH_OAI211X1 U16393 ( .A(n17607), .B(n15368), .C(n15367), .D(n15366), 
        .Z(n15372) );
  HS65_LH_NAND2X2 U16394 ( .A(n15370), .B(n15369), .Z(n15371) );
  HS65_LH_NOR4ABX2 U16395 ( .A(n15373), .B(n15372), .C(n38565), .D(n15371), 
        .Z(n15375) );
  HS65_LH_CBI4I1X3 U16396 ( .A(n15377), .B(n15376), .C(n15375), .D(n17473), 
        .Z(n15378) );
  HS65_LH_CBI4I6X2 U16397 ( .A(n17475), .B(n15379), .C(n15378), .D(n17328), 
        .Z(n15382) );
  HS65_LH_AOI22X1 U16398 ( .A(n17266), .B(n15382), .C(n15529), .D(n15381), .Z(
        n15383) );
  HS65_LH_NAND2X2 U16399 ( .A(n15391), .B(n15390), .Z(n15721) );
  HS65_LH_NAND2X2 U16400 ( .A(n33227), .B(n15721), .Z(n15719) );
  HS65_LH_PAOI2X1 U16402 ( .A(n40560), .B(n15395), .P(n15394), .Z(n15718) );
  HS65_LH_OAI21X2 U16403 ( .A(n17463), .B(n17307), .C(n17599), .Z(n15424) );
  HS65_LH_OAI22X1 U16404 ( .A(n38568), .B(n17638), .C(n15399), .D(n15398), .Z(
        n15420) );
  HS65_LH_NAND4ABX3 U16405 ( .A(n15403), .B(n15402), .C(n15401), .D(n15400), 
        .Z(n15406) );
  HS65_LH_AOI22X1 U16406 ( .A(n15499), .B(n15406), .C(n15405), .D(n15404), .Z(
        n15416) );
  HS65_LH_OAI22X1 U16407 ( .A(n15717), .B(n17471), .C(n17607), .D(n35213), .Z(
        n15413) );
  HS65_LH_OAI22X1 U16408 ( .A(n15717), .B(n17523), .C(n15410), .D(n15409), .Z(
        n15412) );
  HS65_LH_CBI4I6X2 U16409 ( .A(n17515), .B(n15413), .C(n38579), .D(n15412), 
        .Z(n15415) );
  HS65_LH_OAI211X1 U16410 ( .A(n15418), .B(n15417), .C(n15416), .D(n15415), 
        .Z(n15419) );
  HS65_LH_AOI211X1 U16411 ( .A(n29624), .B(n15421), .C(n15420), .D(n15419), 
        .Z(n15423) );
  HS65_LH_CBI4I1X3 U16412 ( .A(n17307), .B(n17463), .C(n15424), .D(n17272), 
        .Z(n15425) );
  HS65_LH_CNIVX3 U16413 ( .A(n13887), .Z(n15428) );
  HS65_LH_CNIVX3 U16414 ( .A(n13885), .Z(n15429) );
  HS65_LH_CNIVX3 U16415 ( .A(n13890), .Z(n15430) );
  HS65_LH_CNIVX3 U16416 ( .A(n13646), .Z(n15470) );
  HS65_LH_FA1X4 U16417 ( .A0(n17549), .B0(n18000), .CI(n15471), .CO(n15472), 
        .S0(n14192) );
  HS65_LHS_XOR3X2 U16418 ( .A(n17550), .B(n15472), .C(n17526), .Z(n15473) );
  HS65_LH_CNIVX3 U16419 ( .A(n13650), .Z(n15474) );
  HS65_LH_OAI22X1 U16420 ( .A(n17623), .B(n17707), .C(n17620), .D(n17705), .Z(
        n15479) );
  HS65_LH_AOI212X2 U16421 ( .A(n17623), .B(n17707), .C(n17704), .D(n17620), 
        .E(n15479), .Z(n15480) );
  HS65_LH_OAI212X3 U16422 ( .A(n17497), .B(n40191), .C(n17621), .D(n17702), 
        .E(n15480), .Z(n15481) );
  HS65_LH_AOI212X2 U16423 ( .A(n17650), .B(n40615), .C(n17622), .D(n17709), 
        .E(n15481), .Z(n15482) );
  HS65_LH_CNIVX3 U16424 ( .A(n12382), .Z(n1113) );
  HS65_LH_MUXI21X2 U16425 ( .D0(n40440), .D1(n17694), .S0(n17497), .Z(n15484)
         );
  HS65_LH_AOI212X2 U16426 ( .A(n17698), .B(n17623), .C(n40236), .D(n17499), 
        .E(n15484), .Z(n15486) );
  HS65_LH_OAI212X3 U16427 ( .A(n17492), .B(n40170), .C(n17624), .D(n17701), 
        .E(n15486), .Z(n15487) );
  HS65_LH_AOI212X2 U16428 ( .A(n17651), .B(n27626), .C(n17620), .D(n17696), 
        .E(n15487), .Z(n15489) );
  HS65_LH_AOI22X1 U16429 ( .A(n39479), .B(n39477), .C(n15483), .D(n39476), .Z(
        n137) );
  HS65_LH_NAND2X2 U16430 ( .A(n17591), .B(n15492), .Z(n15494) );
  HS65_LH_CBI4I6X2 U16431 ( .A(n32759), .B(n15512), .C(n15494), .D(n15515), 
        .Z(n15535) );
  HS65_LH_AOI22X1 U16432 ( .A(n15499), .B(n15498), .C(n15497), .D(n15496), .Z(
        n15504) );
  HS65_LH_OAI211X1 U16433 ( .A(n17606), .B(n15502), .C(n17314), .D(n15500), 
        .Z(n15503) );
  HS65_LH_NOR2X2 U16434 ( .A(n15508), .B(n15507), .Z(n15527) );
  HS65_LH_NAND3X2 U16435 ( .A(n15511), .B(n15510), .C(n15509), .Z(n15526) );
  HS65_LH_AOI22X1 U16436 ( .A(n32629), .B(n15513), .C(n17590), .D(n15512), .Z(
        n15523) );
  HS65_LH_IVX2 U16437 ( .A(n15515), .Z(n15521) );
  HS65_LH_AOI22X1 U16438 ( .A(n13892), .B(n15518), .C(n15517), .D(n15516), .Z(
        n15520) );
  HS65_LH_CBI4I1X3 U16439 ( .A(n15523), .B(n17638), .C(n15521), .D(n15520), 
        .Z(n15524) );
  HS65_LH_CBI4I6X2 U16440 ( .A(n15527), .B(n15526), .C(n15525), .D(n15524), 
        .Z(n15533) );
  HS65_LH_NOR2X2 U16441 ( .A(n14037), .B(n15528), .Z(n15531) );
  HS65_LH_CBI4I1X3 U16442 ( .A(n32353), .B(n15531), .C(n15530), .D(n15529), 
        .Z(n15532) );
  HS65_LH_NAND4ABX3 U16443 ( .A(n15535), .B(n15534), .C(n15533), .D(n15532), 
        .Z(n15536) );
  HS65_LH_NOR3X1 U16444 ( .A(n33858), .B(n33796), .C(n32999), .Z(n15539) );
  HS65_LH_NAND4ABX3 U16445 ( .A(n32506), .B(n33732), .C(n33562), .D(n15539), 
        .Z(n15543) );
  HS65_LH_NOR4ABX2 U16446 ( .A(n33616), .B(n33520), .C(n33259), .D(n15543), 
        .Z(n15547) );
  HS65_LH_NAND4ABX3 U16447 ( .A(n33477), .B(n33689), .C(n32930), .D(n15547), 
        .Z(n15553) );
  HS65_LH_NAND4ABX3 U16448 ( .A(n33020), .B(n15553), .C(n32774), .D(n32880), 
        .Z(n15555) );
  HS65_LH_NOR4ABX2 U16449 ( .A(n15558), .B(n32637), .C(n15556), .D(n15555), 
        .Z(n15561) );
  HS65_LH_NOR4ABX2 U16450 ( .A(n15562), .B(n15561), .C(n32517), .D(n32710), 
        .Z(n15565) );
  HS65_LH_NOR4ABX2 U16451 ( .A(n15566), .B(n15565), .C(n15564), .D(n15563), 
        .Z(n15569) );
  HS65_LH_NOR4ABX2 U16452 ( .A(n17273), .B(n17271), .C(n17282), .D(n17318), 
        .Z(n15571) );
  HS65_LH_NAND4ABX3 U16453 ( .A(n17276), .B(n17275), .C(n15572), .D(n15571), 
        .Z(n15575) );
  HS65_LH_NOR2X2 U16454 ( .A(n15641), .B(n14111), .Z(n15640) );
  HS65_LHS_XOR3X2 U16455 ( .A(n29692), .B(n17550), .C(n15579), .Z(n15580) );
  HS65_LH_FA1X4 U16456 ( .A0(n29693), .B0(n17549), .CI(n15581), .CO(n15579), 
        .S0(n15582) );
  HS65_LH_FA1X4 U16457 ( .A0(n29692), .B0(n17548), .CI(n15583), .CO(n15581), 
        .S0(n15584) );
  HS65_LH_FA1X4 U16458 ( .A0(n29693), .B0(n17547), .CI(n15585), .CO(n15583), 
        .S0(n15586) );
  HS65_LH_FA1X4 U16459 ( .A0(n29692), .B0(n17546), .CI(n15587), .CO(n15585), 
        .S0(n15588) );
  HS65_LH_FA1X4 U16460 ( .A0(n29693), .B0(n17545), .CI(n15589), .CO(n15587), 
        .S0(n15590) );
  HS65_LH_FA1X4 U16461 ( .A0(n29692), .B0(n17544), .CI(n15591), .CO(n15589), 
        .S0(n15592) );
  HS65_LH_FA1X4 U16462 ( .A0(n29693), .B0(n17543), .CI(n15593), .CO(n15591), 
        .S0(n15594) );
  HS65_LH_FA1X4 U16463 ( .A0(n29692), .B0(n17542), .CI(n15595), .CO(n15593), 
        .S0(n15596) );
  HS65_LH_FA1X4 U16464 ( .A0(n29693), .B0(n17541), .CI(n15597), .CO(n15595), 
        .S0(n15598) );
  HS65_LH_FA1X4 U16465 ( .A0(n29692), .B0(n17540), .CI(n15599), .CO(n15597), 
        .S0(n15600) );
  HS65_LH_FA1X4 U16466 ( .A0(n29693), .B0(n17539), .CI(n15601), .CO(n15599), 
        .S0(n15602) );
  HS65_LH_FA1X4 U16467 ( .A0(n29692), .B0(n17538), .CI(n15603), .CO(n15601), 
        .S0(n15604) );
  HS65_LH_FA1X4 U16468 ( .A0(n17527), .B0(n17537), .CI(n15605), .CO(n15603), 
        .S0(n15606) );
  HS65_LH_FA1X4 U16469 ( .A0(n17527), .B0(n17536), .CI(n15607), .CO(n15605), 
        .S0(n15608) );
  HS65_LH_FA1X4 U16470 ( .A0(n17527), .B0(n17535), .CI(n15609), .CO(n15607), 
        .S0(n15610) );
  HS65_LH_FA1X4 U16471 ( .A0(n18158), .B0(n17534), .CI(n15611), .CO(n15609), 
        .S0(n15612) );
  HS65_LH_FA1X4 U16472 ( .A0(n17560), .B0(n17533), .CI(n15613), .CO(n15611), 
        .S0(n15614) );
  HS65_LH_FA1X4 U16473 ( .A0(n17559), .B0(n17532), .CI(n15615), .CO(n15613), 
        .S0(n15616) );
  HS65_LH_FA1X4 U16474 ( .A0(n17558), .B0(n17531), .CI(n15617), .CO(n15615), 
        .S0(n15618) );
  HS65_LH_FA1X4 U16475 ( .A0(n17557), .B0(n17530), .CI(n15619), .CO(n15617), 
        .S0(n15620) );
  HS65_LH_FA1X4 U16476 ( .A0(n17556), .B0(n17529), .CI(n17270), .CO(n15619), 
        .S0(n15622) );
  HS65_LH_FA1X4 U16477 ( .A0(\u_DataPath/u_idexreg/N34 ), .B0(
        \u_DataPath/pc_4_to_ex_i [9]), .CI(n15623), .CO(n15621), .S0(n15624)
         );
  HS65_LH_FA1X4 U16478 ( .A0(\u_DataPath/u_idexreg/N33 ), .B0(
        \u_DataPath/pc_4_to_ex_i [8]), .CI(n15625), .CO(n15623), .S0(n15626)
         );
  HS65_LH_FA1X4 U16479 ( .A0(\u_DataPath/u_idexreg/N32 ), .B0(
        \u_DataPath/pc_4_to_ex_i [7]), .CI(n15627), .CO(n15625), .S0(n15628)
         );
  HS65_LH_FA1X4 U16480 ( .A0(\u_DataPath/u_idexreg/N31 ), .B0(
        \u_DataPath/pc_4_to_ex_i [6]), .CI(n15629), .CO(n15627), .S0(n15630)
         );
  HS65_LH_FA1X4 U16481 ( .A0(\u_DataPath/u_idexreg/N30 ), .B0(
        \u_DataPath/pc_4_to_ex_i [5]), .CI(n15631), .CO(n15629), .S0(n15632)
         );
  HS65_LH_FA1X4 U16482 ( .A0(\u_DataPath/u_idexreg/N29 ), .B0(
        \u_DataPath/pc_4_to_ex_i [4]), .CI(n15633), .CO(n15631), .S0(n15634)
         );
  HS65_LH_FA1X4 U16483 ( .A0(\u_DataPath/u_idexreg/N28 ), .B0(
        \u_DataPath/pc_4_to_ex_i [3]), .CI(n15635), .CO(n15633), .S0(n15636)
         );
  HS65_LH_FA1X4 U16484 ( .A0(\u_DataPath/u_idexreg/N27 ), .B0(
        \u_DataPath/pc_4_to_ex_i [2]), .CI(n15637), .CO(n15635), .S0(n15638)
         );
  HS65_LH_FA1X4 U16485 ( .A0(\u_DataPath/u_idexreg/N26 ), .B0(
        \u_DataPath/u_execute/link_value_i [1]), .CI(n15640), .CO(n15637), 
        .S0(n15639) );
  HS65_LH_CNIVX3 U16486 ( .A(n13879), .Z(n15643) );
  HS65_LH_CNIVX3 U16487 ( .A(n15711), .Z(n15712) );
  HS65_LH_CNIVX3 U16488 ( .A(n15714), .Z(n15710) );
  HS65_LH_NAND3X5 U16489 ( .A(n15670), .B(n15712), .C(n15710), .Z(n111) );
  HS65_LH_NOR2AX3 U16490 ( .A(\u_DataPath/mem_writedata_out_i [11]), .B(n15694), .Z(n15672) );
  HS65_LH_NOR2AX3 U16491 ( .A(\u_DataPath/mem_writedata_out_i [15]), .B(n15694), .Z(n15675) );
  HS65_LH_NOR2AX3 U16492 ( .A(\u_DataPath/mem_writedata_out_i [9]), .B(n15694), 
        .Z(n15677) );
  HS65_LH_NOR2AX3 U16493 ( .A(\u_DataPath/mem_writedata_out_i [12]), .B(n15694), .Z(n15679) );
  HS65_LH_NOR2AX3 U16494 ( .A(\u_DataPath/mem_writedata_out_i [13]), .B(n15694), .Z(n15681) );
  HS65_LH_NOR2AX3 U16495 ( .A(\u_DataPath/mem_writedata_out_i [14]), .B(n15694), .Z(n15683) );
  HS65_LH_NOR2AX3 U16496 ( .A(\u_DataPath/mem_writedata_out_i [8]), .B(n15694), 
        .Z(n15685) );
  HS65_LH_NOR2AX3 U16497 ( .A(\u_DataPath/mem_writedata_out_i [10]), .B(n15694), .Z(n15688) );
  HS65_LL_AND2ABX18 U16498 ( .A(n14078), .B(n15697), .Z(Address_toRAM_18) );
  HS65_LL_AND2ABX18 U16499 ( .A(n14078), .B(n15698), .Z(Address_toRAM_12) );
  HS65_LL_AND2ABX18 U16500 ( .A(n15700), .B(n15699), .Z(Address_toRAM_0) );
  HS65_LL_NOR2AX25 U16501 ( .A(\u_DataPath/mem_writedata_out_i [26]), .B(
        n14072), .Z(Data_in_26) );
  HS65_LL_NOR2AX25 U16502 ( .A(\u_DataPath/mem_writedata_out_i [25]), .B(
        n14072), .Z(Data_in_25) );
  HS65_LL_NOR2AX25 U16503 ( .A(\u_DataPath/mem_writedata_out_i [24]), .B(
        n14072), .Z(Data_in_24) );
  HS65_LL_NOR2AX25 U16504 ( .A(\u_DataPath/mem_writedata_out_i [23]), .B(
        n14072), .Z(Data_in_23) );
  HS65_LH_NOR2X3 U16505 ( .A(n10732), .B(n14026), .Z(n17198) );
  HS65_LL_OR2X18 U16506 ( .A(n17198), .B(n15750), .Z(\nibble[1]_snps_wire ) );
  HS65_LL_AND2X18 U16507 ( .A(\u_DataPath/mem_writedata_out_i [3]), .B(
        write_op_snps_wire), .Z(Data_in_3) );
  HS65_LL_AND2X18 U16508 ( .A(\u_DataPath/mem_writedata_out_i [4]), .B(
        write_op_snps_wire), .Z(Data_in_4) );
  HS65_LL_AND2X18 U16509 ( .A(\u_DataPath/mem_writedata_out_i [1]), .B(
        write_op_snps_wire), .Z(Data_in_1) );
  HS65_LL_AND2X18 U16510 ( .A(\u_DataPath/mem_writedata_out_i [2]), .B(
        write_op_snps_wire), .Z(Data_in_2) );
  HS65_LL_AND2X18 U16511 ( .A(\u_DataPath/mem_writedata_out_i [5]), .B(
        write_op_snps_wire), .Z(Data_in_5) );
  HS65_LL_AND2X18 U16512 ( .A(\u_DataPath/mem_writedata_out_i [6]), .B(
        write_op_snps_wire), .Z(Data_in_6) );
  HS65_LH_NAND2X2 U16514 ( .A(n13646), .B(n13879), .Z(n278) );
  HS65_LH_NAND2X2 U16515 ( .A(n13639), .B(n258), .Z(n282) );
  HS65_LH_CNIVX3 U16516 ( .A(n12482), .Z(n191) );
  HS65_LH_NOR3X1 U16517 ( .A(n15475), .B(n282), .C(n191), .Z(n17205) );
  HS65_LH_NOR2X2 U16518 ( .A(n15470), .B(n15474), .Z(n17204) );
  HS65_LH_CNIVX3 U16519 ( .A(n13639), .Z(n15741) );
  HS65_LH_NAND3X2 U16520 ( .A(n13654), .B(n15741), .C(n258), .Z(n17202) );
  HS65_LH_NOR2X2 U16521 ( .A(n191), .B(n282), .Z(n15763) );
  HS65_LH_NAND2X2 U16522 ( .A(n15475), .B(n15763), .Z(n15758) );
  HS65_LH_OAI32X2 U16523 ( .A(n15643), .B(n17204), .C(n17202), .D(n13879), .E(
        n15758), .Z(n15708) );
  HS65_LH_NOR2X2 U16527 ( .A(n17246), .B(n17469), .Z(
        \u_DataPath/u_execute/EXALU/N810 ) );
  HS65_LH_OAI212X3 U16529 ( .A(n15718), .B(n15717), .C(n25922), .D(n29559), 
        .E(n17590), .Z(n15727) );
  HS65_LH_IVX2 U16530 ( .A(n15719), .Z(n15725) );
  HS65_LH_AOI21X2 U16531 ( .A(n15722), .B(n15721), .C(n17467), .Z(n15723) );
  HS65_LH_OAI21X2 U16532 ( .A(n15725), .B(n15724), .C(n15723), .Z(n15726) );
  HS65_LH_CBI4I6X2 U16533 ( .A(n15728), .B(n15727), .C(n15726), .D(n17246), 
        .Z(\u_DataPath/u_execute/EXALU/N811 ) );
  HS65_LH_NOR3X1 U16534 ( .A(n11699), .B(n11747), .C(n11723), .Z(n277) );
  HS65_LH_NAND2X2 U16535 ( .A(n12481), .B(n258), .Z(n15732) );
  HS65_LH_NAND2X2 U16536 ( .A(n17204), .B(n15643), .Z(n15740) );
  HS65_LH_NOR3X1 U16537 ( .A(n13654), .B(n15643), .C(n282), .Z(n17203) );
  HS65_LH_NAND2X2 U16538 ( .A(n17203), .B(n15475), .Z(n15731) );
  HS65_LH_NOR2X2 U16539 ( .A(n15474), .B(n17202), .Z(n280) );
  HS65_LH_AOI21X2 U16540 ( .A(n15474), .B(n278), .C(n258), .Z(n15729) );
  HS65_LH_NAND3X2 U16541 ( .A(n13654), .B(n10454), .C(n15729), .Z(n15753) );
  HS65_LH_CNIVX3 U16542 ( .A(n15753), .Z(n17207) );
  HS65_LH_OAI32X2 U16543 ( .A(n17644), .B(n17305), .C(n17440), .D(n17573), .E(
        n17577), .Z(n15730) );
  HS65_LH_NAND3X2 U16545 ( .A(n13890), .B(n11649), .C(n11644), .Z(n15737) );
  HS65_LH_CNIVX3 U16546 ( .A(n15737), .Z(n15756) );
  HS65_LH_CNIVX3 U16547 ( .A(n11649), .Z(n1101) );
  HS65_LH_NAND2X2 U16548 ( .A(n13887), .B(n13885), .Z(n243) );
  HS65_LH_CNIVX3 U16549 ( .A(n243), .Z(n15743) );
  HS65_LH_CNIVX3 U16550 ( .A(n9480), .Z(n1103) );
  HS65_LH_NAND3X2 U16551 ( .A(n196), .B(n15743), .C(n1103), .Z(n15734) );
  HS65_LH_NOR2X2 U16552 ( .A(n15430), .B(n15734), .Z(n15745) );
  HS65_LH_AOI31X2 U16553 ( .A(n15756), .B(n13887), .C(n13885), .D(n15745), .Z(
        n217) );
  HS65_LH_NAND3X2 U16554 ( .A(n196), .B(n15428), .C(n13890), .Z(n15733) );
  HS65_LH_NOR2X2 U16555 ( .A(n15733), .B(n9480), .Z(n15735) );
  HS65_LH_CNIVX3 U16556 ( .A(n15735), .Z(n239) );
  HS65_LH_NOR3X1 U16557 ( .A(n1103), .B(n15428), .C(n15737), .Z(n15755) );
  HS65_LH_NOR2X2 U16558 ( .A(n13885), .B(n15733), .Z(n15746) );
  HS65_LH_NOR2X2 U16559 ( .A(n15755), .B(n15746), .Z(n17210) );
  HS65_LH_NOR2X2 U16560 ( .A(n13890), .B(n15734), .Z(n17209) );
  HS65_LH_AOI21X2 U16561 ( .A(n13885), .B(n15735), .C(n17209), .Z(n15747) );
  HS65_LH_NOR2X2 U16562 ( .A(n13890), .B(n1103), .Z(n242) );
  HS65_LH_NOR2X2 U16563 ( .A(n11649), .B(n11644), .Z(n200) );
  HS65_LH_NAND3X2 U16564 ( .A(n242), .B(n200), .C(n236), .Z(n15738) );
  HS65_LH_NOR2X2 U16565 ( .A(n13887), .B(n15429), .Z(n15736) );
  HS65_LH_MUX21X4 U16566 ( .D0(n15738), .D1(n15737), .S0(n15736), .Z(n15739)
         );
  HS65_LH_NAND3X2 U16567 ( .A(n17210), .B(n15747), .C(n15739), .Z(n198) );
  HS65_LH_NOR2X2 U16568 ( .A(n13639), .B(n258), .Z(n192) );
  HS65_LH_CNIVX3 U16569 ( .A(n15740), .Z(n209) );
  HS65_LH_NAND2X2 U16570 ( .A(n15741), .B(n15474), .Z(n15742) );
  HS65_LH_NOR2X2 U16571 ( .A(n13887), .B(n15430), .Z(n15744) );
  HS65_LH_NOR3X1 U16572 ( .A(n9480), .B(n15744), .C(n15743), .Z(n224) );
  HS65_LH_AOI21X2 U16573 ( .A(n15746), .B(n9480), .C(n15745), .Z(n240) );
  HS65_LH_NAND2X2 U16574 ( .A(n15747), .B(n240), .Z(n225) );
  HS65_LH_CNIVX3 U16575 ( .A(n15748), .Z(n15751) );
  HS65_LH_NOR3X1 U16576 ( .A(n15751), .B(n13639), .C(n15475), .Z(n15749) );
  HS65_LH_NAND3X2 U16577 ( .A(n15749), .B(n191), .C(n258), .Z(n226) );
  HS65_LH_CNIVX3 U16578 ( .A(n17197), .Z(n312) );
  HS65_LH_IVX2 U16579 ( .A(Data_out_fromRAM[30]), .Z(n293) );
  HS65_LH_IVX2 U16580 ( .A(Data_out_fromRAM[27]), .Z(n296) );
  HS65_LH_IVX2 U16581 ( .A(Data_out_fromRAM[25]), .Z(n298) );
  HS65_LH_IVX2 U16582 ( .A(Data_out_fromRAM[24]), .Z(n299) );
  HS65_LH_IVX2 U16583 ( .A(Data_out_fromRAM[18]), .Z(n305) );
  HS65_LH_IVX2 U16584 ( .A(Data_out_fromRAM[28]), .Z(n295) );
  HS65_LH_IVX2 U16585 ( .A(Data_out_fromRAM[20]), .Z(n303) );
  HS65_LH_IVX2 U16586 ( .A(Data_out_fromRAM[23]), .Z(n300) );
  HS65_LH_IVX2 U16587 ( .A(Data_out_fromRAM[19]), .Z(n304) );
  HS65_LH_IVX2 U16588 ( .A(Data_out_fromRAM[17]), .Z(n306) );
  HS65_LH_IVX2 U16589 ( .A(Data_out_fromRAM[21]), .Z(n302) );
  HS65_LH_IVX2 U16590 ( .A(Data_out_fromRAM[16]), .Z(n308) );
  HS65_LH_IVX2 U16591 ( .A(Data_out_fromRAM[29]), .Z(n294) );
  HS65_LH_IVX2 U16592 ( .A(Data_out_fromRAM[26]), .Z(n297) );
  HS65_LH_IVX2 U16593 ( .A(Data_out_fromRAM[22]), .Z(n301) );
  HS65_LH_IVX2 U16594 ( .A(Data_out_fromRAM[31]), .Z(n292) );
  HS65_LH_CNIVX3 U16595 ( .A(n278), .Z(n15757) );
  HS65_LH_NOR2X2 U16596 ( .A(n17202), .B(n15751), .Z(n15761) );
  HS65_LH_NOR3X1 U16598 ( .A(n13879), .B(n15470), .C(n17202), .Z(n15759) );
  HS65_LH_CBI4I6X2 U16599 ( .A(n17630), .B(n17577), .C(n17302), .D(n17296), 
        .Z(n15754) );
  HS65_LH_AOI21X2 U16602 ( .A(n15756), .B(n13885), .C(n15755), .Z(n251) );
  HS65_LH_CNIVX3 U16604 ( .A(n15758), .Z(n15760) );
  HS65_LH_NAND2X2 U16605 ( .A(n13646), .B(n15643), .Z(n17208) );
  HS65_LH_CNIVX3 U16606 ( .A(n17208), .Z(n15762) );
  HS65_LH_AOI21X2 U16607 ( .A(n15763), .B(n15762), .C(n15761), .Z(n230) );
  HS65_LH_NAND3X2 U16608 ( .A(n12324), .B(n15179), .C(n1928), .Z(n15767) );
  HS65_LH_NOR2X5 U16609 ( .A(n15781), .B(n15767), .Z(n16395) );
  HS65_LH_NAND3X2 U16610 ( .A(n12324), .B(n12338), .C(n15179), .Z(n15766) );
  HS65_LH_NOR2X5 U16611 ( .A(n15791), .B(n15766), .Z(n16367) );
  HS65_LH_AOI22X1 U16612 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][0] ), .B(n36264), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][0] ), .D(
        n17431), .Z(n15765) );
  HS65_LH_NAND3X2 U16613 ( .A(n12338), .B(n15179), .C(n14053), .Z(n15773) );
  HS65_LH_NOR2X5 U16614 ( .A(n15773), .B(n15786), .Z(n16368) );
  HS65_LH_NOR2X5 U16615 ( .A(n15791), .B(n15773), .Z(n16393) );
  HS65_LH_AOI22X1 U16616 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][0] ), .B(n17430), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[8][0] ), .D(
        n29554), .Z(n15764) );
  HS65_LH_NAND2X2 U16618 ( .A(n11878), .B(n1913), .Z(n15789) );
  HS65_LH_NOR2X5 U16619 ( .A(n15789), .B(n15766), .Z(n16317) );
  HS65_LH_BFX4 U16620 ( .A(n36385), .Z(n16446) );
  HS65_LH_NOR2X5 U16621 ( .A(n15773), .B(n15781), .Z(n16437) );
  HS65_LH_AO22X4 U16622 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][0] ), .B(n16446), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][0] ), .D(
        n17427), .Z(n15771) );
  HS65_LH_NAND3X2 U16623 ( .A(n15179), .B(n14053), .C(n1928), .Z(n15772) );
  HS65_LH_NOR2X5 U16624 ( .A(n15789), .B(n15767), .Z(n16394) );
  HS65_LH_AO22X4 U16626 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][0] ), .B(n18125), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][0] ), .D(
        n17426), .Z(n15770) );
  HS65_LH_NOR2X5 U16627 ( .A(n15786), .B(n15766), .Z(n16436) );
  HS65_LH_NOR2X5 U16629 ( .A(n15786), .B(n15767), .Z(n16400) );
  HS65_LH_AOI22X1 U16630 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][0] ), .B(n35786), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][0] ), .D(
        n29561), .Z(n15769) );
  HS65_LH_NOR2X5 U16631 ( .A(n15781), .B(n15766), .Z(n16405) );
  HS65_LH_NOR2X5 U16633 ( .A(n15791), .B(n15767), .Z(n16392) );
  HS65_LH_AOI22X1 U16635 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][0] ), .B(n17423), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][0] ), .D(
        n17422), .Z(n15768) );
  HS65_LH_NAND4ABX3 U16636 ( .A(n15771), .B(n15770), .C(n15769), .D(n15768), 
        .Z(n15776) );
  HS65_LH_NOR2X5 U16638 ( .A(n15772), .B(n15786), .Z(n16429) );
  HS65_LH_BFX4 U16639 ( .A(n17421), .Z(n16342) );
  HS65_LH_AOI22X1 U16640 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][0] ), .B(n18122), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][0] ), .D(
        n16342), .Z(n15775) );
  HS65_LH_NOR2X5 U16641 ( .A(n15791), .B(n15772), .Z(n16447) );
  HS65_LH_NOR2X5 U16643 ( .A(n15789), .B(n15773), .Z(n16439) );
  HS65_LH_BFX4 U16644 ( .A(n36958), .Z(n16406) );
  HS65_LH_AOI22X1 U16645 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][0] ), .B(n17420), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[9][0] ), .D(
        n16406), .Z(n15774) );
  HS65_LH_NAND4ABX3 U16646 ( .A(n15777), .B(n15776), .C(n15775), .D(n15774), 
        .Z(n2726) );
  HS65_LH_NAND3X2 U16647 ( .A(n12324), .B(n12370), .C(n1928), .Z(n15780) );
  HS65_LH_NOR2X5 U16648 ( .A(n15791), .B(n15780), .Z(n16411) );
  HS65_LH_NAND3X2 U16649 ( .A(n12370), .B(n12338), .C(n14053), .Z(n15788) );
  HS65_LH_NOR2X5 U16650 ( .A(n15791), .B(n15788), .Z(n16377) );
  HS65_LH_AOI22X1 U16651 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][0] ), .B(n17418), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][0] ), .D(
        n17417), .Z(n15779) );
  HS65_LH_NAND3X2 U16652 ( .A(n12370), .B(n14053), .C(n1928), .Z(n15790) );
  HS65_LH_NOR2X5 U16653 ( .A(n15789), .B(n15790), .Z(n16455) );
  HS65_LH_NOR2X5 U16655 ( .A(n15786), .B(n15790), .Z(n16456) );
  HS65_LH_AOI22X1 U16656 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][0] ), .B(n29606), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][0] ), .D(
        n17415), .Z(n15778) );
  HS65_LH_NAND2X2 U16657 ( .A(n15779), .B(n15778), .Z(n15795) );
  HS65_LH_NOR2X5 U16658 ( .A(n15781), .B(n15788), .Z(n16461) );
  HS65_LH_NAND3X2 U16659 ( .A(n12370), .B(n12324), .C(n12338), .Z(n15787) );
  HS65_LH_NOR2X5 U16660 ( .A(n15791), .B(n15787), .Z(n16351) );
  HS65_LH_BFX4 U16661 ( .A(n36561), .Z(n16474) );
  HS65_LH_AO22X4 U16662 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][0] ), .B(n17414), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][0] ), .D(
        n16474), .Z(n15785) );
  HS65_LH_NOR2X5 U16663 ( .A(n15786), .B(n15780), .Z(n16387) );
  HS65_LH_NOR2X5 U16665 ( .A(n15789), .B(n15780), .Z(n16352) );
  HS65_LH_AO22X4 U16667 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][0] ), .B(n17412), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][0] ), .D(
        n17411), .Z(n15784) );
  HS65_LH_NOR2X5 U16668 ( .A(n15781), .B(n15787), .Z(n16417) );
  HS65_LH_AOI22X1 U16670 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][0] ), .B(n40993), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][0] ), .D(
        n36571), .Z(n15783) );
  HS65_LH_NOR2X5 U16671 ( .A(n15786), .B(n15787), .Z(n16464) );
  HS65_LH_NOR2X5 U16672 ( .A(n15781), .B(n15790), .Z(n16466) );
  HS65_LH_AOI22X1 U16673 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][0] ), .B(n17409), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][0] ), .D(
        n17408), .Z(n15782) );
  HS65_LH_NAND4ABX3 U16674 ( .A(n15785), .B(n15784), .C(n15783), .D(n15782), 
        .Z(n15794) );
  HS65_LH_NOR2X5 U16675 ( .A(n15786), .B(n15788), .Z(n16412) );
  HS65_LH_AOI22X1 U16678 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][0] ), .B(n17407), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][0] ), .D(
        n29602), .Z(n15793) );
  HS65_LH_NOR2X5 U16679 ( .A(n15789), .B(n15788), .Z(n16457) );
  HS65_LH_NOR2X5 U16681 ( .A(n15791), .B(n15790), .Z(n16473) );
  HS65_LH_AOI22X1 U16683 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][0] ), .B(n17406), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[16][0] ), .D(
        n17405), .Z(n15792) );
  HS65_LH_NAND4ABX3 U16684 ( .A(n15795), .B(n15794), .C(n15793), .D(n15792), 
        .Z(n2727) );
  HS65_LH_AOI22X1 U16685 ( .A(n17431), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][1] ), .C(n17426), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][1] ), .Z(
        n15797) );
  HS65_LH_AOI22X1 U16687 ( .A(n29620), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][1] ), .C(n17424), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][1] ), .Z(
        n15796) );
  HS65_LH_AO22X4 U16690 ( .A(n16342), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][1] ), .C(n29543), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][1] ), .Z(
        n15801) );
  HS65_LH_AO22X4 U16691 ( .A(n16446), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][1] ), .C(n17422), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][1] ), .Z(
        n15800) );
  HS65_LH_AOI22X1 U16692 ( .A(n18122), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][1] ), .C(n17423), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][1] ), .Z(
        n15799) );
  HS65_LH_AOI22X1 U16694 ( .A(n36264), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][1] ), .C(n18125), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][1] ), .Z(
        n15798) );
  HS65_LH_NAND4ABX3 U16695 ( .A(n15801), .B(n15800), .C(n15799), .D(n15798), 
        .Z(n15804) );
  HS65_LH_AOI22X1 U16697 ( .A(n17420), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][1] ), .C(n35698), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[8][1] ), .Z(
        n15803) );
  HS65_LH_AOI22X1 U16698 ( .A(n16406), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][1] ), .C(n35786), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][1] ), .Z(
        n15802) );
  HS65_LH_NAND4ABX3 U16699 ( .A(n15805), .B(n15804), .C(n15803), .D(n15802), 
        .Z(n2669) );
  HS65_LH_AOI22X1 U16700 ( .A(n36561), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][1] ), .C(n17409), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][1] ), .Z(
        n15807) );
  HS65_LH_BFX4 U16701 ( .A(n17415), .Z(n16379) );
  HS65_LH_AOI22X1 U16702 ( .A(n16379), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][1] ), .C(n17417), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][1] ), .Z(
        n15806) );
  HS65_LH_NAND2X2 U16703 ( .A(n15807), .B(n15806), .Z(n15815) );
  HS65_LH_AO22X4 U16705 ( .A(n17412), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][1] ), .C(n17408), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][1] ), .Z(
        n15811) );
  HS65_LH_AO22X4 U16706 ( .A(n29606), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][1] ), .C(n29553), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][1] ), .Z(
        n15810) );
  HS65_LH_AOI22X1 U16707 ( .A(n17406), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][1] ), .C(n17407), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][1] ), .Z(
        n15809) );
  HS65_LH_AOI22X1 U16709 ( .A(n17418), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][1] ), .C(n17414), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[27][1] ), .Z(
        n15808) );
  HS65_LH_NAND4ABX3 U16710 ( .A(n15811), .B(n15810), .C(n15809), .D(n15808), 
        .Z(n15814) );
  HS65_LH_AOI22X1 U16711 ( .A(n29602), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][1] ), .C(n40993), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[31][1] ), .Z(
        n15813) );
  HS65_LH_AOI22X1 U16713 ( .A(n17405), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][1] ), .C(n29560), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][1] ), .Z(
        n15812) );
  HS65_LH_NAND4ABX3 U16714 ( .A(n15815), .B(n15814), .C(n15813), .D(n15812), 
        .Z(n2670) );
  HS65_LH_AOI22X1 U16715 ( .A(n36958), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][2] ), .C(n20433), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][2] ), .Z(
        n15817) );
  HS65_LH_AOI22X1 U16716 ( .A(n29603), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][2] ), .C(n29551), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][2] ), .Z(
        n15816) );
  HS65_LH_AO22X4 U16718 ( .A(n18348), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][2] ), .C(n17421), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][2] ), .Z(
        n15821) );
  HS65_LH_AO22X4 U16719 ( .A(n20916), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][2] ), .C(n17424), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][2] ), .Z(
        n15820) );
  HS65_LH_AOI22X1 U16721 ( .A(n17430), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][2] ), .C(n29549), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][2] ), .Z(
        n15819) );
  HS65_LH_AOI22X1 U16723 ( .A(n17427), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][2] ), .C(n17422), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][2] ), .Z(
        n15818) );
  HS65_LH_NAND4ABX3 U16724 ( .A(n15821), .B(n15820), .C(n15819), .D(n15818), 
        .Z(n15824) );
  HS65_LH_AOI22X1 U16725 ( .A(n16446), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][2] ), .C(n20342), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][2] ), .Z(
        n15823) );
  HS65_LH_AOI22X1 U16726 ( .A(n35698), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][2] ), .C(n29542), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][2] ), .Z(
        n15822) );
  HS65_LH_NAND4ABX3 U16727 ( .A(n35671), .B(n35670), .C(n15823), .D(n15822), 
        .Z(n2645) );
  HS65_LH_AOI22X1 U16728 ( .A(n29606), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][2] ), .C(n16474), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][2] ), .Z(
        n15827) );
  HS65_LH_AOI22X1 U16729 ( .A(n29616), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][2] ), .C(n17405), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[16][2] ), .Z(
        n15826) );
  HS65_LH_NAND2X2 U16730 ( .A(n15827), .B(n15826), .Z(n15835) );
  HS65_LH_AO22X4 U16731 ( .A(n16379), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][2] ), .C(n17410), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[31][2] ), .Z(
        n15831) );
  HS65_LH_AO22X4 U16732 ( .A(n18123), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][2] ), .C(n17408), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][2] ), .Z(
        n15830) );
  HS65_LH_AOI22X1 U16733 ( .A(n29622), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][2] ), .C(n17414), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[27][2] ), .Z(
        n15829) );
  HS65_LH_BFX4 U16734 ( .A(n17409), .Z(n16415) );
  HS65_LH_AOI22X1 U16735 ( .A(n29610), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][2] ), .C(n16415), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][2] ), .Z(
        n15828) );
  HS65_LH_NAND4ABX3 U16736 ( .A(n15831), .B(n15830), .C(n15829), .D(n15828), 
        .Z(n15834) );
  HS65_LH_AOI22X1 U16737 ( .A(n40995), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][2] ), .C(n29560), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][2] ), .Z(
        n15833) );
  HS65_LH_AOI22X1 U16739 ( .A(n29552), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][2] ), .C(n29553), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][2] ), .Z(
        n15832) );
  HS65_LH_NAND4ABX3 U16740 ( .A(n15835), .B(n15834), .C(n15833), .D(n15832), 
        .Z(n2646) );
  HS65_LH_AOI22X1 U16741 ( .A(n17423), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][3] ), .C(n17424), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][3] ), .Z(
        n15837) );
  HS65_LH_AOI22X1 U16742 ( .A(n16342), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][3] ), .C(n29554), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[8][3] ), .Z(
        n15836) );
  HS65_LH_NAND2X2 U16743 ( .A(n15837), .B(n15836), .Z(n15845) );
  HS65_LH_AO22X4 U16744 ( .A(n17420), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][3] ), .C(n16406), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[9][3] ), .Z(
        n15841) );
  HS65_LH_AO22X4 U16745 ( .A(n16446), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][3] ), .C(n17422), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][3] ), .Z(
        n15840) );
  HS65_LH_AOI22X1 U16746 ( .A(n18122), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][3] ), .C(n18125), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][3] ), .Z(
        n15839) );
  HS65_LH_AOI22X1 U16747 ( .A(n29549), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][3] ), .C(n17426), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][3] ), .Z(
        n15838) );
  HS65_LH_NAND4ABX3 U16748 ( .A(n15841), .B(n15840), .C(n15839), .D(n15838), 
        .Z(n15844) );
  HS65_LH_AOI22X1 U16750 ( .A(n17430), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][3] ), .C(n17431), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][3] ), .Z(
        n15843) );
  HS65_LH_AOI22X1 U16751 ( .A(n17427), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][3] ), .C(n35786), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][3] ), .Z(
        n15842) );
  HS65_LH_NAND4ABX3 U16752 ( .A(n15845), .B(n15844), .C(n15843), .D(n15842), 
        .Z(n2621) );
  HS65_LH_AOI22X1 U16753 ( .A(n17409), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][3] ), .C(n17410), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[31][3] ), .Z(
        n15847) );
  HS65_LH_AOI22X1 U16754 ( .A(n36759), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][3] ), .C(n17415), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][3] ), .Z(
        n15846) );
  HS65_LH_NAND2X2 U16755 ( .A(n15847), .B(n15846), .Z(n15855) );
  HS65_LH_AO22X4 U16756 ( .A(n18123), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][3] ), .C(n36571), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][3] ), .Z(
        n15851) );
  HS65_LH_AO22X4 U16757 ( .A(n17417), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][3] ), .C(n16474), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][3] ), .Z(
        n15850) );
  HS65_LH_AOI22X1 U16758 ( .A(n17407), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][3] ), .C(n17418), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][3] ), .Z(
        n15849) );
  HS65_LH_AOI22X1 U16759 ( .A(n17406), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][3] ), .C(n17411), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][3] ), .Z(
        n15848) );
  HS65_LH_NAND4ABX3 U16760 ( .A(n15851), .B(n15850), .C(n15849), .D(n15848), 
        .Z(n15854) );
  HS65_LH_AOI22X1 U16761 ( .A(n17414), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][3] ), .C(n40994), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][3] ), .Z(
        n15853) );
  HS65_LH_AOI22X1 U16762 ( .A(n17405), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][3] ), .C(n29622), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][3] ), .Z(
        n15852) );
  HS65_LH_NAND4ABX3 U16763 ( .A(n15855), .B(n15854), .C(n15853), .D(n15852), 
        .Z(n2622) );
  HS65_LH_AOI22X1 U16764 ( .A(n16342), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][4] ), .C(n35698), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[8][4] ), .Z(
        n15857) );
  HS65_LH_AOI22X1 U16765 ( .A(n29603), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][4] ), .C(n18125), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][4] ), .Z(
        n15856) );
  HS65_LH_NAND2X2 U16766 ( .A(n15857), .B(n15856), .Z(n15865) );
  HS65_LH_AO22X4 U16767 ( .A(n16406), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][4] ), .C(n17430), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][4] ), .Z(
        n15861) );
  HS65_LH_AO22X4 U16768 ( .A(n17423), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][4] ), .C(n17422), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][4] ), .Z(
        n15860) );
  HS65_LH_AOI22X1 U16769 ( .A(n29549), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][4] ), .C(n17427), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][4] ), .Z(
        n15859) );
  HS65_LH_AOI22X1 U16770 ( .A(n20916), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][4] ), .C(n18122), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][4] ), .Z(
        n15858) );
  HS65_LH_NAND4ABX3 U16771 ( .A(n15861), .B(n15860), .C(n15859), .D(n15858), 
        .Z(n15864) );
  HS65_LH_AOI22X1 U16772 ( .A(n29551), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][4] ), .C(n16446), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][4] ), .Z(
        n15863) );
  HS65_LH_AOI22X1 U16773 ( .A(n35786), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][4] ), .C(n17424), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][4] ), .Z(
        n15862) );
  HS65_LH_NAND4ABX3 U16774 ( .A(n15865), .B(n15864), .C(n15863), .D(n15862), 
        .Z(n2597) );
  HS65_LH_AOI22X1 U16776 ( .A(n29610), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][4] ), .C(n40995), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][4] ), .Z(
        n15867) );
  HS65_LH_AOI22X1 U16777 ( .A(n29616), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][4] ), .C(n16379), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][4] ), .Z(
        n15866) );
  HS65_LH_NAND2X2 U16778 ( .A(n15867), .B(n15866), .Z(n15875) );
  HS65_LH_AO22X4 U16779 ( .A(n29602), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][4] ), .C(n29560), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][4] ), .Z(
        n15871) );
  HS65_LH_AO22X4 U16780 ( .A(n40994), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][4] ), .C(n17410), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[31][4] ), .Z(
        n15870) );
  HS65_LH_AOI22X1 U16781 ( .A(n29547), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][4] ), .C(n16474), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][4] ), .Z(
        n15869) );
  HS65_LH_AOI22X1 U16782 ( .A(n29622), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][4] ), .C(n29553), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][4] ), .Z(
        n15868) );
  HS65_LH_NAND4ABX3 U16783 ( .A(n15871), .B(n33305), .C(n15869), .D(n15868), 
        .Z(n15874) );
  HS65_LH_AOI22X1 U16784 ( .A(n29606), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][4] ), .C(n16415), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][4] ), .Z(
        n15873) );
  HS65_LH_AOI22X1 U16785 ( .A(n29618), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][4] ), .C(n29552), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][4] ), .Z(
        n15872) );
  HS65_LH_NAND4ABX3 U16786 ( .A(n15875), .B(n15874), .C(n15873), .D(n15872), 
        .Z(n2598) );
  HS65_LH_AOI22X1 U16787 ( .A(n29543), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][5] ), .C(n17424), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][5] ), .Z(
        n15877) );
  HS65_LH_AOI22X1 U16788 ( .A(n17429), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][5] ), .C(n29603), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][5] ), .Z(
        n15876) );
  HS65_LH_AO22X4 U16790 ( .A(n18348), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][5] ), .C(n17426), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][5] ), .Z(
        n15881) );
  HS65_LH_AO22X4 U16791 ( .A(n17423), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][5] ), .C(n29604), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][5] ), .Z(
        n15880) );
  HS65_LH_AOI22X1 U16792 ( .A(n20916), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][5] ), .C(n16342), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][5] ), .Z(
        n15879) );
  HS65_LH_AOI22X1 U16793 ( .A(n29549), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][5] ), .C(n29542), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][5] ), .Z(
        n15878) );
  HS65_LH_NAND4ABX3 U16794 ( .A(n15881), .B(n15880), .C(n15879), .D(n15878), 
        .Z(n15884) );
  HS65_LH_AOI22X1 U16795 ( .A(n16406), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][5] ), .C(n16446), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][5] ), .Z(
        n15883) );
  HS65_LH_AOI22X1 U16796 ( .A(n29620), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][5] ), .C(n20433), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][5] ), .Z(
        n15882) );
  HS65_LH_NAND4ABX3 U16797 ( .A(n36158), .B(n15884), .C(n15883), .D(n15882), 
        .Z(n2573) );
  HS65_LH_AOI22X1 U16798 ( .A(n29606), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][5] ), .C(n16415), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][5] ), .Z(
        n15887) );
  HS65_LH_AOI22X1 U16799 ( .A(n36561), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][5] ), .C(n40993), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[31][5] ), .Z(
        n15886) );
  HS65_LH_NAND2X2 U16800 ( .A(n15887), .B(n15886), .Z(n15895) );
  HS65_LH_AO22X4 U16801 ( .A(n17406), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][5] ), .C(n17414), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[27][5] ), .Z(
        n15891) );
  HS65_LH_AO22X4 U16802 ( .A(n17411), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][5] ), .C(n17408), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][5] ), .Z(
        n15890) );
  HS65_LH_AOI22X1 U16803 ( .A(n18123), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][5] ), .C(n29552), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][5] ), .Z(
        n15889) );
  HS65_LH_AOI22X1 U16804 ( .A(n17415), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][5] ), .C(n29622), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][5] ), .Z(
        n15888) );
  HS65_LH_NAND4ABX3 U16805 ( .A(n15891), .B(n15890), .C(n15889), .D(n15888), 
        .Z(n15894) );
  HS65_LH_AOI22X1 U16806 ( .A(n17405), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][5] ), .C(n29560), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][5] ), .Z(
        n15893) );
  HS65_LH_AOI22X1 U16807 ( .A(n29610), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][5] ), .C(n40995), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][5] ), .Z(
        n15892) );
  HS65_LH_AOI22X1 U16809 ( .A(n36958), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][6] ), .C(n29603), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][6] ), .Z(
        n15897) );
  HS65_LH_AOI22X1 U16810 ( .A(n29551), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][6] ), .C(n29561), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][6] ), .Z(
        n15896) );
  HS65_LH_AO22X4 U16812 ( .A(n18348), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][6] ), .C(n29543), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][6] ), .Z(
        n15901) );
  HS65_LH_AO22X4 U16813 ( .A(n16342), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][6] ), .C(n29604), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][6] ), .Z(
        n15900) );
  HS65_LH_AOI22X1 U16814 ( .A(n20916), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][6] ), .C(n36385), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][6] ), .Z(
        n15899) );
  HS65_LH_AOI22X1 U16815 ( .A(n29554), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][6] ), .C(n20342), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][6] ), .Z(
        n15898) );
  HS65_LH_NAND4ABX3 U16816 ( .A(n15901), .B(n15900), .C(n15899), .D(n15898), 
        .Z(n15904) );
  HS65_LH_AOI22X1 U16817 ( .A(n29549), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][6] ), .C(n29620), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][6] ), .Z(
        n15903) );
  HS65_LH_AOI22X1 U16818 ( .A(n29542), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][6] ), .C(n20433), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][6] ), .Z(
        n15902) );
  HS65_LH_NAND4ABX3 U16819 ( .A(n35789), .B(n15904), .C(n15903), .D(n15902), 
        .Z(n2549) );
  HS65_LH_AOI22X1 U16820 ( .A(n17412), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][6] ), .C(n40994), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][6] ), .Z(
        n15907) );
  HS65_LH_AOI22X1 U16821 ( .A(n29616), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][6] ), .C(n29553), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][6] ), .Z(
        n15906) );
  HS65_LH_AO22X4 U16823 ( .A(n17405), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][6] ), .C(n17417), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][6] ), .Z(
        n15911) );
  HS65_LH_AO22X4 U16824 ( .A(n36759), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][6] ), .C(n29560), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][6] ), .Z(
        n15910) );
  HS65_LH_AOI22X1 U16825 ( .A(n29602), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][6] ), .C(n16415), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][6] ), .Z(
        n15909) );
  HS65_LH_AOI22X1 U16826 ( .A(n29610), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][6] ), .C(n29552), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][6] ), .Z(
        n15908) );
  HS65_LH_NAND4ABX3 U16827 ( .A(n15911), .B(n15910), .C(n15909), .D(n15908), 
        .Z(n15914) );
  HS65_LH_AOI22X1 U16828 ( .A(n16379), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][6] ), .C(n16474), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][6] ), .Z(
        n15913) );
  HS65_LH_AOI22X1 U16829 ( .A(n29547), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][6] ), .C(n40993), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[31][6] ), .Z(
        n15912) );
  HS65_LH_NAND4ABX3 U16830 ( .A(n15915), .B(n15914), .C(n15913), .D(n15912), 
        .Z(n2550) );
  HS65_LH_AOI22X1 U16831 ( .A(n17429), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][7] ), .C(n17423), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][7] ), .Z(
        n15917) );
  HS65_LH_AOI22X1 U16832 ( .A(n36958), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][7] ), .C(n17422), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][7] ), .Z(
        n15916) );
  HS65_LH_AO22X4 U16834 ( .A(n18122), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][7] ), .C(n18125), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][7] ), .Z(
        n15921) );
  HS65_LH_AO22X4 U16835 ( .A(n16342), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][7] ), .C(n17432), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][7] ), .Z(
        n15920) );
  HS65_LH_AOI22X1 U16836 ( .A(n17431), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][7] ), .C(n17425), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][7] ), .Z(
        n15919) );
  HS65_LH_AOI22X1 U16837 ( .A(n16446), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][7] ), .C(n17427), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][7] ), .Z(
        n15918) );
  HS65_LH_NAND4ABX3 U16838 ( .A(n15921), .B(n15920), .C(n15919), .D(n15918), 
        .Z(n15924) );
  HS65_LH_AOI22X1 U16839 ( .A(n17430), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][7] ), .C(n17424), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][7] ), .Z(
        n15923) );
  HS65_LH_AOI22X1 U16840 ( .A(n17420), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][7] ), .C(n17426), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][7] ), .Z(
        n15922) );
  HS65_LH_NAND4ABX3 U16841 ( .A(n15925), .B(n15924), .C(n15923), .D(n15922), 
        .Z(n2525) );
  HS65_LH_AOI22X1 U16842 ( .A(n17418), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][7] ), .C(n16415), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][7] ), .Z(
        n15927) );
  HS65_LH_AOI22X1 U16843 ( .A(n17412), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][7] ), .C(n17411), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][7] ), .Z(
        n15926) );
  HS65_LH_NAND2X2 U16844 ( .A(n15927), .B(n15926), .Z(n15935) );
  HS65_LH_AO22X4 U16845 ( .A(n18123), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][7] ), .C(n17408), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][7] ), .Z(
        n15931) );
  HS65_LH_AO22X4 U16846 ( .A(n17405), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][7] ), .C(n16474), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][7] ), .Z(
        n15930) );
  HS65_LH_AOI22X1 U16847 ( .A(n36759), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][7] ), .C(n18126), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][7] ), .Z(
        n15929) );
  HS65_LH_AOI22X1 U16848 ( .A(n17415), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][7] ), .C(n40993), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[31][7] ), .Z(
        n15928) );
  HS65_LH_NAND4ABX3 U16849 ( .A(n15931), .B(n15930), .C(n15929), .D(n15928), 
        .Z(n15934) );
  HS65_LH_AOI22X1 U16850 ( .A(n17406), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][7] ), .C(n40995), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][7] ), .Z(
        n15933) );
  HS65_LH_AOI22X1 U16851 ( .A(n29610), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][7] ), .C(n29547), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[27][7] ), .Z(
        n15932) );
  HS65_LH_AOI22X1 U16853 ( .A(n17432), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][8] ), .C(n18125), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][8] ), .Z(
        n15937) );
  HS65_LH_AOI22X1 U16854 ( .A(n16406), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][8] ), .C(n17424), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][8] ), .Z(
        n15936) );
  HS65_LH_NAND2X2 U16855 ( .A(n15937), .B(n15936), .Z(n15945) );
  HS65_LH_AO22X4 U16856 ( .A(n17430), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][8] ), .C(n17425), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][8] ), .Z(
        n15941) );
  HS65_LH_AO22X4 U16857 ( .A(n17420), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][8] ), .C(n17427), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][8] ), .Z(
        n15940) );
  HS65_LH_AOI22X1 U16858 ( .A(n16342), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][8] ), .C(n17431), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][8] ), .Z(
        n15939) );
  HS65_LH_AOI22X1 U16859 ( .A(n17426), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][8] ), .C(n17422), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][8] ), .Z(
        n15938) );
  HS65_LH_NAND4ABX3 U16860 ( .A(n15941), .B(n15940), .C(n15939), .D(n15938), 
        .Z(n15944) );
  HS65_LH_AOI22X1 U16861 ( .A(n16446), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][8] ), .C(n20342), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][8] ), .Z(
        n15943) );
  HS65_LH_AOI22X1 U16862 ( .A(n18122), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][8] ), .C(n17429), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[8][8] ), .Z(
        n15942) );
  HS65_LH_NAND4ABX3 U16863 ( .A(n15945), .B(n15944), .C(n15943), .D(n36755), 
        .Z(n2501) );
  HS65_LH_AOI22X1 U16864 ( .A(n17405), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][8] ), .C(n17417), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][8] ), .Z(
        n15947) );
  HS65_LH_AOI22X1 U16865 ( .A(n17409), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][8] ), .C(n18126), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][8] ), .Z(
        n15946) );
  HS65_LH_NAND2X2 U16866 ( .A(n15947), .B(n15946), .Z(n15955) );
  HS65_LH_AO22X4 U16867 ( .A(n18123), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][8] ), .C(n17408), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][8] ), .Z(
        n15951) );
  HS65_LH_AO22X4 U16868 ( .A(n17418), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][8] ), .C(n17411), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][8] ), .Z(
        n15950) );
  HS65_LH_AOI22X1 U16869 ( .A(n17407), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][8] ), .C(n16474), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][8] ), .Z(
        n15949) );
  HS65_LH_AOI22X1 U16870 ( .A(n17406), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][8] ), .C(n17415), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][8] ), .Z(
        n15948) );
  HS65_LH_NAND4ABX3 U16871 ( .A(n15951), .B(n15950), .C(n15949), .D(n15948), 
        .Z(n15954) );
  HS65_LH_AOI22X1 U16872 ( .A(n17412), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][8] ), .C(n17414), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[27][8] ), .Z(
        n15953) );
  HS65_LH_AOI22X1 U16873 ( .A(n36759), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][8] ), .C(n40993), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[31][8] ), .Z(
        n15952) );
  HS65_LH_AOI22X1 U16875 ( .A(n29603), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][9] ), .C(n17422), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][9] ), .Z(
        n15957) );
  HS65_LH_AOI22X1 U16876 ( .A(n20916), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][9] ), .C(n18348), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][9] ), .Z(
        n15956) );
  HS65_LH_NAND2X2 U16877 ( .A(n15957), .B(n15956), .Z(n15965) );
  HS65_LH_AO22X4 U16878 ( .A(n16342), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][9] ), .C(n17427), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][9] ), .Z(
        n15961) );
  HS65_LH_AO22X4 U16879 ( .A(n17423), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][9] ), .C(n29561), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][9] ), .Z(
        n15960) );
  HS65_LH_AOI22X1 U16880 ( .A(n29551), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][9] ), .C(n36385), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][9] ), .Z(
        n15959) );
  HS65_LH_AOI22X1 U16881 ( .A(n29554), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][9] ), .C(n36264), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][9] ), .Z(
        n15958) );
  HS65_LH_NAND4ABX3 U16882 ( .A(n15961), .B(n15960), .C(n15959), .D(n15958), 
        .Z(n15964) );
  HS65_LH_AOI22X1 U16883 ( .A(n16406), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][9] ), .C(n20433), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][9] ), .Z(
        n15963) );
  HS65_LH_AOI22X1 U16884 ( .A(n17430), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][9] ), .C(n18125), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][9] ), .Z(
        n15962) );
  HS65_LH_NAND4ABX3 U16885 ( .A(n15965), .B(n15964), .C(n15963), .D(n15962), 
        .Z(n2477) );
  HS65_LH_AOI22X1 U16886 ( .A(n18123), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][9] ), .C(n17417), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][9] ), .Z(
        n15967) );
  HS65_LH_AOI22X1 U16887 ( .A(n29618), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][9] ), .C(n29606), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[17][9] ), .Z(
        n15966) );
  HS65_LH_NAND2X2 U16888 ( .A(n15967), .B(n15966), .Z(n15975) );
  HS65_LH_AO22X4 U16889 ( .A(n16379), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][9] ), .C(n17410), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[31][9] ), .Z(
        n15971) );
  HS65_LH_AO22X4 U16890 ( .A(n36561), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][9] ), .C(n36571), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][9] ), .Z(
        n15970) );
  HS65_LH_AOI22X1 U16891 ( .A(n29610), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][9] ), .C(n17408), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][9] ), .Z(
        n15969) );
  HS65_LH_AOI22X1 U16892 ( .A(n29616), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][9] ), .C(n16415), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][9] ), .Z(
        n15968) );
  HS65_LH_NAND4ABX3 U16893 ( .A(n15971), .B(n15970), .C(n15969), .D(n15968), 
        .Z(n15974) );
  HS65_LH_AOI22X1 U16894 ( .A(n29553), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][9] ), .C(n17414), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[27][9] ), .Z(
        n15973) );
  HS65_LH_AOI22X1 U16895 ( .A(n17418), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][9] ), .C(n29622), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][9] ), .Z(
        n15972) );
  HS65_LH_NAND4ABX3 U16896 ( .A(n15975), .B(n15974), .C(n15973), .D(n15972), 
        .Z(n2478) );
  HS65_LH_AOI22X1 U16897 ( .A(n20916), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][10] ), .C(n17427), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][10] ), .Z(
        n15977) );
  HS65_LH_AOI22X1 U16898 ( .A(n17430), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][10] ), .C(n17428), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][10] ), .Z(n15976)
         );
  HS65_LH_AO22X4 U16900 ( .A(n17429), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][10] ), .C(n29561), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][10] ), .Z(
        n15981) );
  HS65_LH_AO22X4 U16901 ( .A(n17423), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][10] ), .C(n17425), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][10] ), .Z(n15980)
         );
  HS65_LH_AOI22X1 U16902 ( .A(n17431), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][10] ), .C(n18125), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][10] ), .Z(n15979) );
  HS65_LH_AOI22X1 U16903 ( .A(n18122), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][10] ), .C(n16342), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][10] ), .Z(
        n15978) );
  HS65_LH_NAND4ABX3 U16904 ( .A(n15981), .B(n15980), .C(n15979), .D(n15978), 
        .Z(n15984) );
  HS65_LH_AOI22X1 U16905 ( .A(n17432), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][10] ), .C(n17422), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][10] ), .Z(
        n15983) );
  HS65_LH_AOI22X1 U16906 ( .A(n16406), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][10] ), .C(n29551), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][10] ), .Z(
        n15982) );
  HS65_LH_NAND4ABX3 U16907 ( .A(n15985), .B(n15984), .C(n15983), .D(n15982), 
        .Z(n2453) );
  HS65_LH_AOI22X1 U16908 ( .A(n17418), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][10] ), .C(n16415), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][10] ), .Z(n15987)
         );
  HS65_LH_AOI22X1 U16909 ( .A(n17406), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][10] ), .C(n17410), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[31][10] ), .Z(n15986)
         );
  HS65_LH_NAND2X2 U16910 ( .A(n15987), .B(n15986), .Z(n15995) );
  HS65_LH_AO22X4 U16911 ( .A(n17408), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][10] ), .C(n18126), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][10] ), .Z(n15991)
         );
  HS65_LH_AO22X4 U16912 ( .A(n17417), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][10] ), .C(n17413), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][10] ), .Z(n15990)
         );
  HS65_LH_AOI22X1 U16913 ( .A(n17405), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][10] ), .C(n18123), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][10] ), .Z(n15989)
         );
  HS65_LH_AOI22X1 U16914 ( .A(n17415), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][10] ), .C(n17414), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[27][10] ), .Z(n15988)
         );
  HS65_LH_NAND4ABX3 U16915 ( .A(n15991), .B(n15990), .C(n15989), .D(n15988), 
        .Z(n15994) );
  HS65_LH_AOI22X1 U16916 ( .A(n17407), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][10] ), .C(n17416), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[17][10] ), .Z(n15993)
         );
  HS65_LH_AOI22X1 U16917 ( .A(n17412), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][10] ), .C(n29553), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][10] ), .Z(n15992)
         );
  HS65_LH_NAND4ABX3 U16918 ( .A(n15995), .B(n15994), .C(n15993), .D(n15992), 
        .Z(n2454) );
  HS65_LH_AOI22X1 U16919 ( .A(n29554), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][11] ), .C(n16446), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][11] ), .Z(
        n15997) );
  HS65_LH_AOI22X1 U16920 ( .A(n18122), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][11] ), .C(n17422), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][11] ), .Z(
        n15996) );
  HS65_LH_NAND2X2 U16921 ( .A(n15997), .B(n15996), .Z(n16005) );
  HS65_LH_AO22X4 U16922 ( .A(n16406), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][11] ), .C(n17427), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][11] ), .Z(
        n16001) );
  HS65_LH_AO22X4 U16923 ( .A(n16342), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][11] ), .C(n17431), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][11] ), .Z(
        n16000) );
  HS65_LH_AOI22X1 U16924 ( .A(n20916), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][11] ), .C(n17425), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][11] ), .Z(
        n15999) );
  HS65_LH_AOI22X1 U16925 ( .A(n29543), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][11] ), .C(n17424), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][11] ), .Z(n15998) );
  HS65_LH_NAND4ABX3 U16926 ( .A(n16001), .B(n16000), .C(n15999), .D(n15998), 
        .Z(n16004) );
  HS65_LH_AOI22X1 U16927 ( .A(n17432), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][11] ), .C(n20342), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][11] ), .Z(
        n16003) );
  HS65_LH_AOI22X1 U16928 ( .A(n29542), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][11] ), .C(n17426), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][11] ), .Z(
        n16002) );
  HS65_LH_NAND4ABX3 U16929 ( .A(n16005), .B(n16004), .C(n16003), .D(n16002), 
        .Z(n2429) );
  HS65_LH_AOI22X1 U16930 ( .A(n17411), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][11] ), .C(n36571), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][11] ), .Z(n16007)
         );
  HS65_LH_AOI22X1 U16931 ( .A(n17407), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][11] ), .C(n17417), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][11] ), .Z(n16006)
         );
  HS65_LH_NAND2X2 U16932 ( .A(n16007), .B(n16006), .Z(n16015) );
  HS65_LH_AO22X4 U16933 ( .A(n16379), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][11] ), .C(n16415), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][11] ), .Z(n16011)
         );
  HS65_LH_AO22X4 U16934 ( .A(n17414), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][11] ), .C(n36561), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][11] ), .Z(n16010)
         );
  HS65_LH_AOI22X1 U16935 ( .A(n17418), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][11] ), .C(n29622), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][11] ), .Z(n16009)
         );
  HS65_LH_AOI22X1 U16936 ( .A(n29618), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][11] ), .C(n17410), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[31][11] ), .Z(n16008)
         );
  HS65_LH_AOI22X1 U16939 ( .A(n29616), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][11] ), .C(n36759), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[17][11] ), .Z(n16012)
         );
  HS65_LH_NAND4ABX3 U16940 ( .A(n16015), .B(n36488), .C(n36563), .D(n16012), 
        .Z(n2430) );
  HS65_LH_AOI22X1 U16941 ( .A(n29554), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][12] ), .C(n18125), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][12] ), .Z(
        n16017) );
  HS65_LH_AOI22X1 U16942 ( .A(n17430), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][12] ), .C(n16446), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][12] ), .Z(n16016)
         );
  HS65_LH_NAND2X2 U16943 ( .A(n16017), .B(n16016), .Z(n16025) );
  HS65_LH_AO22X4 U16944 ( .A(n20916), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][12] ), .C(n17432), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][12] ), .Z(
        n16021) );
  HS65_LH_AO22X4 U16945 ( .A(n17423), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][12] ), .C(n17424), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][12] ), .Z(n16020) );
  HS65_LH_AOI22X1 U16946 ( .A(n18122), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][12] ), .C(n17426), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][12] ), .Z(
        n16019) );
  HS65_LH_AOI22X1 U16947 ( .A(n16406), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][12] ), .C(n17422), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][12] ), .Z(
        n16018) );
  HS65_LH_NAND4ABX3 U16948 ( .A(n16021), .B(n16020), .C(n16019), .D(n16018), 
        .Z(n16024) );
  HS65_LH_AOI22X1 U16949 ( .A(n17431), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][12] ), .C(n17425), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][12] ), .Z(n16023)
         );
  HS65_LH_AOI22X1 U16950 ( .A(n17421), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][12] ), .C(n17427), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][12] ), .Z(
        n16022) );
  HS65_LH_NAND4ABX3 U16951 ( .A(n16025), .B(n16024), .C(n16023), .D(n36478), 
        .Z(n2405) );
  HS65_LH_AOI22X1 U16952 ( .A(n17411), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][12] ), .C(n36571), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][12] ), .Z(n16027)
         );
  HS65_LH_AOI22X1 U16953 ( .A(n40995), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][12] ), .C(n40994), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][12] ), .Z(n16026)
         );
  HS65_LH_NAND2X2 U16954 ( .A(n16027), .B(n16026), .Z(n16035) );
  HS65_LH_AO22X4 U16955 ( .A(n17406), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][12] ), .C(n16379), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][12] ), .Z(n16031)
         );
  HS65_LH_AO22X4 U16956 ( .A(n17407), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][12] ), .C(n18123), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][12] ), .Z(n16030)
         );
  HS65_LH_AOI22X1 U16957 ( .A(n29618), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][12] ), .C(n16474), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][12] ), .Z(n16029)
         );
  HS65_LH_AOI22X1 U16958 ( .A(n29606), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][12] ), .C(n40993), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[31][12] ), .Z(n16028)
         );
  HS65_LH_NAND4ABX3 U16959 ( .A(n16031), .B(n16030), .C(n16029), .D(n16028), 
        .Z(n16034) );
  HS65_LH_AOI22X1 U16960 ( .A(n17418), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][12] ), .C(n29622), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][12] ), .Z(n16033)
         );
  HS65_LH_AOI22X1 U16961 ( .A(n17414), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][12] ), .C(n16415), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][12] ), .Z(n16032)
         );
  HS65_LH_NAND4ABX3 U16962 ( .A(n16035), .B(n16034), .C(n36469), .D(n36472), 
        .Z(n2406) );
  HS65_LH_AOI22X1 U16963 ( .A(n29551), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][13] ), .C(n17427), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][13] ), .Z(
        n16037) );
  HS65_LH_AOI22X1 U16964 ( .A(n17429), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][13] ), .C(n20342), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][13] ), .Z(
        n16036) );
  HS65_LH_AO22X4 U16966 ( .A(n17430), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][13] ), .C(n20433), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][13] ), .Z(n16041)
         );
  HS65_LH_AO22X4 U16967 ( .A(n29542), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][13] ), .C(n17424), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][13] ), .Z(
        n16040) );
  HS65_LH_AOI22X1 U16968 ( .A(n29549), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][13] ), .C(n17428), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][13] ), .Z(
        n16039) );
  HS65_LH_AOI22X1 U16969 ( .A(n18122), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][13] ), .C(n29603), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][13] ), .Z(
        n16038) );
  HS65_LH_NAND4ABX3 U16970 ( .A(n16041), .B(n16040), .C(n16039), .D(n16038), 
        .Z(n16044) );
  HS65_LH_AOI22X1 U16971 ( .A(n16406), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][13] ), .C(n16342), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][13] ), .Z(
        n16043) );
  HS65_LH_AOI22X1 U16972 ( .A(n20916), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][13] ), .C(n17422), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][13] ), .Z(
        n16042) );
  HS65_LH_NAND4ABX3 U16973 ( .A(n29538), .B(n16044), .C(n16043), .D(n36646), 
        .Z(n2381) );
  HS65_LH_AOI22X1 U16974 ( .A(n29610), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][13] ), .C(n29602), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][13] ), .Z(n16047)
         );
  HS65_LH_AOI22X1 U16975 ( .A(n17411), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][13] ), .C(n17414), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[27][13] ), .Z(n16046)
         );
  HS65_LH_AO22X4 U16977 ( .A(n17406), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][13] ), .C(n17408), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][13] ), .Z(n16051)
         );
  HS65_LH_AO22X4 U16978 ( .A(n17413), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][13] ), .C(n17409), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][13] ), .Z(n16050)
         );
  HS65_LH_AOI22X1 U16979 ( .A(n17412), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][13] ), .C(n40993), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[31][13] ), .Z(n16049)
         );
  HS65_LH_AOI22X1 U16980 ( .A(n29618), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][13] ), .C(n16379), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][13] ), .Z(n16048)
         );
  HS65_LH_NAND4ABX3 U16981 ( .A(n16051), .B(n16050), .C(n16049), .D(n16048), 
        .Z(n16054) );
  HS65_LH_AOI22X1 U16982 ( .A(n40995), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][13] ), .C(n36571), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][13] ), .Z(n16053)
         );
  HS65_LH_AOI22X1 U16983 ( .A(n36759), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][13] ), .C(n29552), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][13] ), .Z(n16052)
         );
  HS65_LH_NAND4ABX3 U16984 ( .A(n16055), .B(n16054), .C(n36650), .D(n16052), 
        .Z(n2382) );
  HS65_LH_AOI22X1 U16985 ( .A(n35698), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][14] ), .C(n17422), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][14] ), .Z(
        n16057) );
  HS65_LH_AOI22X1 U16986 ( .A(n36385), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][14] ), .C(n29561), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][14] ), .Z(n16056) );
  HS65_LH_NAND2X2 U16987 ( .A(n16057), .B(n16056), .Z(n16065) );
  HS65_LH_AO22X4 U16988 ( .A(n16342), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][14] ), .C(n20433), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][14] ), .Z(
        n16061) );
  HS65_LH_AO22X4 U16989 ( .A(n29603), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][14] ), .C(n17423), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][14] ), .Z(n16060)
         );
  HS65_LH_AOI22X1 U16990 ( .A(n17420), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][14] ), .C(n17427), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][14] ), .Z(
        n16059) );
  HS65_LH_AOI22X1 U16991 ( .A(n36264), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][14] ), .C(n18125), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][14] ), .Z(
        n16058) );
  HS65_LH_NAND4ABX3 U16992 ( .A(n16061), .B(n16060), .C(n16059), .D(n16058), 
        .Z(n16064) );
  HS65_LH_AOI22X1 U16993 ( .A(n29543), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][14] ), .C(n17426), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][14] ), .Z(n16063) );
  HS65_LH_AOI22X1 U16994 ( .A(n16406), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][14] ), .C(n18348), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][14] ), .Z(
        n16062) );
  HS65_LH_NAND4ABX3 U16995 ( .A(n16065), .B(n16064), .C(n16063), .D(n16062), 
        .Z(n2357) );
  HS65_LH_AOI22X1 U16996 ( .A(n17417), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][14] ), .C(n29547), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[27][14] ), .Z(n16067)
         );
  HS65_LH_AOI22X1 U16997 ( .A(n17407), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][14] ), .C(n17408), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][14] ), .Z(n16066)
         );
  HS65_LH_AO22X4 U16999 ( .A(n16379), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][14] ), .C(n17411), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][14] ), .Z(n16071)
         );
  HS65_LH_AO22X4 U17000 ( .A(n36759), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][14] ), .C(n16415), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][14] ), .Z(n16070)
         );
  HS65_LH_AOI22X1 U17001 ( .A(n29618), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][14] ), .C(n29560), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][14] ), .Z(n16069)
         );
  HS65_LH_AOI22X1 U17002 ( .A(n29552), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][14] ), .C(n16474), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][14] ), .Z(n16068)
         );
  HS65_LH_NAND4ABX3 U17003 ( .A(n16071), .B(n16070), .C(n16069), .D(n16068), 
        .Z(n16074) );
  HS65_LH_AOI22X1 U17004 ( .A(n29616), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][14] ), .C(n29602), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][14] ), .Z(n16073)
         );
  HS65_LH_AOI22X1 U17005 ( .A(n17412), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][14] ), .C(n17410), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[31][14] ), .Z(n16072)
         );
  HS65_LH_NAND4ABX3 U17006 ( .A(n16075), .B(n16074), .C(n16073), .D(n16072), 
        .Z(n2358) );
  HS65_LH_AOI22X1 U17007 ( .A(n17421), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][15] ), .C(n17432), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][15] ), .Z(
        n16077) );
  HS65_LH_AOI22X1 U17008 ( .A(n18122), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][15] ), .C(n29551), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][15] ), .Z(
        n16076) );
  HS65_LH_NAND2X2 U17009 ( .A(n16077), .B(n16076), .Z(n16085) );
  HS65_LH_AO22X4 U17010 ( .A(n17429), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][15] ), .C(n17431), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][15] ), .Z(
        n16081) );
  HS65_LH_AO22X4 U17011 ( .A(n17430), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][15] ), .C(n20342), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][15] ), .Z(n16080)
         );
  HS65_LH_AOI22X1 U17012 ( .A(n17427), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][15] ), .C(n29561), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][15] ), .Z(n16079) );
  HS65_LH_AOI22X1 U17013 ( .A(n16406), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][15] ), .C(n29542), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][15] ), .Z(
        n16078) );
  HS65_LH_NAND4ABX3 U17014 ( .A(n16081), .B(n16080), .C(n16079), .D(n16078), 
        .Z(n16084) );
  HS65_LH_AOI22X1 U17015 ( .A(n36385), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][15] ), .C(n29604), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][15] ), .Z(n16083) );
  HS65_LH_AOI22X1 U17016 ( .A(n17420), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][15] ), .C(n20433), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][15] ), .Z(
        n16082) );
  HS65_LH_NAND4ABX3 U17017 ( .A(n16085), .B(n16084), .C(n36387), .D(n16082), 
        .Z(n2333) );
  HS65_LH_AOI22X1 U17018 ( .A(n16379), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][15] ), .C(n29622), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][15] ), .Z(n16087)
         );
  HS65_LH_AOI22X1 U17019 ( .A(n29552), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][15] ), .C(n36571), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][15] ), .Z(n16086)
         );
  HS65_LH_NAND2X2 U17020 ( .A(n16087), .B(n16086), .Z(n16095) );
  HS65_LH_AO22X4 U17021 ( .A(n17417), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][15] ), .C(n40993), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[31][15] ), .Z(n16091)
         );
  HS65_LH_AO22X4 U17022 ( .A(n29602), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][15] ), .C(n17408), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][15] ), .Z(n16090)
         );
  HS65_LH_AOI22X1 U17023 ( .A(n36759), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][15] ), .C(n17409), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][15] ), .Z(n16089)
         );
  HS65_LH_AOI22X1 U17024 ( .A(n29618), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][15] ), .C(n29610), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][15] ), .Z(n16088)
         );
  HS65_LH_NAND4ABX3 U17025 ( .A(n16091), .B(n16090), .C(n16089), .D(n16088), 
        .Z(n16094) );
  HS65_LH_AOI22X1 U17026 ( .A(n29616), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][15] ), .C(n29553), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][15] ), .Z(n16093)
         );
  HS65_LH_AOI22X1 U17027 ( .A(n17414), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][15] ), .C(n16474), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][15] ), .Z(n16092)
         );
  HS65_LH_NAND4ABX3 U17028 ( .A(n16095), .B(n16094), .C(n16093), .D(n16092), 
        .Z(n2334) );
  HS65_LH_AOI22X1 U17029 ( .A(n17421), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][16] ), .C(n29554), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[8][16] ), .Z(
        n16097) );
  HS65_LH_AOI22X1 U17030 ( .A(n29542), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][16] ), .C(n29604), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][16] ), .Z(
        n16096) );
  HS65_LH_AO22X4 U17032 ( .A(n29551), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][16] ), .C(n16446), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][16] ), .Z(
        n16101) );
  HS65_LH_AO22X4 U17033 ( .A(n29549), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][16] ), .C(n20433), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][16] ), .Z(
        n16100) );
  HS65_LH_AOI22X1 U17034 ( .A(n17420), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][16] ), .C(n16406), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[9][16] ), .Z(
        n16099) );
  HS65_LH_AOI22X1 U17035 ( .A(n18348), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][16] ), .C(n29603), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][16] ), .Z(
        n16098) );
  HS65_LH_NAND4ABX3 U17036 ( .A(n16101), .B(n16100), .C(n16099), .D(n16098), 
        .Z(n16104) );
  HS65_LH_AOI22X1 U17037 ( .A(n29620), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][16] ), .C(n29561), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][16] ), .Z(n16103) );
  HS65_LH_AOI22X1 U17038 ( .A(n29543), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][16] ), .C(n20342), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][16] ), .Z(n16102)
         );
  HS65_LH_NAND4ABX3 U17039 ( .A(n35839), .B(n16104), .C(n16103), .D(n16102), 
        .Z(n2309) );
  HS65_LH_AOI22X1 U17040 ( .A(n17409), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][16] ), .C(n17408), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][16] ), .Z(n16107)
         );
  HS65_LH_AOI22X1 U17041 ( .A(n17407), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][16] ), .C(n29622), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][16] ), .Z(n16106)
         );
  HS65_LH_AO22X4 U17043 ( .A(n17411), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][16] ), .C(n36571), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][16] ), .Z(n16111)
         );
  HS65_LH_AO22X4 U17044 ( .A(n17406), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][16] ), .C(n17417), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][16] ), .Z(n16110)
         );
  HS65_LH_AOI22X1 U17045 ( .A(n17405), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][16] ), .C(n16379), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][16] ), .Z(n16109)
         );
  HS65_LH_AOI22X1 U17046 ( .A(n29606), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][16] ), .C(n36561), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][16] ), .Z(n16108)
         );
  HS65_LH_NAND4ABX3 U17047 ( .A(n16111), .B(n16110), .C(n16109), .D(n16108), 
        .Z(n16114) );
  HS65_LH_AOI22X1 U17048 ( .A(n18123), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][16] ), .C(n29547), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[27][16] ), .Z(n16113)
         );
  HS65_LH_AOI22X1 U17049 ( .A(n29552), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][16] ), .C(n17410), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[31][16] ), .Z(n16112)
         );
  HS65_LH_AOI22X1 U17051 ( .A(n29542), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][17] ), .C(n36385), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][17] ), .Z(
        n16117) );
  HS65_LH_AOI22X1 U17052 ( .A(n29554), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][17] ), .C(n29620), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][17] ), .Z(
        n16116) );
  HS65_LH_NAND2X2 U17053 ( .A(n16117), .B(n16116), .Z(n16125) );
  HS65_LH_AO22X4 U17054 ( .A(n17430), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][17] ), .C(n17431), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][17] ), .Z(n16121)
         );
  HS65_LH_AO22X4 U17055 ( .A(n16342), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][17] ), .C(n29561), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][17] ), .Z(
        n16120) );
  HS65_LH_AOI22X1 U17056 ( .A(n17420), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][17] ), .C(n36958), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[9][17] ), .Z(
        n16119) );
  HS65_LH_AOI22X1 U17057 ( .A(n18348), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][17] ), .C(n20433), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][17] ), .Z(
        n16118) );
  HS65_LH_NAND4ABX3 U17058 ( .A(n16121), .B(n16120), .C(n16119), .D(n16118), 
        .Z(n16124) );
  HS65_LH_AOI22X1 U17059 ( .A(n36264), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][17] ), .C(n20342), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][17] ), .Z(
        n16123) );
  HS65_LH_AOI22X1 U17060 ( .A(n29551), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][17] ), .C(n29604), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][17] ), .Z(
        n16122) );
  HS65_LH_NAND4ABX3 U17061 ( .A(n16125), .B(n16124), .C(n36266), .D(n16122), 
        .Z(n2285) );
  HS65_LH_AOI22X1 U17062 ( .A(n29606), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][17] ), .C(n29547), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[27][17] ), .Z(n16127)
         );
  HS65_LH_AOI22X1 U17063 ( .A(n29616), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][17] ), .C(n29618), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[16][17] ), .Z(n16126)
         );
  HS65_LH_NAND2X2 U17064 ( .A(n16127), .B(n16126), .Z(n16135) );
  HS65_LH_AO22X4 U17065 ( .A(n17412), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][17] ), .C(n16474), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][17] ), .Z(n16131)
         );
  HS65_LH_AO22X4 U17066 ( .A(n17407), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][17] ), .C(n40995), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][17] ), .Z(n16130)
         );
  HS65_LH_AOI22X1 U17067 ( .A(n16415), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][17] ), .C(n29560), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][17] ), .Z(n16129)
         );
  HS65_LH_AOI22X1 U17068 ( .A(n29553), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][17] ), .C(n40994), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][17] ), .Z(n16128)
         );
  HS65_LH_NAND4ABX3 U17069 ( .A(n16131), .B(n16130), .C(n16129), .D(n16128), 
        .Z(n16134) );
  HS65_LH_AOI22X1 U17070 ( .A(n29602), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][17] ), .C(n17410), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[31][17] ), .Z(n16133)
         );
  HS65_LH_AOI22X1 U17071 ( .A(n16379), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][17] ), .C(n29552), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][17] ), .Z(n16132)
         );
  HS65_LH_NAND4ABX3 U17072 ( .A(n16135), .B(n16134), .C(n16133), .D(n16132), 
        .Z(n2286) );
  HS65_LH_AOI22X1 U17073 ( .A(n36958), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][18] ), .C(n18125), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][18] ), .Z(
        n16137) );
  HS65_LH_AOI22X1 U17074 ( .A(n17426), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][18] ), .C(n16446), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][18] ), .Z(
        n16136) );
  HS65_LH_NAND2X2 U17075 ( .A(n16137), .B(n16136), .Z(n16145) );
  HS65_LH_AO22X4 U17076 ( .A(n17420), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][18] ), .C(n17432), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][18] ), .Z(
        n16141) );
  HS65_LH_AO22X4 U17077 ( .A(n18122), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][18] ), .C(n29604), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][18] ), .Z(
        n16140) );
  HS65_LH_AOI22X1 U17079 ( .A(n17430), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][18] ), .C(n17423), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][18] ), .Z(n16138)
         );
  HS65_LH_NAND4ABX3 U17080 ( .A(n16141), .B(n16140), .C(n16139), .D(n16138), 
        .Z(n16144) );
  HS65_LH_AOI22X1 U17081 ( .A(n17431), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][18] ), .C(n17427), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][18] ), .Z(n16143)
         );
  HS65_LH_AOI22X1 U17082 ( .A(n17421), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][18] ), .C(n17429), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[8][18] ), .Z(
        n16142) );
  HS65_LH_NAND4ABX3 U17083 ( .A(n16145), .B(n16144), .C(n16143), .D(n16142), 
        .Z(n2261) );
  HS65_LH_AOI22X1 U17084 ( .A(n17412), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][18] ), .C(n17408), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][18] ), .Z(n16147)
         );
  HS65_LH_AOI22X1 U17085 ( .A(n17409), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][18] ), .C(n18126), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][18] ), .Z(n16146)
         );
  HS65_LH_AO22X4 U17087 ( .A(n17411), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][18] ), .C(n16474), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][18] ), .Z(n16151)
         );
  HS65_LH_AO22X4 U17088 ( .A(n17418), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][18] ), .C(n17414), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[27][18] ), .Z(n16150)
         );
  HS65_LH_AOI22X1 U17089 ( .A(n17406), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][18] ), .C(n40993), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[31][18] ), .Z(n16149)
         );
  HS65_LH_AOI22X1 U17090 ( .A(n17415), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][18] ), .C(n17417), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][18] ), .Z(n16148)
         );
  HS65_LH_NAND4ABX3 U17091 ( .A(n16151), .B(n16150), .C(n16149), .D(n16148), 
        .Z(n16154) );
  HS65_LH_AOI22X1 U17092 ( .A(n18123), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][18] ), .C(n17416), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[17][18] ), .Z(n16153)
         );
  HS65_LH_AOI22X1 U17093 ( .A(n17405), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][18] ), .C(n29610), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][18] ), .Z(n16152)
         );
  HS65_LH_NAND4ABX3 U17094 ( .A(n16155), .B(n16154), .C(n16153), .D(n16152), 
        .Z(n2262) );
  HS65_LH_AOI22X1 U17095 ( .A(n17421), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][19] ), .C(n36385), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][19] ), .Z(
        n16157) );
  HS65_LH_AOI22X1 U17096 ( .A(n36958), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][19] ), .C(n29603), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][19] ), .Z(
        n16156) );
  HS65_LH_AO22X4 U17098 ( .A(n17426), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][19] ), .C(n20433), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][19] ), .Z(
        n16161) );
  HS65_LH_AO22X4 U17099 ( .A(n29620), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][19] ), .C(n17423), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][19] ), .Z(n16160)
         );
  HS65_LH_AOI22X1 U17100 ( .A(n17422), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][19] ), .C(n17424), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][19] ), .Z(
        n16159) );
  HS65_LH_AOI22X1 U17101 ( .A(n29549), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][19] ), .C(n29542), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][19] ), .Z(
        n16158) );
  HS65_LH_NAND4ABX3 U17102 ( .A(n16161), .B(n16160), .C(n16159), .D(n16158), 
        .Z(n16164) );
  HS65_LH_AOI22X1 U17103 ( .A(n18122), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][19] ), .C(n29543), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][19] ), .Z(
        n16163) );
  HS65_LH_AOI22X1 U17104 ( .A(n20916), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][19] ), .C(n36045), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[8][19] ), .Z(
        n16162) );
  HS65_LH_NAND4ABX3 U17105 ( .A(n16165), .B(n16164), .C(n16163), .D(n16162), 
        .Z(n2237) );
  HS65_LH_AOI22X1 U17106 ( .A(n29616), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][19] ), .C(n29606), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[17][19] ), .Z(n16167)
         );
  HS65_LH_AOI22X1 U17107 ( .A(n18123), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][19] ), .C(n36561), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][19] ), .Z(n16166)
         );
  HS65_LH_NAND2X2 U17108 ( .A(n16167), .B(n16166), .Z(n16175) );
  HS65_LH_AO22X4 U17109 ( .A(n17417), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][19] ), .C(n17412), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][19] ), .Z(n16171)
         );
  HS65_LH_AO22X4 U17110 ( .A(n16415), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][19] ), .C(n40994), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][19] ), .Z(n16170)
         );
  HS65_LH_AOI22X1 U17111 ( .A(n17407), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][19] ), .C(n17418), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][19] ), .Z(n16169)
         );
  HS65_LH_AOI22X1 U17112 ( .A(n17411), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][19] ), .C(n29560), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][19] ), .Z(n16168)
         );
  HS65_LH_NAND4ABX3 U17113 ( .A(n16171), .B(n16170), .C(n16169), .D(n16168), 
        .Z(n16174) );
  HS65_LH_AOI22X1 U17114 ( .A(n29618), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][19] ), .C(n16379), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][19] ), .Z(n16173)
         );
  HS65_LH_AOI22X1 U17115 ( .A(n29547), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][19] ), .C(n17410), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[31][19] ), .Z(n16172)
         );
  HS65_LH_NAND4ABX3 U17116 ( .A(n16175), .B(n16174), .C(n16173), .D(n16172), 
        .Z(n2238) );
  HS65_LH_AOI22X1 U17117 ( .A(n29620), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][20] ), .C(n17422), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][20] ), .Z(n16177) );
  HS65_LH_AOI22X1 U17118 ( .A(n29549), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][20] ), .C(n16446), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][20] ), .Z(
        n16176) );
  HS65_LH_NAND2X2 U17119 ( .A(n16177), .B(n16176), .Z(n16185) );
  HS65_LH_AO22X4 U17120 ( .A(n16342), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][20] ), .C(n17424), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][20] ), .Z(
        n16181) );
  HS65_LH_AO22X4 U17121 ( .A(n16406), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][20] ), .C(n17431), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][20] ), .Z(
        n16180) );
  HS65_LH_AOI22X1 U17122 ( .A(n18348), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][20] ), .C(n17430), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][20] ), .Z(
        n16179) );
  HS65_LH_AOI22X1 U17123 ( .A(n17420), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][20] ), .C(n29542), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][20] ), .Z(
        n16178) );
  HS65_LH_NAND4ABX3 U17124 ( .A(n16181), .B(n16180), .C(n16179), .D(n16178), 
        .Z(n16184) );
  HS65_LH_AOI22X1 U17125 ( .A(n29551), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][20] ), .C(n17425), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][20] ), .Z(
        n16183) );
  HS65_LH_AOI22X1 U17126 ( .A(n17429), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][20] ), .C(n20342), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][20] ), .Z(
        n16182) );
  HS65_LH_AOI22X1 U17128 ( .A(n29618), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][20] ), .C(n17415), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][20] ), .Z(n16187)
         );
  HS65_LH_AOI22X1 U17129 ( .A(n29602), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][20] ), .C(n36561), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][20] ), .Z(n16186)
         );
  HS65_LH_AO22X4 U17131 ( .A(n17412), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][20] ), .C(n17410), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[31][20] ), .Z(n16191)
         );
  HS65_LH_AO22X4 U17132 ( .A(n40995), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][20] ), .C(n29560), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][20] ), .Z(n16190)
         );
  HS65_LH_AOI22X1 U17133 ( .A(n29547), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][20] ), .C(n40994), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][20] ), .Z(n16189)
         );
  HS65_LH_AOI22X1 U17134 ( .A(n29616), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][20] ), .C(n29606), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[17][20] ), .Z(n16188)
         );
  HS65_LH_NAND4ABX3 U17135 ( .A(n16191), .B(n16190), .C(n16189), .D(n16188), 
        .Z(n16194) );
  HS65_LH_AOI22X1 U17136 ( .A(n29610), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][20] ), .C(n16415), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][20] ), .Z(n16193)
         );
  HS65_LH_AOI22X1 U17137 ( .A(n29552), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][20] ), .C(n29553), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][20] ), .Z(n16192)
         );
  HS65_LH_NAND4ABX3 U17138 ( .A(n36275), .B(n16194), .C(n16193), .D(n16192), 
        .Z(n2214) );
  HS65_LH_AOI22X1 U17139 ( .A(n17421), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][21] ), .C(n17423), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][21] ), .Z(
        n16197) );
  HS65_LH_AOI22X1 U17140 ( .A(n29554), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][21] ), .C(n16446), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][21] ), .Z(
        n16196) );
  HS65_LH_NAND2X2 U17141 ( .A(n16197), .B(n16196), .Z(n16205) );
  HS65_LH_AO22X4 U17142 ( .A(n17431), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][21] ), .C(n18125), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][21] ), .Z(n16201) );
  HS65_LH_AO22X4 U17143 ( .A(n18122), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][21] ), .C(n17422), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][21] ), .Z(
        n16200) );
  HS65_LH_AOI22X1 U17144 ( .A(n17427), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][21] ), .C(n17424), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][21] ), .Z(n16199) );
  HS65_LH_AOI22X1 U17145 ( .A(n36958), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][21] ), .C(n17426), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][21] ), .Z(
        n16198) );
  HS65_LH_NAND4ABX3 U17146 ( .A(n16201), .B(n16200), .C(n16199), .D(n16198), 
        .Z(n16204) );
  HS65_LH_AOI22X1 U17147 ( .A(n29543), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][21] ), .C(n29549), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][21] ), .Z(n16203) );
  HS65_LH_AOI22X1 U17148 ( .A(n17420), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][21] ), .C(n17425), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][21] ), .Z(
        n16202) );
  HS65_LH_NAND4ABX3 U17149 ( .A(n16205), .B(n16204), .C(n16203), .D(n16202), 
        .Z(n2189) );
  HS65_LH_AOI22X1 U17150 ( .A(n29606), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][21] ), .C(n29622), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][21] ), .Z(n16207)
         );
  HS65_LH_AOI22X1 U17151 ( .A(n17415), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][21] ), .C(n17408), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][21] ), .Z(n16206)
         );
  HS65_LH_NAND2X2 U17152 ( .A(n16207), .B(n16206), .Z(n16215) );
  HS65_LH_AO22X4 U17153 ( .A(n17407), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][21] ), .C(n18123), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][21] ), .Z(n16211)
         );
  HS65_LH_AO22X4 U17154 ( .A(n17405), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][21] ), .C(n17414), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[27][21] ), .Z(n16210)
         );
  HS65_LH_AOI22X1 U17155 ( .A(n17406), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][21] ), .C(n16474), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][21] ), .Z(n16209)
         );
  HS65_LH_AOI22X1 U17156 ( .A(n17409), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][21] ), .C(n17410), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[31][21] ), .Z(n16208)
         );
  HS65_LH_NAND4ABX3 U17157 ( .A(n16211), .B(n16210), .C(n16209), .D(n16208), 
        .Z(n16214) );
  HS65_LH_AOI22X1 U17158 ( .A(n40995), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][21] ), .C(n29553), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][21] ), .Z(n16213)
         );
  HS65_LH_AOI22X1 U17159 ( .A(n17418), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][21] ), .C(n36571), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][21] ), .Z(n16212)
         );
  HS65_LH_NAND4ABX3 U17160 ( .A(n16215), .B(n16214), .C(n16213), .D(n16212), 
        .Z(n2190) );
  HS65_LH_AOI22X1 U17161 ( .A(n17426), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][22] ), .C(n17423), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][22] ), .Z(
        n16217) );
  HS65_LH_AOI22X1 U17162 ( .A(n36958), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][22] ), .C(n29604), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][22] ), .Z(
        n16216) );
  HS65_LH_NAND2X2 U17163 ( .A(n16217), .B(n16216), .Z(n16225) );
  HS65_LH_AO22X4 U17164 ( .A(n17432), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][22] ), .C(n17431), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][22] ), .Z(
        n16221) );
  HS65_LH_AO22X4 U17165 ( .A(n20916), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][22] ), .C(n17429), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[8][22] ), .Z(
        n16220) );
  HS65_LH_AOI22X1 U17166 ( .A(n17421), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][22] ), .C(n18125), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][22] ), .Z(
        n16219) );
  HS65_LH_AOI22X1 U17167 ( .A(n18122), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][22] ), .C(n17425), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][22] ), .Z(
        n16218) );
  HS65_LH_NAND4ABX3 U17168 ( .A(n16221), .B(n16220), .C(n16219), .D(n16218), 
        .Z(n16224) );
  HS65_LH_AOI22X1 U17169 ( .A(n29543), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][22] ), .C(n17428), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][22] ), .Z(n16223)
         );
  HS65_LH_AOI22X1 U17170 ( .A(n29620), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][22] ), .C(n29561), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][22] ), .Z(n16222) );
  HS65_LH_AOI22X1 U17172 ( .A(n17407), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][22] ), .C(n17415), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][22] ), .Z(n16227)
         );
  HS65_LH_AOI22X1 U17173 ( .A(n40993), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][22] ), .C(n36571), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][22] ), .Z(n16226)
         );
  HS65_LH_NAND2X2 U17174 ( .A(n16227), .B(n16226), .Z(n16235) );
  HS65_LH_AO22X4 U17175 ( .A(n17414), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][22] ), .C(n16415), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][22] ), .Z(n16231)
         );
  HS65_LH_AO22X4 U17176 ( .A(n18123), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][22] ), .C(n17411), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][22] ), .Z(n16230)
         );
  HS65_LH_AOI22X1 U17177 ( .A(n17406), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][22] ), .C(n17408), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][22] ), .Z(n16229)
         );
  HS65_LH_AOI22X1 U17178 ( .A(n17418), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][22] ), .C(n29622), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][22] ), .Z(n16228)
         );
  HS65_LH_NAND4ABX3 U17179 ( .A(n16231), .B(n16230), .C(n16229), .D(n16228), 
        .Z(n16234) );
  HS65_LH_AOI22X1 U17180 ( .A(n29618), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][22] ), .C(n36759), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[17][22] ), .Z(n16233)
         );
  HS65_LH_NAND4ABX3 U17182 ( .A(n16235), .B(n16234), .C(n16233), .D(n16232), 
        .Z(n2166) );
  HS65_LH_AOI22X1 U17183 ( .A(n29543), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][23] ), .C(n29561), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][23] ), .Z(n16237) );
  HS65_LH_AOI22X1 U17184 ( .A(n36385), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][23] ), .C(n29620), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][23] ), .Z(n16236)
         );
  HS65_LH_NAND2X2 U17185 ( .A(n16237), .B(n16236), .Z(n16245) );
  HS65_LH_AO22X4 U17186 ( .A(n17421), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][23] ), .C(n29542), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][23] ), .Z(
        n16241) );
  HS65_LH_AO22X4 U17187 ( .A(n20916), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][23] ), .C(n20433), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][23] ), .Z(
        n16240) );
  HS65_LH_AOI22X1 U17188 ( .A(n36958), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][23] ), .C(n20342), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][23] ), .Z(
        n16239) );
  HS65_LH_AOI22X1 U17189 ( .A(n17431), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][23] ), .C(n17426), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][23] ), .Z(n16238) );
  HS65_LH_AOI22X1 U17191 ( .A(n36045), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][23] ), .C(n36264), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][23] ), .Z(
        n16243) );
  HS65_LH_AOI22X1 U17192 ( .A(n18348), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][23] ), .C(n29604), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][23] ), .Z(
        n16242) );
  HS65_LH_NAND4ABX3 U17193 ( .A(n16245), .B(n16244), .C(n16243), .D(n16242), 
        .Z(n2141) );
  HS65_LH_AOI22X1 U17194 ( .A(n29616), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][23] ), .C(n17405), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[16][23] ), .Z(n16247)
         );
  HS65_LH_AOI22X1 U17195 ( .A(n17418), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][23] ), .C(n36571), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][23] ), .Z(n16246)
         );
  HS65_LH_AO22X4 U17197 ( .A(n29606), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][23] ), .C(n17412), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][23] ), .Z(n16251)
         );
  HS65_LH_AO22X4 U17198 ( .A(n17411), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][23] ), .C(n17410), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[31][23] ), .Z(n16250)
         );
  HS65_LH_AOI22X1 U17199 ( .A(n17415), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][23] ), .C(n17408), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][23] ), .Z(n16249)
         );
  HS65_LH_AOI22X1 U17200 ( .A(n17407), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][23] ), .C(n36561), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][23] ), .Z(n16248)
         );
  HS65_LH_NAND4ABX3 U17201 ( .A(n16251), .B(n16250), .C(n16249), .D(n16248), 
        .Z(n16254) );
  HS65_LH_AOI22X1 U17202 ( .A(n40995), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][23] ), .C(n16415), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][23] ), .Z(n16253)
         );
  HS65_LH_AOI22X1 U17203 ( .A(n18123), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][23] ), .C(n29547), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[27][23] ), .Z(n16252)
         );
  HS65_LH_NAND4ABX3 U17204 ( .A(n16255), .B(n16254), .C(n16253), .D(n16252), 
        .Z(n2142) );
  HS65_LH_AOI22X1 U17205 ( .A(n36958), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][24] ), .C(n29603), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][24] ), .Z(
        n16257) );
  HS65_LH_AOI22X1 U17206 ( .A(n29554), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][24] ), .C(n29620), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][24] ), .Z(
        n16256) );
  HS65_LH_NAND2X2 U17207 ( .A(n16257), .B(n16256), .Z(n16265) );
  HS65_LH_AO22X4 U17208 ( .A(n17421), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][24] ), .C(n17423), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][24] ), .Z(
        n16261) );
  HS65_LH_AO22X4 U17209 ( .A(n17420), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][24] ), .C(n36264), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][24] ), .Z(
        n16260) );
  HS65_LH_AOI22X1 U17210 ( .A(n17426), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][24] ), .C(n36385), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][24] ), .Z(
        n16259) );
  HS65_LH_AOI22X1 U17211 ( .A(n18348), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][24] ), .C(n29543), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][24] ), .Z(
        n16258) );
  HS65_LH_NAND4ABX3 U17212 ( .A(n16261), .B(n16260), .C(n16259), .D(n16258), 
        .Z(n16264) );
  HS65_LH_AOI22X1 U17213 ( .A(n29542), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][24] ), .C(n29604), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][24] ), .Z(
        n16263) );
  HS65_LH_AOI22X1 U17214 ( .A(n17425), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][24] ), .C(n29561), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][24] ), .Z(n16262) );
  HS65_LH_NAND4ABX3 U17215 ( .A(n16265), .B(n16264), .C(n16263), .D(n35936), 
        .Z(n2117) );
  HS65_LH_AOI22X1 U17216 ( .A(n17412), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][24] ), .C(n17410), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[31][24] ), .Z(n16267)
         );
  HS65_LH_AOI22X1 U17217 ( .A(n17411), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][24] ), .C(n17414), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[27][24] ), .Z(n16266)
         );
  HS65_LH_NAND2X2 U17218 ( .A(n16267), .B(n16266), .Z(n16275) );
  HS65_LH_AO22X4 U17219 ( .A(n17407), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][24] ), .C(n16474), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][24] ), .Z(n16271)
         );
  HS65_LH_AO22X4 U17220 ( .A(n17417), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][24] ), .C(n17408), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][24] ), .Z(n16270)
         );
  HS65_LH_AOI22X1 U17221 ( .A(n17406), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][24] ), .C(n17409), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][24] ), .Z(n16269)
         );
  HS65_LH_AOI22X1 U17222 ( .A(n17418), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][24] ), .C(n29560), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][24] ), .Z(n16268)
         );
  HS65_LH_NAND4ABX3 U17223 ( .A(n16271), .B(n16270), .C(n16269), .D(n16268), 
        .Z(n16274) );
  HS65_LH_AOI22X1 U17224 ( .A(n36759), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][24] ), .C(n16379), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][24] ), .Z(n16273)
         );
  HS65_LH_AOI22X1 U17225 ( .A(n17405), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][24] ), .C(n29602), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][24] ), .Z(n16272)
         );
  HS65_LH_NAND4ABX3 U17226 ( .A(n16275), .B(n16274), .C(n16273), .D(n16272), 
        .Z(n2118) );
  HS65_LH_AOI22X1 U17227 ( .A(n17428), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][25] ), .C(n17427), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][25] ), .Z(n16277)
         );
  HS65_LH_AOI22X1 U17228 ( .A(n17421), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][25] ), .C(n17425), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][25] ), .Z(
        n16276) );
  HS65_LH_NAND2X2 U17229 ( .A(n16277), .B(n16276), .Z(n16285) );
  HS65_LH_AO22X4 U17230 ( .A(n17429), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][25] ), .C(n17423), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][25] ), .Z(
        n16281) );
  HS65_LH_AO22X4 U17231 ( .A(n16406), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][25] ), .C(n18348), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][25] ), .Z(
        n16280) );
  HS65_LH_AOI22X1 U17232 ( .A(n17420), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][25] ), .C(n29603), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][25] ), .Z(
        n16279) );
  HS65_LH_AOI22X1 U17233 ( .A(n17430), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][25] ), .C(n17424), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][25] ), .Z(n16278) );
  HS65_LH_AOI22X1 U17235 ( .A(n29549), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][25] ), .C(n29551), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][25] ), .Z(
        n16283) );
  HS65_LH_AOI22X1 U17236 ( .A(n29542), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][25] ), .C(n29604), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][25] ), .Z(
        n16282) );
  HS65_LH_NAND4ABX3 U17237 ( .A(n36857), .B(n16284), .C(n16283), .D(n16282), 
        .Z(n2093) );
  HS65_LH_AOI22X1 U17238 ( .A(n29552), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][25] ), .C(n16415), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][25] ), .Z(n16287)
         );
  HS65_LH_AOI22X1 U17239 ( .A(n29547), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][25] ), .C(n17410), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[31][25] ), .Z(n16286)
         );
  HS65_LH_NAND2X2 U17240 ( .A(n16287), .B(n16286), .Z(n16295) );
  HS65_LH_AO22X4 U17241 ( .A(n29602), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][25] ), .C(n17417), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][25] ), .Z(n16291)
         );
  HS65_LH_AO22X4 U17242 ( .A(n17416), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][25] ), .C(n17415), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][25] ), .Z(n16290)
         );
  HS65_LH_AOI22X1 U17243 ( .A(n29553), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][25] ), .C(n17408), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][25] ), .Z(n16289)
         );
  HS65_LH_AOI22X1 U17244 ( .A(n29616), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][25] ), .C(n16474), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][25] ), .Z(n16288)
         );
  HS65_LH_NAND4ABX3 U17245 ( .A(n16291), .B(n16290), .C(n16289), .D(n16288), 
        .Z(n16294) );
  HS65_LH_AOI22X1 U17246 ( .A(n17407), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][25] ), .C(n29560), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][25] ), .Z(n16293)
         );
  HS65_LH_AOI22X1 U17247 ( .A(n17405), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][25] ), .C(n29622), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][25] ), .Z(n16292)
         );
  HS65_LH_NAND4ABX3 U17248 ( .A(n16295), .B(n16294), .C(n16293), .D(n16292), 
        .Z(n2094) );
  HS65_LH_AOI22X1 U17249 ( .A(n29554), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][26] ), .C(n17424), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][26] ), .Z(
        n16297) );
  HS65_LH_AOI22X1 U17250 ( .A(n17423), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][26] ), .C(n20433), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][26] ), .Z(n16296)
         );
  HS65_LH_NAND2X2 U17251 ( .A(n16297), .B(n16296), .Z(n16305) );
  HS65_LH_AO22X4 U17252 ( .A(n16406), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][26] ), .C(n18125), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][26] ), .Z(
        n16301) );
  HS65_LH_AO22X4 U17253 ( .A(n17420), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][26] ), .C(n17422), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][26] ), .Z(
        n16300) );
  HS65_LH_AOI22X1 U17254 ( .A(n16446), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][26] ), .C(n17427), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][26] ), .Z(n16299)
         );
  HS65_LH_AOI22X1 U17255 ( .A(n18348), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][26] ), .C(n29543), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][26] ), .Z(
        n16298) );
  HS65_LH_AOI22X1 U17258 ( .A(n16342), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][26] ), .C(n29551), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][26] ), .Z(
        n16302) );
  HS65_LH_NAND4ABX3 U17259 ( .A(n16305), .B(n16304), .C(n29535), .D(n16302), 
        .Z(n2069) );
  HS65_LH_AOI22X1 U17260 ( .A(n29606), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][26] ), .C(n40995), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][26] ), .Z(n16307)
         );
  HS65_LH_AOI22X1 U17261 ( .A(n29618), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][26] ), .C(n29547), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[27][26] ), .Z(n16306)
         );
  HS65_LH_NAND2X2 U17262 ( .A(n16307), .B(n16306), .Z(n16316) );
  HS65_LH_AO22X4 U17263 ( .A(n17406), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][26] ), .C(n17407), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][26] ), .Z(n16312)
         );
  HS65_LH_AO22X4 U17264 ( .A(n17411), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][26] ), .C(n17408), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][26] ), .Z(n16311)
         );
  HS65_LH_AOI22X1 U17265 ( .A(n16415), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][26] ), .C(n40993), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[31][26] ), .Z(n16310)
         );
  HS65_LH_AOI22X1 U17266 ( .A(n29622), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][26] ), .C(n36571), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][26] ), .Z(n16309)
         );
  HS65_LH_AOI22X1 U17268 ( .A(n29602), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][26] ), .C(n16379), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][26] ), .Z(n16314)
         );
  HS65_LH_AOI22X1 U17269 ( .A(n17418), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][26] ), .C(n36561), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][26] ), .Z(n16313)
         );
  HS65_LH_NAND4ABX3 U17270 ( .A(n16316), .B(n16315), .C(n16314), .D(n16313), 
        .Z(n2070) );
  HS65_LH_AOI22X1 U17271 ( .A(n29542), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][27] ), .C(n36385), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][27] ), .Z(
        n16319) );
  HS65_LH_AOI22X1 U17272 ( .A(n16342), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][27] ), .C(n29561), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][27] ), .Z(
        n16318) );
  HS65_LH_NAND2X2 U17273 ( .A(n16319), .B(n16318), .Z(n16328) );
  HS65_LH_AO22X4 U17274 ( .A(n36045), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][27] ), .C(n17422), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][27] ), .Z(
        n16323) );
  HS65_LH_AO22X4 U17275 ( .A(n17426), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][27] ), .C(n29620), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][27] ), .Z(
        n16322) );
  HS65_LH_AOI22X1 U17276 ( .A(n18122), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][27] ), .C(n17423), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][27] ), .Z(
        n16321) );
  HS65_LH_AOI22X1 U17277 ( .A(n17430), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][27] ), .C(n35786), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][27] ), .Z(n16320)
         );
  HS65_LH_AOI22X1 U17279 ( .A(n20916), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][27] ), .C(n17431), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][27] ), .Z(
        n16326) );
  HS65_LH_AOI22X1 U17280 ( .A(n16406), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][27] ), .C(n29549), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][27] ), .Z(
        n16325) );
  HS65_LH_NAND4ABX3 U17281 ( .A(n16328), .B(n16327), .C(n35732), .D(n16325), 
        .Z(n2045) );
  HS65_LH_AOI22X1 U17282 ( .A(n17411), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][27] ), .C(n17414), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[27][27] ), .Z(n16330)
         );
  HS65_LH_AOI22X1 U17283 ( .A(n17407), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][27] ), .C(n29552), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][27] ), .Z(n16329)
         );
  HS65_LH_NAND2X2 U17284 ( .A(n16330), .B(n16329), .Z(n16338) );
  HS65_LH_AO22X4 U17285 ( .A(n17406), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][27] ), .C(n17405), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[16][27] ), .Z(n16334)
         );
  HS65_LH_AO22X4 U17286 ( .A(n17412), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][27] ), .C(n17410), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[31][27] ), .Z(n16333)
         );
  HS65_LH_AOI22X1 U17287 ( .A(n17417), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][27] ), .C(n17409), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][27] ), .Z(n16332)
         );
  HS65_LH_AOI22X1 U17288 ( .A(n16474), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][27] ), .C(n40994), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][27] ), .Z(n16331)
         );
  HS65_LH_NAND4ABX3 U17289 ( .A(n16334), .B(n16333), .C(n16332), .D(n16331), 
        .Z(n16337) );
  HS65_LH_AOI22X1 U17290 ( .A(n18123), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][27] ), .C(n16379), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][27] ), .Z(n16336)
         );
  HS65_LH_AOI22X1 U17291 ( .A(n36759), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][27] ), .C(n36571), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][27] ), .Z(n16335)
         );
  HS65_LH_NAND4ABX3 U17292 ( .A(n16338), .B(n16337), .C(n16336), .D(n16335), 
        .Z(n2046) );
  HS65_LH_AOI22X1 U17293 ( .A(n29554), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][28] ), .C(n17425), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][28] ), .Z(
        n16340) );
  HS65_LH_AOI22X1 U17294 ( .A(n29551), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][28] ), .C(n29620), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][28] ), .Z(
        n16339) );
  HS65_LH_NAND2X2 U17295 ( .A(n16340), .B(n16339), .Z(n16350) );
  HS65_LH_AO22X4 U17296 ( .A(n29603), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][28] ), .C(n17424), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][28] ), .Z(n16346) );
  HS65_LH_AO22X4 U17297 ( .A(n29549), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][28] ), .C(n29542), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][28] ), .Z(
        n16345) );
  HS65_LH_AOI22X1 U17298 ( .A(n36958), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][28] ), .C(n20342), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][28] ), .Z(
        n16344) );
  HS65_LH_AOI22X1 U17299 ( .A(n17420), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][28] ), .C(n16342), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][28] ), .Z(
        n16343) );
  HS65_LH_NAND4ABX3 U17300 ( .A(n16346), .B(n16345), .C(n16344), .D(n16343), 
        .Z(n16349) );
  HS65_LH_AOI22X1 U17301 ( .A(n29543), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][28] ), .C(n16446), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][28] ), .Z(n16348)
         );
  HS65_LH_AOI22X1 U17302 ( .A(n18122), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][28] ), .C(n29604), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][28] ), .Z(
        n16347) );
  HS65_LH_NAND4ABX3 U17303 ( .A(n16350), .B(n16349), .C(n16348), .D(n16347), 
        .Z(n2021) );
  HS65_LH_AOI22X1 U17304 ( .A(n29610), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][28] ), .C(n17409), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][28] ), .Z(n16354)
         );
  HS65_LH_AOI22X1 U17305 ( .A(n17411), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][28] ), .C(n36561), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][28] ), .Z(n16353)
         );
  HS65_LH_NAND2X2 U17306 ( .A(n16354), .B(n16353), .Z(n16363) );
  HS65_LH_AO22X4 U17307 ( .A(n16379), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][28] ), .C(n17418), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][28] ), .Z(n16358)
         );
  HS65_LH_AO22X4 U17308 ( .A(n17412), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][28] ), .C(n17410), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[31][28] ), .Z(n16357)
         );
  HS65_LH_AOI22X1 U17309 ( .A(n17406), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][28] ), .C(n29547), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[27][28] ), .Z(n16356)
         );
  HS65_LH_AOI22X1 U17310 ( .A(n29618), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][28] ), .C(n40994), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][28] ), .Z(n16355)
         );
  HS65_LH_NAND4ABX3 U17311 ( .A(n16358), .B(n16357), .C(n16356), .D(n16355), 
        .Z(n16362) );
  HS65_LH_AOI22X1 U17312 ( .A(n36759), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][28] ), .C(n29560), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][28] ), .Z(n16361)
         );
  HS65_LH_AOI22X1 U17313 ( .A(n18123), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][28] ), .C(n40995), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][28] ), .Z(n16360)
         );
  HS65_LH_NAND4ABX3 U17314 ( .A(n16363), .B(n16362), .C(n16361), .D(n16360), 
        .Z(n2022) );
  HS65_LH_AOI22X1 U17315 ( .A(n18348), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][29] ), .C(n17424), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][29] ), .Z(
        n16365) );
  HS65_LH_AOI22X1 U17316 ( .A(n17426), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][29] ), .C(n17425), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][29] ), .Z(
        n16364) );
  HS65_LH_NAND2X2 U17317 ( .A(n16365), .B(n16364), .Z(n16376) );
  HS65_LH_AO22X4 U17318 ( .A(n17420), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][29] ), .C(n17427), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][29] ), .Z(
        n16372) );
  HS65_LH_AO22X4 U17319 ( .A(n17431), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][29] ), .C(n16446), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][29] ), .Z(n16371)
         );
  HS65_LH_AOI22X1 U17320 ( .A(n17421), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][29] ), .C(n18125), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][29] ), .Z(
        n16370) );
  HS65_LH_AOI22X1 U17321 ( .A(n17430), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][29] ), .C(n36045), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[8][29] ), .Z(n16369) );
  HS65_LH_NAND4ABX3 U17322 ( .A(n16372), .B(n16371), .C(n16370), .D(n16369), 
        .Z(n16375) );
  HS65_LH_AOI22X1 U17323 ( .A(n20342), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][29] ), .C(n29604), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][29] ), .Z(n16374) );
  HS65_LH_AOI22X1 U17324 ( .A(n16406), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][29] ), .C(n29549), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][29] ), .Z(
        n16373) );
  HS65_LH_NAND4ABX3 U17325 ( .A(n16376), .B(n16375), .C(n16374), .D(n16373), 
        .Z(n1997) );
  HS65_LH_AOI22X1 U17326 ( .A(n40995), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][29] ), .C(n17409), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][29] ), .Z(n16381)
         );
  HS65_LH_AOI22X1 U17327 ( .A(n16379), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][29] ), .C(n36571), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][29] ), .Z(n16380)
         );
  HS65_LH_AO22X4 U17329 ( .A(n29547), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][29] ), .C(n16474), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][29] ), .Z(n16386)
         );
  HS65_LH_AO22X4 U17330 ( .A(n29606), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][29] ), .C(n29553), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][29] ), .Z(n16385)
         );
  HS65_LH_AOI22X1 U17331 ( .A(n29602), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][29] ), .C(n17410), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[31][29] ), .Z(n16384)
         );
  HS65_LH_AOI22X1 U17332 ( .A(n29616), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][29] ), .C(n40994), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][29] ), .Z(n16383)
         );
  HS65_LH_NAND4ABX3 U17333 ( .A(n16386), .B(n16385), .C(n16384), .D(n16383), 
        .Z(n16390) );
  HS65_LH_AOI22X1 U17334 ( .A(n17405), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][29] ), .C(n29622), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][29] ), .Z(n16389)
         );
  HS65_LH_AOI22X1 U17335 ( .A(n29610), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][29] ), .C(n29552), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][29] ), .Z(n16388)
         );
  HS65_LH_NAND4ABX3 U17336 ( .A(n16391), .B(n16390), .C(n16389), .D(n16388), 
        .Z(n1998) );
  HS65_LH_AOI22X1 U17337 ( .A(n29554), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][30] ), .C(n29604), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][30] ), .Z(
        n16397) );
  HS65_LH_AOI22X1 U17338 ( .A(n36264), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][30] ), .C(n17426), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][30] ), .Z(
        n16396) );
  HS65_LH_NAND2X2 U17339 ( .A(n16397), .B(n16396), .Z(n16410) );
  HS65_LH_AO22X4 U17340 ( .A(n17430), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][30] ), .C(n17431), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][30] ), .Z(n16404)
         );
  HS65_LH_AO22X4 U17341 ( .A(n18122), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][30] ), .C(n20433), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][30] ), .Z(
        n16403) );
  HS65_LH_AOI22X1 U17342 ( .A(n29620), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][30] ), .C(n17424), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][30] ), .Z(n16402) );
  HS65_LH_AOI22X1 U17343 ( .A(n17421), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][30] ), .C(n18125), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][30] ), .Z(
        n16401) );
  HS65_LH_NAND4ABX3 U17344 ( .A(n16404), .B(n16403), .C(n16402), .D(n16401), 
        .Z(n16409) );
  HS65_LH_AOI22X1 U17345 ( .A(n17420), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][30] ), .C(n16446), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][30] ), .Z(
        n16408) );
  HS65_LH_NAND4ABX3 U17347 ( .A(n16410), .B(n16409), .C(n16408), .D(n29536), 
        .Z(n1973) );
  HS65_LH_AOI22X1 U17348 ( .A(n17414), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][30] ), .C(n29560), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][30] ), .Z(n16414)
         );
  HS65_LH_AOI22X1 U17349 ( .A(n29610), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][30] ), .C(n17418), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][30] ), .Z(n16413)
         );
  HS65_LH_NAND2X2 U17350 ( .A(n16414), .B(n16413), .Z(n16427) );
  HS65_LH_AO22X4 U17351 ( .A(n18123), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][30] ), .C(n16415), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][30] ), .Z(n16421)
         );
  HS65_LH_AO22X4 U17352 ( .A(n17406), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][30] ), .C(n17412), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][30] ), .Z(n16420)
         );
  HS65_LH_AOI22X1 U17353 ( .A(n17415), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][30] ), .C(n16474), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][30] ), .Z(n16419)
         );
  HS65_LH_AOI22X1 U17354 ( .A(n17417), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][30] ), .C(n17410), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[31][30] ), .Z(n16418)
         );
  HS65_LH_NAND4ABX3 U17355 ( .A(n16421), .B(n16420), .C(n16419), .D(n16418), 
        .Z(n16426) );
  HS65_LH_AOI22X1 U17356 ( .A(n17405), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][30] ), .C(n40994), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][30] ), .Z(n16425)
         );
  HS65_LH_AOI22X1 U17357 ( .A(n36759), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][30] ), .C(n29553), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][30] ), .Z(n16424)
         );
  HS65_LH_AOI22X1 U17359 ( .A(n17421), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][31] ), .C(n17422), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][31] ), .Z(
        n16433) );
  HS65_LH_AOI22X1 U17360 ( .A(n17430), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][31] ), .C(n17431), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][31] ), .Z(n16432)
         );
  HS65_LH_NAND2X2 U17361 ( .A(n16433), .B(n16432), .Z(n16453) );
  HS65_LH_AO22X4 U17362 ( .A(n17429), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][31] ), .C(n18125), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][31] ), .Z(
        n16445) );
  HS65_LH_AO22X4 U17363 ( .A(n17427), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][31] ), .C(n17425), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][31] ), .Z(n16444)
         );
  HS65_LH_AOI22X1 U17364 ( .A(n36958), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][31] ), .C(n17424), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][31] ), .Z(
        n16443) );
  HS65_LH_AOI22X1 U17365 ( .A(n18122), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][31] ), .C(n29549), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][31] ), .Z(
        n16442) );
  HS65_LH_NAND4ABX3 U17366 ( .A(n16445), .B(n16444), .C(n16443), .D(n16442), 
        .Z(n16452) );
  HS65_LH_AOI22X1 U17368 ( .A(n17426), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][31] ), .C(n20342), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][31] ), .Z(
        n16450) );
  HS65_LH_NAND4ABX3 U17369 ( .A(n16453), .B(n16452), .C(n40988), .D(n16450), 
        .Z(n1949) );
  HS65_LH_AOI22X1 U17370 ( .A(n17416), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][31] ), .C(n17417), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][31] ), .Z(n16459)
         );
  HS65_LH_AOI22X1 U17371 ( .A(n17406), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][31] ), .C(n17415), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][31] ), .Z(n16458)
         );
  HS65_LH_NAND2X2 U17372 ( .A(n16459), .B(n16458), .Z(n16479) );
  HS65_LH_AO22X4 U17373 ( .A(n17414), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][31] ), .C(n18126), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][31] ), .Z(n16471)
         );
  HS65_LH_AO22X4 U17374 ( .A(n17418), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][31] ), .C(n40993), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[31][31] ), .Z(n16470)
         );
  HS65_LH_AOI22X1 U17375 ( .A(n17411), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][31] ), .C(n17409), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][31] ), .Z(n16469)
         );
  HS65_LH_AOI22X1 U17376 ( .A(n18123), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][31] ), .C(n40994), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][31] ), .Z(n16468)
         );
  HS65_LH_NAND4ABX3 U17377 ( .A(n16471), .B(n16470), .C(n16469), .D(n16468), 
        .Z(n16478) );
  HS65_LH_AOI22X1 U17378 ( .A(n17405), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][31] ), .C(n17407), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][31] ), .Z(n16477)
         );
  HS65_LH_AOI22X1 U17379 ( .A(n17412), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][31] ), .C(n16474), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][31] ), .Z(n16476)
         );
  HS65_LH_NAND4ABX3 U17380 ( .A(n16479), .B(n16478), .C(n16477), .D(n16476), 
        .Z(n1950) );
  HS65_LH_NAND3X2 U17381 ( .A(n15169), .B(n15167), .C(n15170), .Z(n16482) );
  HS65_LH_NOR2X5 U17382 ( .A(n16503), .B(n16482), .Z(n17153) );
  HS65_LH_NAND3X2 U17383 ( .A(n12426), .B(n12446), .C(n15170), .Z(n16489) );
  HS65_LH_NOR2X5 U17384 ( .A(n16489), .B(n16503), .Z(n17066) );
  HS65_LH_AOI22X1 U17385 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][0] ), .B(n29623), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][0] ), .D(
        n17403), .Z(n16481) );
  HS65_LH_NOR2X5 U17386 ( .A(n16507), .B(n16482), .Z(n17090) );
  HS65_LH_NAND3X2 U17387 ( .A(n12446), .B(n15167), .C(n15170), .Z(n16488) );
  HS65_LH_AOI22X1 U17388 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][0] ), .B(n17402), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][0] ), .D(
        n18124), .Z(n16480) );
  HS65_LH_NAND2X2 U17389 ( .A(n16481), .B(n16480), .Z(n16494) );
  HS65_LH_NOR2X5 U17390 ( .A(n16505), .B(n16482), .Z(n17114) );
  HS65_LH_NOR2X5 U17391 ( .A(n16489), .B(n16507), .Z(n17147) );
  HS65_LH_AO22X4 U17392 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][0] ), .B(n17401), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][0] ), .D(
        n17400), .Z(n16487) );
  HS65_LH_NOR2X5 U17393 ( .A(n16505), .B(n16488), .Z(n17158) );
  HS65_LH_BFX4 U17394 ( .A(n17399), .Z(n17121) );
  HS65_LH_NOR2X5 U17395 ( .A(n16489), .B(n16497), .Z(n17156) );
  HS65_LH_BFX4 U17396 ( .A(n17398), .Z(n17065) );
  HS65_LH_AO22X4 U17397 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][0] ), .B(n17121), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][0] ), .D(
        n17065), .Z(n16486) );
  HS65_LH_NOR2X5 U17398 ( .A(n16482), .B(n16497), .Z(n17060) );
  HS65_LH_NAND3X2 U17399 ( .A(n12426), .B(n15169), .C(n15170), .Z(n16490) );
  HS65_LH_BFX4 U17400 ( .A(n18121), .Z(n17120) );
  HS65_LH_AOI22X1 U17401 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][0] ), .B(n17397), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][0] ), .D(
        n17120), .Z(n16485) );
  HS65_LH_NOR2X5 U17402 ( .A(n16488), .B(n16507), .Z(n17110) );
  HS65_LH_NOR2X2 U17403 ( .A(n16490), .B(n16507), .Z(n16483) );
  HS65_LH_BFX4 U17404 ( .A(n16483), .Z(n17035) );
  HS65_LH_AOI22X1 U17405 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][0] ), .B(n21638), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][0] ), .D(
        n17565), .Z(n16484) );
  HS65_LH_NAND4ABX3 U17406 ( .A(n16487), .B(n16486), .C(n16485), .D(n16484), 
        .Z(n16493) );
  HS65_LH_NOR2X5 U17407 ( .A(n16503), .B(n16488), .Z(n17146) );
  HS65_LH_BFX4 U17408 ( .A(n17394), .Z(n17057) );
  HS65_LH_NOR2X5 U17409 ( .A(n16490), .B(n16503), .Z(n17083) );
  HS65_LH_BFX4 U17410 ( .A(n17393), .Z(n17166) );
  HS65_LH_AOI22X1 U17411 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][0] ), .B(n17057), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][0] ), .D(
        n17166), .Z(n16492) );
  HS65_LH_NOR2X5 U17412 ( .A(n16505), .B(n16489), .Z(n17111) );
  HS65_LH_NOR2X5 U17413 ( .A(n16505), .B(n16490), .Z(n17092) );
  HS65_LH_BFX4 U17414 ( .A(n17391), .Z(n17148) );
  HS65_LH_AOI22X1 U17415 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][0] ), .B(n17392), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][0] ), .D(
        n17148), .Z(n16491) );
  HS65_LH_NAND4ABX3 U17416 ( .A(n16494), .B(n16493), .C(n16492), .D(n16491), 
        .Z(n1896) );
  HS65_LH_NAND3X2 U17417 ( .A(n12446), .B(n12471), .C(n15167), .Z(n16506) );
  HS65_LH_NOR2X5 U17418 ( .A(n16497), .B(n16506), .Z(n17045) );
  HS65_LH_NAND3X2 U17419 ( .A(n12426), .B(n12471), .C(n15169), .Z(n16504) );
  HS65_LH_NOR2X5 U17420 ( .A(n16497), .B(n16504), .Z(n17178) );
  HS65_LH_BFX4 U17421 ( .A(n17389), .Z(n17073) );
  HS65_LH_AOI22X1 U17422 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][0] ), .B(n17390), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][0] ), .D(
        n17073), .Z(n16496) );
  HS65_LH_NOR2X5 U17423 ( .A(n16503), .B(n16504), .Z(n17048) );
  HS65_LH_NOR2X5 U17424 ( .A(n16503), .B(n16506), .Z(n17174) );
  HS65_LH_AOI22X1 U17425 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][0] ), .B(n17388), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][0] ), .D(
        n17387), .Z(n16495) );
  HS65_LH_NAND2X2 U17426 ( .A(n16496), .B(n16495), .Z(n16512) );
  HS65_LH_NAND3X2 U17427 ( .A(n12471), .B(n15169), .C(n15167), .Z(n16508) );
  HS65_LH_NOR2X5 U17428 ( .A(n16505), .B(n16508), .Z(n17132) );
  HS65_LH_NAND3X2 U17429 ( .A(n12446), .B(n12426), .C(n12471), .Z(n16498) );
  HS65_LH_NOR2X5 U17430 ( .A(n16497), .B(n16498), .Z(n17171) );
  HS65_LH_BFX4 U17431 ( .A(n17385), .Z(n17140) );
  HS65_LH_AO22X4 U17432 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][0] ), .B(n17386), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[31][0] ), .D(
        n17140), .Z(n16502) );
  HS65_LH_NOR2X5 U17433 ( .A(n16507), .B(n16504), .Z(n17173) );
  HS65_LH_BFX4 U17434 ( .A(n17384), .Z(n17141) );
  HS65_LH_NOR2X5 U17435 ( .A(n16503), .B(n16498), .Z(n17184) );
  HS65_LH_BFX4 U17436 ( .A(n17383), .Z(n17074) );
  HS65_LH_AO22X4 U17437 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][0] ), .B(n17141), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][0] ), .D(
        n17074), .Z(n16501) );
  HS65_LH_NOR2X5 U17438 ( .A(n16505), .B(n16498), .Z(n17101) );
  HS65_LH_AOI22X1 U17439 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][0] ), .B(n17517), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][0] ), .D(
        n17382), .Z(n16500) );
  HS65_LH_NOR2X5 U17440 ( .A(n16505), .B(n16506), .Z(n17134) );
  HS65_LH_NOR2X5 U17441 ( .A(n16507), .B(n16498), .Z(n17133) );
  HS65_LH_AOI22X1 U17442 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][0] ), .B(n17381), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][0] ), .D(
        n17380), .Z(n16499) );
  HS65_LH_NAND4ABX3 U17443 ( .A(n16502), .B(n16501), .C(n16500), .D(n16499), 
        .Z(n16511) );
  HS65_LH_BFX4 U17444 ( .A(n17182), .Z(n17097) );
  HS65_LH_NOR2X5 U17445 ( .A(n16505), .B(n16504), .Z(n17172) );
  HS65_LH_AOI22X1 U17446 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][0] ), .B(n17564), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][0] ), .D(
        n17379), .Z(n16510) );
  HS65_LH_NOR2X5 U17447 ( .A(n16507), .B(n16506), .Z(n17139) );
  HS65_LH_NOR2X5 U17448 ( .A(n16497), .B(n16508), .Z(n17127) );
  HS65_LH_AOI22X1 U17449 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][0] ), .B(n17378), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][0] ), .D(
        n17377), .Z(n16509) );
  HS65_LH_NAND4ABX3 U17450 ( .A(n16512), .B(n16511), .C(n16510), .D(n16509), 
        .Z(n1897) );
  HS65_LH_BFX4 U17451 ( .A(n17397), .Z(n17149) );
  HS65_LH_AOI22X1 U17452 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][1] ), .B(n17392), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][1] ), .D(
        n17149), .Z(n16514) );
  HS65_LH_BFX4 U17453 ( .A(n17400), .Z(n17040) );
  HS65_LH_AOI22X1 U17454 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][1] ), .B(n17391), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][1] ), .D(
        n17040), .Z(n16513) );
  HS65_LH_AO22X4 U17456 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][1] ), .B(n18124), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][1] ), .D(
        n18121), .Z(n16518) );
  HS65_LH_BFX4 U17457 ( .A(n17403), .Z(n17152) );
  HS65_LH_BFX4 U17458 ( .A(n17401), .Z(n17165) );
  HS65_LH_AO22X4 U17459 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][1] ), .B(n17152), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][1] ), .D(
        n17165), .Z(n16517) );
  HS65_LH_BFX4 U17460 ( .A(n17402), .Z(n17154) );
  HS65_LH_AOI22X1 U17461 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][1] ), .B(n17121), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][1] ), .D(
        n17154), .Z(n16516) );
  HS65_LH_BFX4 U17462 ( .A(n16483), .Z(n17122) );
  HS65_LH_AOI22X1 U17463 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][1] ), .B(n17563), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][1] ), .D(
        n17393), .Z(n16515) );
  HS65_LH_AOI22X1 U17466 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][1] ), .B(n17057), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][1] ), .D(
        n29623), .Z(n16520) );
  HS65_LH_AOI22X1 U17468 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][1] ), .B(n21638), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][1] ), .D(
        n17065), .Z(n16519) );
  HS65_LH_NAND4ABX3 U17469 ( .A(n37931), .B(n37930), .C(n16520), .D(n16519), 
        .Z(n1840) );
  HS65_LH_BFX4 U17470 ( .A(n17387), .Z(n17130) );
  HS65_LH_AOI22X1 U17471 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][1] ), .B(n17516), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][1] ), .D(
        n17130), .Z(n16524) );
  HS65_LH_BFX4 U17472 ( .A(n17379), .Z(n17100) );
  HS65_LH_AOI22X1 U17473 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][1] ), .B(n17380), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][1] ), .D(
        n17100), .Z(n16523) );
  HS65_LH_NAND2X2 U17474 ( .A(n16524), .B(n16523), .Z(n16532) );
  HS65_LH_BFX4 U17475 ( .A(n17382), .Z(n17179) );
  HS65_LH_AO22X4 U17476 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][1] ), .B(n17179), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][1] ), .D(
        n17383), .Z(n16528) );
  HS65_LH_BFX4 U17477 ( .A(n17390), .Z(n17177) );
  HS65_LH_AO22X4 U17478 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][1] ), .B(n17177), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][1] ), .D(
        n17388), .Z(n16527) );
  HS65_LH_AOI22X1 U17479 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][1] ), .B(n17389), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][1] ), .D(
        n17384), .Z(n16526) );
  HS65_LH_BFX4 U17480 ( .A(n17381), .Z(n17180) );
  HS65_LH_AOI22X1 U17481 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][1] ), .B(n17385), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][1] ), .D(
        n17180), .Z(n16525) );
  HS65_LH_NAND4ABX3 U17482 ( .A(n16528), .B(n16527), .C(n16526), .D(n16525), 
        .Z(n16531) );
  HS65_LH_BFX4 U17483 ( .A(n17386), .Z(n17190) );
  HS65_LH_BFX4 U17484 ( .A(n17131), .Z(n17183) );
  HS65_LH_AOI22X1 U17485 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][1] ), .B(n17190), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[17][1] ), .D(
        n17562), .Z(n16530) );
  HS65_LH_BFX4 U17486 ( .A(n17378), .Z(n17192) );
  HS65_LH_AOI22X1 U17487 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][1] ), .B(n17377), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][1] ), .D(
        n17192), .Z(n16529) );
  HS65_LH_NAND4ABX3 U17488 ( .A(n16532), .B(n16531), .C(n16530), .D(n16529), 
        .Z(n1841) );
  HS65_LH_AOI22X1 U17489 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][2] ), .B(n17152), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][2] ), .D(
        n17165), .Z(n16534) );
  HS65_LH_AOI22X1 U17490 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][2] ), .B(n17399), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][2] ), .D(
        n17120), .Z(n16533) );
  HS65_LH_NAND2X2 U17491 ( .A(n16534), .B(n16533), .Z(n16542) );
  HS65_LH_AO22X4 U17492 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][2] ), .B(n17392), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][2] ), .D(
        n17404), .Z(n16538) );
  HS65_LH_AO22X4 U17493 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][2] ), .B(n17057), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][2] ), .D(
        n17393), .Z(n16537) );
  HS65_LH_BFX4 U17494 ( .A(n18124), .Z(n17155) );
  HS65_LH_AOI22X1 U17495 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][2] ), .B(n17397), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][2] ), .D(
        n17155), .Z(n16536) );
  HS65_LH_AOI22X1 U17496 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][2] ), .B(n21638), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][2] ), .D(
        n17148), .Z(n16535) );
  HS65_LH_NAND4ABX3 U17497 ( .A(n16538), .B(n16537), .C(n16536), .D(n16535), 
        .Z(n16541) );
  HS65_LH_AOI22X1 U17498 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][2] ), .B(n17040), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][2] ), .D(
        n17065), .Z(n16540) );
  HS65_LH_AOI22X1 U17499 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][2] ), .B(n17402), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][2] ), .D(
        n17565), .Z(n16539) );
  HS65_LH_NAND4ABX3 U17500 ( .A(n16542), .B(n16541), .C(n16540), .D(n38428), 
        .Z(n1817) );
  HS65_LH_AOI22X1 U17501 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][2] ), .B(n17517), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][2] ), .D(
        n17180), .Z(n16544) );
  HS65_LH_BFX4 U17502 ( .A(n17388), .Z(n17181) );
  HS65_LH_BFX4 U17503 ( .A(n17377), .Z(n17189) );
  HS65_LH_AOI22X1 U17504 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][2] ), .B(n17181), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][2] ), .D(
        n17189), .Z(n16543) );
  HS65_LH_NAND2X2 U17505 ( .A(n16544), .B(n16543), .Z(n16552) );
  HS65_LH_BFX4 U17506 ( .A(n17380), .Z(n17191) );
  HS65_LH_AO22X4 U17507 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][2] ), .B(n17191), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][2] ), .D(
        n17179), .Z(n16548) );
  HS65_LH_AO22X4 U17508 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][2] ), .B(n17074), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][2] ), .D(
        n17100), .Z(n16547) );
  HS65_LH_AOI22X1 U17509 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][2] ), .B(n17141), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[31][2] ), .D(
        n17140), .Z(n16546) );
  HS65_LH_AOI22X1 U17510 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][2] ), .B(n17389), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[27][2] ), .D(
        n17390), .Z(n16545) );
  HS65_LH_NAND4ABX3 U17511 ( .A(n16548), .B(n16547), .C(n16546), .D(n16545), 
        .Z(n16551) );
  HS65_LH_AOI22X1 U17512 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][2] ), .B(n17564), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][2] ), .D(
        n17190), .Z(n16550) );
  HS65_LH_AOI22X1 U17513 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][2] ), .B(n17387), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][2] ), .D(
        n17192), .Z(n16549) );
  HS65_LH_NAND4ABX3 U17514 ( .A(n16552), .B(n16551), .C(n16550), .D(n16549), 
        .Z(n1818) );
  HS65_LH_AOI22X1 U17515 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][3] ), .B(n29623), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][3] ), .D(
        n17395), .Z(n16554) );
  HS65_LH_AOI22X1 U17516 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][3] ), .B(n17152), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][3] ), .D(
        n17149), .Z(n16553) );
  HS65_LH_AO22X4 U17518 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][3] ), .B(n17121), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[9][3] ), .D(
        n17396), .Z(n16558) );
  HS65_LH_AO22X4 U17519 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][3] ), .B(n17166), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][3] ), .D(
        n17400), .Z(n16557) );
  HS65_LH_AOI22X1 U17520 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][3] ), .B(n17392), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][3] ), .D(
        n17120), .Z(n16556) );
  HS65_LH_AOI22X1 U17521 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][3] ), .B(n17165), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[8][3] ), .D(
        n17394), .Z(n16555) );
  HS65_LH_NAND4ABX3 U17522 ( .A(n16558), .B(n16557), .C(n16556), .D(n16555), 
        .Z(n16561) );
  HS65_LH_AOI22X1 U17523 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][3] ), .B(n18124), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][3] ), .D(
        n17402), .Z(n16560) );
  HS65_LH_AOI22X1 U17524 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][3] ), .B(n17065), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][3] ), .D(
        n17148), .Z(n16559) );
  HS65_LH_NAND4ABX3 U17525 ( .A(n38440), .B(n16561), .C(n16560), .D(n16559), 
        .Z(n1794) );
  HS65_LH_AOI22X1 U17526 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][3] ), .B(n17383), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][3] ), .D(
        n17384), .Z(n16564) );
  HS65_LH_AOI22X1 U17527 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][3] ), .B(n17379), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][3] ), .D(
        n17130), .Z(n16563) );
  HS65_LH_NAND2X2 U17528 ( .A(n16564), .B(n16563), .Z(n16572) );
  HS65_LH_AO22X4 U17529 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][3] ), .B(n17377), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][3] ), .D(
        n17378), .Z(n16568) );
  HS65_LH_AO22X4 U17530 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][3] ), .B(n17177), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][3] ), .D(
        n17381), .Z(n16567) );
  HS65_LH_AOI22X1 U17531 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][3] ), .B(n17386), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][3] ), .D(
        n17382), .Z(n16566) );
  HS65_LH_AOI22X1 U17532 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][3] ), .B(n17564), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][3] ), .D(
        n17073), .Z(n16565) );
  HS65_LH_NAND4ABX3 U17533 ( .A(n16568), .B(n16567), .C(n16566), .D(n16565), 
        .Z(n16571) );
  HS65_LH_AOI22X1 U17534 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][3] ), .B(n17140), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][3] ), .D(
        n17191), .Z(n16570) );
  HS65_LH_AOI22X1 U17535 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][3] ), .B(n17562), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][3] ), .D(
        n17181), .Z(n16569) );
  HS65_LH_NAND4ABX3 U17536 ( .A(n16572), .B(n16571), .C(n16570), .D(n16569), 
        .Z(n1795) );
  HS65_LH_AOI22X1 U17537 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][4] ), .B(n17563), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][4] ), .D(
        n17403), .Z(n16574) );
  HS65_LH_AOI22X1 U17538 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][4] ), .B(n17404), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][4] ), .D(
        n17120), .Z(n16573) );
  HS65_LH_AO22X4 U17540 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][4] ), .B(n17148), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[8][4] ), .D(
        n17057), .Z(n16578) );
  HS65_LH_AO22X4 U17541 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][4] ), .B(n17400), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][4] ), .D(
        n17154), .Z(n16577) );
  HS65_LH_AOI22X1 U17542 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][4] ), .B(n17396), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][4] ), .D(
        n17397), .Z(n16576) );
  HS65_LH_AOI22X1 U17543 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][4] ), .B(n17065), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][4] ), .D(
        n17121), .Z(n16575) );
  HS65_LH_NAND4ABX3 U17544 ( .A(n16578), .B(n16577), .C(n16576), .D(n16575), 
        .Z(n16581) );
  HS65_LH_AOI22X1 U17545 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][4] ), .B(n17392), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][4] ), .D(
        n17165), .Z(n16580) );
  HS65_LH_AOI22X1 U17546 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][4] ), .B(n17166), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][4] ), .D(
        n17155), .Z(n16579) );
  HS65_LH_NAND4ABX3 U17547 ( .A(n16582), .B(n16581), .C(n38087), .D(n16579), 
        .Z(n1771) );
  HS65_LH_AOI22X1 U17548 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][4] ), .B(n17385), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][4] ), .D(
        n17100), .Z(n16584) );
  HS65_LH_AOI22X1 U17549 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][4] ), .B(n17181), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][4] ), .D(
        n17074), .Z(n16583) );
  HS65_LH_NAND2X2 U17550 ( .A(n16584), .B(n16583), .Z(n16592) );
  HS65_LH_AO22X4 U17551 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][4] ), .B(n17191), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][4] ), .D(
        n17073), .Z(n16588) );
  HS65_LH_AO22X4 U17552 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][4] ), .B(n17386), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[27][4] ), .D(
        n17177), .Z(n16587) );
  HS65_LH_AOI22X1 U17553 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][4] ), .B(n17179), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][4] ), .D(
        n17130), .Z(n16586) );
  HS65_LH_AOI22X1 U17554 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][4] ), .B(n17517), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][4] ), .D(
        n17180), .Z(n16585) );
  HS65_LH_NAND4ABX3 U17555 ( .A(n16588), .B(n16587), .C(n16586), .D(n16585), 
        .Z(n16591) );
  HS65_LH_AOI22X1 U17556 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][4] ), .B(n17564), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][4] ), .D(
        n17189), .Z(n16590) );
  HS65_LH_AOI22X1 U17557 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][4] ), .B(n17192), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][4] ), .D(
        n17141), .Z(n16589) );
  HS65_LH_AOI22X1 U17559 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][5] ), .B(n17399), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][5] ), .D(
        n17120), .Z(n16594) );
  HS65_LH_AOI22X1 U17560 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][5] ), .B(n21638), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][5] ), .D(
        n17149), .Z(n16593) );
  HS65_LH_AO22X4 U17562 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][5] ), .B(n17392), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][5] ), .D(
        n17404), .Z(n16598) );
  HS65_LH_AO22X4 U17563 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][5] ), .B(n17155), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][5] ), .D(
        n17400), .Z(n16597) );
  HS65_LH_AOI22X1 U17564 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][5] ), .B(n17057), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][5] ), .D(
        n17165), .Z(n16596) );
  HS65_LH_AOI22X1 U17565 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][5] ), .B(n17152), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][5] ), .D(
        n17154), .Z(n16595) );
  HS65_LH_NAND4ABX3 U17566 ( .A(n16598), .B(n16597), .C(n16596), .D(n16595), 
        .Z(n16601) );
  HS65_LH_AOI22X1 U17567 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][5] ), .B(n17391), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][5] ), .D(
        n17565), .Z(n16600) );
  HS65_LH_AOI22X1 U17568 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][5] ), .B(n17166), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][5] ), .D(
        n17065), .Z(n16599) );
  HS65_LH_NAND4ABX3 U17569 ( .A(n16602), .B(n16601), .C(n37249), .D(n16599), 
        .Z(n1748) );
  HS65_LH_AOI22X1 U17570 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][5] ), .B(n17192), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][5] ), .D(
        n17181), .Z(n16604) );
  HS65_LH_AOI22X1 U17571 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][5] ), .B(n17140), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][5] ), .D(
        n17382), .Z(n16603) );
  HS65_LH_NAND2X2 U17572 ( .A(n16604), .B(n16603), .Z(n16612) );
  HS65_LH_AO22X4 U17573 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][5] ), .B(n17516), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[17][5] ), .D(
        n17517), .Z(n16608) );
  HS65_LH_AO22X4 U17574 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][5] ), .B(n17379), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][5] ), .D(
        n17386), .Z(n16607) );
  HS65_LH_AOI22X1 U17575 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][5] ), .B(n17141), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][5] ), .D(
        n17189), .Z(n16606) );
  HS65_LH_AOI22X1 U17576 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][5] ), .B(n17387), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][5] ), .D(
        n17191), .Z(n16605) );
  HS65_LH_NAND4ABX3 U17577 ( .A(n16608), .B(n16607), .C(n16606), .D(n16605), 
        .Z(n16611) );
  HS65_LH_AOI22X1 U17578 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][5] ), .B(n17381), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][5] ), .D(
        n17073), .Z(n16610) );
  HS65_LH_AOI22X1 U17579 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][5] ), .B(n17074), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[27][5] ), .D(
        n17177), .Z(n16609) );
  HS65_LH_AOI22X1 U17581 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][6] ), .B(n17399), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][6] ), .D(
        n17040), .Z(n16614) );
  HS65_LH_AOI22X1 U17582 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][6] ), .B(n17563), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][6] ), .D(
        n17398), .Z(n16613) );
  HS65_LH_NAND2X2 U17583 ( .A(n16614), .B(n16613), .Z(n16622) );
  HS65_LH_AO22X4 U17584 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][6] ), .B(n17402), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][6] ), .D(
        n18124), .Z(n16618) );
  HS65_LH_AO22X4 U17585 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][6] ), .B(n17391), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][6] ), .D(
        n17404), .Z(n16617) );
  HS65_LH_BFX4 U17586 ( .A(n17392), .Z(n17157) );
  HS65_LH_AOI22X1 U17587 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][6] ), .B(n17157), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][6] ), .D(
        n17166), .Z(n16616) );
  HS65_LH_AOI22X1 U17588 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][6] ), .B(n18121), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[8][6] ), .D(
        n17394), .Z(n16615) );
  HS65_LH_NAND4ABX3 U17589 ( .A(n16618), .B(n16617), .C(n16616), .D(n16615), 
        .Z(n16621) );
  HS65_LH_AOI22X1 U17590 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][6] ), .B(n17152), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][6] ), .D(
        n17165), .Z(n16620) );
  HS65_LH_AOI22X1 U17591 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][6] ), .B(n17396), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][6] ), .D(
        n17149), .Z(n16619) );
  HS65_LH_NAND4ABX3 U17592 ( .A(n16622), .B(n16621), .C(n16620), .D(n16619), 
        .Z(n1725) );
  HS65_LH_AOI22X1 U17593 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][6] ), .B(n17189), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[17][6] ), .D(
        n17562), .Z(n16624) );
  HS65_LH_AOI22X1 U17594 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][6] ), .B(n17390), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][6] ), .D(
        n17180), .Z(n16623) );
  HS65_LH_NAND2X2 U17595 ( .A(n16624), .B(n16623), .Z(n16632) );
  HS65_LH_AO22X4 U17596 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][6] ), .B(n17192), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][6] ), .D(
        n17388), .Z(n16628) );
  HS65_LH_AO22X4 U17597 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][6] ), .B(n17141), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][6] ), .D(
        n17130), .Z(n16627) );
  HS65_LH_AOI22X1 U17598 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][6] ), .B(n17389), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[16][6] ), .D(
        n17564), .Z(n16626) );
  HS65_LH_AOI22X1 U17599 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][6] ), .B(n17140), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][6] ), .D(
        n17100), .Z(n16625) );
  HS65_LH_NAND4ABX3 U17600 ( .A(n16628), .B(n16627), .C(n16626), .D(n16625), 
        .Z(n16631) );
  HS65_LH_AOI22X1 U17601 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][6] ), .B(n17190), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][6] ), .D(
        n17191), .Z(n16630) );
  HS65_LH_AOI22X1 U17602 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][6] ), .B(n17383), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][6] ), .D(
        n17179), .Z(n16629) );
  HS65_LH_NAND4ABX3 U17603 ( .A(n16632), .B(n16631), .C(n16630), .D(n16629), 
        .Z(n1726) );
  HS65_LH_AOI22X1 U17604 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][7] ), .B(n18121), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][7] ), .D(
        n17402), .Z(n16634) );
  HS65_LH_AOI22X1 U17605 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][7] ), .B(n29623), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][7] ), .D(
        n17121), .Z(n16633) );
  HS65_LH_NAND2X2 U17606 ( .A(n16634), .B(n16633), .Z(n16642) );
  HS65_LH_AO22X4 U17607 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][7] ), .B(n17565), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[9][7] ), .D(
        n17396), .Z(n16638) );
  HS65_LH_AO22X4 U17608 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][7] ), .B(n17065), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][7] ), .D(
        n17165), .Z(n16637) );
  HS65_LH_AOI22X1 U17609 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][7] ), .B(n17393), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][7] ), .D(
        n17152), .Z(n16636) );
  HS65_LH_AOI22X1 U17610 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][7] ), .B(n17391), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][7] ), .D(
        n17397), .Z(n16635) );
  HS65_LH_NAND4ABX3 U17611 ( .A(n16638), .B(n16637), .C(n16636), .D(n16635), 
        .Z(n16641) );
  HS65_LH_AOI22X1 U17612 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][7] ), .B(n17057), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][7] ), .D(
        n17155), .Z(n16640) );
  HS65_LH_AOI22X1 U17613 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][7] ), .B(n17040), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][7] ), .D(
        n17157), .Z(n16639) );
  HS65_LH_NAND4ABX3 U17614 ( .A(n16642), .B(n16641), .C(n16640), .D(n16639), 
        .Z(n1702) );
  HS65_LH_AOI22X1 U17615 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][7] ), .B(n17381), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][7] ), .D(
        n17189), .Z(n16644) );
  HS65_LH_AOI22X1 U17616 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][7] ), .B(n17564), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[17][7] ), .D(
        n17562), .Z(n16643) );
  HS65_LH_NAND2X2 U17617 ( .A(n16644), .B(n16643), .Z(n16652) );
  HS65_LH_AO22X4 U17618 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][7] ), .B(n17141), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][7] ), .D(
        n17383), .Z(n16648) );
  HS65_LH_AO22X4 U17619 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][7] ), .B(n17379), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][7] ), .D(
        n17388), .Z(n16647) );
  HS65_LH_AOI22X1 U17620 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][7] ), .B(n17390), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][7] ), .D(
        n17190), .Z(n16646) );
  HS65_LH_AOI22X1 U17621 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][7] ), .B(n17387), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[31][7] ), .D(
        n17385), .Z(n16645) );
  HS65_LH_NAND4ABX3 U17622 ( .A(n16648), .B(n16647), .C(n16646), .D(n16645), 
        .Z(n16651) );
  HS65_LH_AOI22X1 U17623 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][7] ), .B(n17378), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][7] ), .D(
        n17382), .Z(n16650) );
  HS65_LH_AOI22X1 U17624 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][7] ), .B(n17191), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][7] ), .D(
        n17073), .Z(n16649) );
  HS65_LH_NAND4ABX3 U17625 ( .A(n16652), .B(n16651), .C(n16650), .D(n16649), 
        .Z(n1703) );
  HS65_LH_AOI22X1 U17626 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][8] ), .B(n17398), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][8] ), .D(
        n17403), .Z(n16654) );
  HS65_LH_AOI22X1 U17627 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][8] ), .B(n17563), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][8] ), .D(
        n17165), .Z(n16653) );
  HS65_LH_AO22X4 U17629 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][8] ), .B(n17154), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][8] ), .D(
        n17121), .Z(n16658) );
  HS65_LH_AO22X4 U17630 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][8] ), .B(n17057), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][8] ), .D(
        n17120), .Z(n16657) );
  HS65_LH_AOI22X1 U17631 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][8] ), .B(n17148), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][8] ), .D(
        n29623), .Z(n16656) );
  HS65_LH_AOI22X1 U17632 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][8] ), .B(n17040), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[9][8] ), .D(
        n21638), .Z(n16655) );
  HS65_LH_NAND4ABX3 U17633 ( .A(n16658), .B(n16657), .C(n16656), .D(n16655), 
        .Z(n16661) );
  HS65_LH_AOI22X1 U17634 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][8] ), .B(n17149), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][8] ), .D(
        n17155), .Z(n16660) );
  HS65_LH_AOI22X1 U17635 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][8] ), .B(n17157), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][8] ), .D(
        n17166), .Z(n16659) );
  HS65_LH_NAND4ABX3 U17636 ( .A(n33408), .B(n16661), .C(n16660), .D(n16659), 
        .Z(n1679) );
  HS65_LH_AOI22X1 U17637 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][8] ), .B(n17517), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[27][8] ), .D(
        n17390), .Z(n16664) );
  HS65_LH_AOI22X1 U17638 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][8] ), .B(n17379), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][8] ), .D(
        n17074), .Z(n16663) );
  HS65_LH_NAND2X2 U17639 ( .A(n16664), .B(n16663), .Z(n16672) );
  HS65_LH_AO22X4 U17640 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][8] ), .B(n17564), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][8] ), .D(
        n17381), .Z(n16668) );
  HS65_LH_AO22X4 U17641 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][8] ), .B(n17141), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][8] ), .D(
        n17377), .Z(n16667) );
  HS65_LH_AOI22X1 U17642 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][8] ), .B(n17389), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][8] ), .D(
        n17191), .Z(n16666) );
  HS65_LH_AOI22X1 U17643 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][8] ), .B(n17388), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][8] ), .D(
        n17190), .Z(n16665) );
  HS65_LH_NAND4ABX3 U17644 ( .A(n16668), .B(n16667), .C(n16666), .D(n16665), 
        .Z(n16671) );
  HS65_LH_AOI22X1 U17645 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][8] ), .B(n17387), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][8] ), .D(
        n17192), .Z(n16670) );
  HS65_LH_AOI22X1 U17646 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][8] ), .B(n17140), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][8] ), .D(
        n17179), .Z(n16669) );
  HS65_LH_NAND4ABX3 U17647 ( .A(n16672), .B(n16671), .C(n16670), .D(n16669), 
        .Z(n1680) );
  HS65_LH_AOI22X1 U17648 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][9] ), .B(n17057), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][9] ), .D(
        n17565), .Z(n16674) );
  HS65_LH_AOI22X1 U17649 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][9] ), .B(n17397), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][9] ), .D(
        n17166), .Z(n16673) );
  HS65_LH_AO22X4 U17651 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][9] ), .B(n17152), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][9] ), .D(
        n17398), .Z(n16678) );
  HS65_LH_AO22X4 U17652 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][9] ), .B(n17402), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][9] ), .D(
        n17404), .Z(n16677) );
  HS65_LH_AOI22X1 U17653 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][9] ), .B(n17165), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][9] ), .D(
        n17155), .Z(n16676) );
  HS65_LH_AOI22X1 U17654 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][9] ), .B(n17392), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][9] ), .D(
        n17120), .Z(n16675) );
  HS65_LH_NAND4ABX3 U17655 ( .A(n16678), .B(n16677), .C(n16676), .D(n16675), 
        .Z(n16681) );
  HS65_LH_AOI22X1 U17656 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][9] ), .B(n21638), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][9] ), .D(
        n17148), .Z(n16680) );
  HS65_LH_AOI22X1 U17657 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][9] ), .B(n17121), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][9] ), .D(
        n17040), .Z(n16679) );
  HS65_LH_NAND4ABX3 U17658 ( .A(n40989), .B(n16681), .C(n16680), .D(n16679), 
        .Z(n1656) );
  HS65_LH_AOI22X1 U17659 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][9] ), .B(n17390), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][9] ), .D(
        n17380), .Z(n16684) );
  HS65_LH_AOI22X1 U17660 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][9] ), .B(n17385), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][9] ), .D(
        n17190), .Z(n16683) );
  HS65_LH_NAND2X2 U17661 ( .A(n16684), .B(n16683), .Z(n16692) );
  HS65_LH_AO22X4 U17662 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][9] ), .B(n17181), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][9] ), .D(
        n17141), .Z(n16688) );
  HS65_LH_AO22X4 U17663 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][9] ), .B(n17517), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][9] ), .D(
        n17381), .Z(n16687) );
  HS65_LH_AOI22X1 U17664 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][9] ), .B(n17100), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[16][9] ), .D(
        n17564), .Z(n16686) );
  HS65_LH_AOI22X1 U17665 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][9] ), .B(n17383), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][9] ), .D(
        n17382), .Z(n16685) );
  HS65_LH_NAND4ABX3 U17666 ( .A(n16688), .B(n16687), .C(n16686), .D(n16685), 
        .Z(n16691) );
  HS65_LH_AOI22X1 U17667 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][9] ), .B(n17389), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][9] ), .D(
        n17189), .Z(n16690) );
  HS65_LH_AOI22X1 U17668 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][9] ), .B(n17387), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][9] ), .D(
        n17192), .Z(n16689) );
  HS65_LH_AOI22X1 U17670 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][10] ), .B(n29623), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][10] ), .D(
        n17398), .Z(n16694) );
  HS65_LH_AOI22X1 U17671 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][10] ), .B(n17396), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][10] ), .D(
        n17402), .Z(n16693) );
  HS65_LH_NAND2X2 U17672 ( .A(n16694), .B(n16693), .Z(n16702) );
  HS65_LH_AO22X4 U17673 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][10] ), .B(n17121), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][10] ), .D(n17148), 
        .Z(n16698) );
  HS65_LH_AO22X4 U17674 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][10] ), .B(n17155), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][10] ), .D(n17397), 
        .Z(n16697) );
  HS65_LH_AOI22X1 U17675 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][10] ), .B(n17393), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][10] ), .D(
        n17165), .Z(n16696) );
  HS65_LH_AOI22X1 U17676 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][10] ), .B(n17040), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[8][10] ), .D(n17394), 
        .Z(n16695) );
  HS65_LH_NAND4ABX3 U17677 ( .A(n16698), .B(n16697), .C(n16696), .D(n16695), 
        .Z(n16701) );
  HS65_LH_AOI22X1 U17678 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][10] ), .B(n17120), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][10] ), .D(
        n17157), .Z(n16700) );
  HS65_LH_AOI22X1 U17679 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][10] ), .B(n17563), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][10] ), .D(
        n17403), .Z(n16699) );
  HS65_LH_NAND4ABX3 U17680 ( .A(n16702), .B(n16701), .C(n16700), .D(n16699), 
        .Z(n1633) );
  HS65_LH_AOI22X1 U17681 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][10] ), .B(n17141), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[17][10] ), .D(n17562), 
        .Z(n16704) );
  HS65_LH_AOI22X1 U17682 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][10] ), .B(n17383), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[16][10] ), .D(n17564), 
        .Z(n16703) );
  HS65_LH_NAND2X2 U17683 ( .A(n16704), .B(n16703), .Z(n16712) );
  HS65_LH_AO22X4 U17684 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][10] ), .B(n17100), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][10] ), .D(n17189), 
        .Z(n16708) );
  HS65_LH_AO22X4 U17685 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][10] ), .B(n17192), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][10] ), .D(n17386), 
        .Z(n16707) );
  HS65_LH_AOI22X1 U17686 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][10] ), .B(n17179), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][10] ), .D(n17181), 
        .Z(n16706) );
  HS65_LH_AOI22X1 U17687 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][10] ), .B(n17387), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][10] ), .D(n17380), 
        .Z(n16705) );
  HS65_LH_NAND4ABX3 U17688 ( .A(n16708), .B(n16707), .C(n16706), .D(n16705), 
        .Z(n16711) );
  HS65_LH_AOI22X1 U17689 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][10] ), .B(n17140), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[27][10] ), .D(n17177), 
        .Z(n16710) );
  HS65_LH_AOI22X1 U17690 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][10] ), .B(n17180), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][10] ), .D(n17073), 
        .Z(n16709) );
  HS65_LH_NAND4ABX3 U17691 ( .A(n16712), .B(n16711), .C(n16710), .D(n16709), 
        .Z(n1634) );
  HS65_LH_AOI22X1 U17692 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][11] ), .B(n18121), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][11] ), .D(
        n17397), .Z(n16714) );
  HS65_LH_AOI22X1 U17693 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][11] ), .B(n17563), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[8][11] ), .D(
        n17057), .Z(n16713) );
  HS65_LH_NAND2X2 U17694 ( .A(n16714), .B(n16713), .Z(n16722) );
  HS65_LH_AO22X4 U17695 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][11] ), .B(n17065), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[9][11] ), .D(n17396), 
        .Z(n16718) );
  HS65_LH_AO22X4 U17696 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][11] ), .B(n17166), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][11] ), .D(
        n17392), .Z(n16717) );
  HS65_LH_AOI22X1 U17697 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][11] ), .B(n17148), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][11] ), .D(
        n17404), .Z(n16716) );
  HS65_LH_AOI22X1 U17698 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][11] ), .B(n18124), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][11] ), .D(n17399), 
        .Z(n16715) );
  HS65_LH_NAND4ABX3 U17699 ( .A(n16718), .B(n16717), .C(n16716), .D(n16715), 
        .Z(n16721) );
  HS65_LH_AOI22X1 U17700 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][11] ), .B(n17040), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][11] ), .D(n17403), 
        .Z(n16720) );
  HS65_LH_AOI22X1 U17701 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][11] ), .B(n17402), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][11] ), .D(
        n17165), .Z(n16719) );
  HS65_LH_NAND4ABX3 U17702 ( .A(n16722), .B(n16721), .C(n16720), .D(n16719), 
        .Z(n1610) );
  HS65_LH_AOI22X1 U17703 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][11] ), .B(n17192), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[31][11] ), .D(n17140), 
        .Z(n16724) );
  HS65_LH_AOI22X1 U17704 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][11] ), .B(n17383), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][11] ), .D(n17382), 
        .Z(n16723) );
  HS65_LH_NAND2X2 U17705 ( .A(n16724), .B(n16723), .Z(n16732) );
  HS65_LH_AO22X4 U17706 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][11] ), .B(n17562), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][11] ), .D(n17073), 
        .Z(n16728) );
  HS65_LH_AO22X4 U17707 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][11] ), .B(n17191), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][11] ), .D(n17130), 
        .Z(n16727) );
  HS65_LH_AOI22X1 U17708 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][11] ), .B(n17390), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][11] ), .D(n17181), 
        .Z(n16726) );
  HS65_LH_AOI22X1 U17709 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][11] ), .B(n17386), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[16][11] ), .D(n17564), 
        .Z(n16725) );
  HS65_LH_NAND4ABX3 U17710 ( .A(n16728), .B(n16727), .C(n16726), .D(n16725), 
        .Z(n16731) );
  HS65_LH_AOI22X1 U17711 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][11] ), .B(n17381), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][11] ), .D(n17100), 
        .Z(n16730) );
  HS65_LH_AOI22X1 U17712 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][11] ), .B(n17377), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][11] ), .D(n17384), 
        .Z(n16729) );
  HS65_LH_NAND4ABX3 U17713 ( .A(n16732), .B(n16731), .C(n16730), .D(n16729), 
        .Z(n1611) );
  HS65_LH_AOI22X1 U17714 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][12] ), .B(n18121), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][12] ), .D(
        n29623), .Z(n16734) );
  HS65_LH_AOI22X1 U17715 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][12] ), .B(n17399), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][12] ), .D(n17154), 
        .Z(n16733) );
  HS65_LH_NAND2X2 U17716 ( .A(n16734), .B(n16733), .Z(n16742) );
  HS65_LH_AO22X4 U17717 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][12] ), .B(n17401), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][12] ), .D(
        n17148), .Z(n16738) );
  HS65_LH_AO22X4 U17718 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][12] ), .B(n17157), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][12] ), .D(n17393), 
        .Z(n16737) );
  HS65_LH_AOI22X1 U17719 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][12] ), .B(n17403), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][12] ), .D(n17398), 
        .Z(n16736) );
  HS65_LH_AOI22X1 U17720 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][12] ), .B(n17400), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[8][12] ), .D(n17394), 
        .Z(n16735) );
  HS65_LH_NAND4ABX3 U17721 ( .A(n16738), .B(n16737), .C(n16736), .D(n16735), 
        .Z(n16741) );
  HS65_LH_AOI22X1 U17722 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][12] ), .B(n17149), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][12] ), .D(
        n17565), .Z(n16740) );
  HS65_LH_AOI22X1 U17723 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][12] ), .B(n17155), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[9][12] ), .D(n21638), 
        .Z(n16739) );
  HS65_LH_NAND4ABX3 U17724 ( .A(n16742), .B(n16741), .C(n16740), .D(n16739), 
        .Z(n1587) );
  HS65_LH_AOI22X1 U17725 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][12] ), .B(n17380), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[31][12] ), .D(n17140), 
        .Z(n16744) );
  HS65_LH_AOI22X1 U17726 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][12] ), .B(n17390), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][12] ), .D(n17190), 
        .Z(n16743) );
  HS65_LH_NAND2X2 U17727 ( .A(n16744), .B(n16743), .Z(n16752) );
  HS65_LH_AO22X4 U17728 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][12] ), .B(n17389), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][12] ), .D(n17141), 
        .Z(n16748) );
  HS65_LH_AO22X4 U17729 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][12] ), .B(n17387), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][12] ), .D(n17074), 
        .Z(n16747) );
  HS65_LH_AOI22X1 U17730 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][12] ), .B(n17100), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[17][12] ), .D(n17562), 
        .Z(n16746) );
  HS65_LH_AOI22X1 U17731 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][12] ), .B(n17382), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][12] ), .D(n17180), 
        .Z(n16745) );
  HS65_LH_NAND4ABX3 U17732 ( .A(n16748), .B(n16747), .C(n16746), .D(n16745), 
        .Z(n16751) );
  HS65_LH_AOI22X1 U17733 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][12] ), .B(n17377), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][12] ), .D(n17378), 
        .Z(n16750) );
  HS65_LH_AOI22X1 U17734 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][12] ), .B(n17181), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[16][12] ), .D(n17564), 
        .Z(n16749) );
  HS65_LH_AOI22X1 U17736 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][13] ), .B(n17401), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][13] ), .D(
        n17040), .Z(n16754) );
  HS65_LH_AOI22X1 U17737 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][13] ), .B(n17393), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][13] ), .D(
        n17121), .Z(n16753) );
  HS65_LH_NAND2X2 U17738 ( .A(n16754), .B(n16753), .Z(n16762) );
  HS65_LH_AO22X4 U17739 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][13] ), .B(n17402), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][13] ), .D(
        n18121), .Z(n16758) );
  HS65_LH_AO22X4 U17740 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][13] ), .B(n17404), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[8][13] ), .D(
        n17057), .Z(n16757) );
  HS65_LH_AOI22X1 U17741 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][13] ), .B(n17396), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][13] ), .D(
        n17157), .Z(n16756) );
  HS65_LH_AOI22X1 U17742 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][13] ), .B(n17563), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][13] ), .D(
        n17155), .Z(n16755) );
  HS65_LH_NAND4ABX3 U17743 ( .A(n16758), .B(n16757), .C(n16756), .D(n16755), 
        .Z(n16761) );
  HS65_LH_AOI22X1 U17744 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][13] ), .B(n17065), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][13] ), .D(n17403), 
        .Z(n16760) );
  HS65_LH_AOI22X1 U17745 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][13] ), .B(n17391), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][13] ), .D(
        n17149), .Z(n16759) );
  HS65_LH_NAND4ABX3 U17746 ( .A(n16762), .B(n16761), .C(n32843), .D(n16759), 
        .Z(n1564) );
  HS65_LH_AOI22X1 U17747 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][13] ), .B(n17389), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][13] ), .D(n17189), 
        .Z(n16764) );
  HS65_LH_AOI22X1 U17748 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][13] ), .B(n17177), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[16][13] ), .D(n17564), 
        .Z(n16763) );
  HS65_LH_NAND2X2 U17749 ( .A(n16764), .B(n16763), .Z(n16772) );
  HS65_LH_AO22X4 U17750 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][13] ), .B(n17517), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][13] ), .D(n17192), 
        .Z(n16768) );
  HS65_LH_AO22X4 U17751 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][13] ), .B(n17190), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[31][13] ), .D(n17140), 
        .Z(n16767) );
  HS65_LH_AOI22X1 U17752 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][13] ), .B(n17130), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][13] ), .D(n17074), 
        .Z(n16766) );
  HS65_LH_AOI22X1 U17753 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][13] ), .B(n17380), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][13] ), .D(n17100), 
        .Z(n16765) );
  HS65_LH_NAND4ABX3 U17754 ( .A(n16768), .B(n16767), .C(n16766), .D(n16765), 
        .Z(n16771) );
  HS65_LH_AOI22X1 U17755 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][13] ), .B(n17384), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][13] ), .D(n17179), 
        .Z(n16770) );
  HS65_LH_AOI22X1 U17756 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][13] ), .B(n17181), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][13] ), .D(n17180), 
        .Z(n16769) );
  HS65_LH_NAND4ABX3 U17757 ( .A(n16772), .B(n16771), .C(n16770), .D(n16769), 
        .Z(n1565) );
  HS65_LH_AOI22X1 U17758 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][14] ), .B(n17400), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][14] ), .D(n17120), 
        .Z(n16774) );
  HS65_LH_AOI22X1 U17759 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][14] ), .B(n17152), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][14] ), .D(n17155), 
        .Z(n16773) );
  HS65_LH_AO22X4 U17761 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][14] ), .B(n17401), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][14] ), .D(
        n17154), .Z(n16778) );
  HS65_LH_AO22X4 U17762 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][14] ), .B(n17391), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][14] ), .D(
        n17393), .Z(n16777) );
  HS65_LH_AOI22X1 U17763 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][14] ), .B(n17399), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][14] ), .D(n17157), 
        .Z(n16776) );
  HS65_LH_AOI22X1 U17764 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][14] ), .B(n17396), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][14] ), .D(
        n17565), .Z(n16775) );
  HS65_LH_NAND4ABX3 U17765 ( .A(n16778), .B(n16777), .C(n16776), .D(n16775), 
        .Z(n16781) );
  HS65_LH_AOI22X1 U17766 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][14] ), .B(n17065), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][14] ), .D(n17404), 
        .Z(n16780) );
  HS65_LH_AOI22X1 U17767 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][14] ), .B(n17149), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[8][14] ), .D(
        n17057), .Z(n16779) );
  HS65_LH_NAND4ABX3 U17768 ( .A(n16782), .B(n31796), .C(n31802), .D(n16779), 
        .Z(n1541) );
  HS65_LH_AOI22X1 U17769 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][14] ), .B(n17517), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][14] ), .D(n17073), 
        .Z(n16784) );
  HS65_LH_AOI22X1 U17770 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][14] ), .B(n17385), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][14] ), .D(n17180), 
        .Z(n16783) );
  HS65_LH_NAND2X2 U17771 ( .A(n16784), .B(n16783), .Z(n16792) );
  HS65_LH_AO22X4 U17772 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][14] ), .B(n17379), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[16][14] ), .D(n17516), 
        .Z(n16788) );
  HS65_LH_AO22X4 U17773 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][14] ), .B(n17192), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][14] ), .D(n17387), 
        .Z(n16787) );
  HS65_LH_AOI22X1 U17774 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][14] ), .B(n17377), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][14] ), .D(n17181), 
        .Z(n16786) );
  HS65_LH_AOI22X1 U17775 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][14] ), .B(n17177), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][14] ), .D(n17074), 
        .Z(n16785) );
  HS65_LH_NAND4ABX3 U17776 ( .A(n16788), .B(n16787), .C(n16786), .D(n16785), 
        .Z(n16791) );
  HS65_LH_AOI22X1 U17777 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][14] ), .B(n17179), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][14] ), .D(n17384), 
        .Z(n16790) );
  HS65_LH_AOI22X1 U17778 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][14] ), .B(n17191), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][14] ), .D(n17190), 
        .Z(n16789) );
  HS65_LH_AOI22X1 U17780 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][15] ), .B(n29623), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][15] ), .D(
        n17121), .Z(n16794) );
  HS65_LH_AOI22X1 U17781 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][15] ), .B(n17157), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][15] ), .D(n17398), 
        .Z(n16793) );
  HS65_LH_AO22X4 U17783 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][15] ), .B(n17393), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][15] ), .D(
        n17397), .Z(n16798) );
  HS65_LH_AO22X4 U17784 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][15] ), .B(n17563), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][15] ), .D(
        n18121), .Z(n16797) );
  HS65_LH_AOI22X1 U17785 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][15] ), .B(n17152), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][15] ), .D(n17148), 
        .Z(n16796) );
  HS65_LH_AOI22X1 U17786 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][15] ), .B(n17394), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][15] ), .D(
        n17154), .Z(n16795) );
  HS65_LH_AOI22X1 U17788 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][15] ), .B(n17396), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][15] ), .D(
        n17155), .Z(n16800) );
  HS65_LH_AOI22X1 U17789 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][15] ), .B(n17040), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][15] ), .D(n17165), 
        .Z(n16799) );
  HS65_LH_NAND4ABX3 U17790 ( .A(n16802), .B(n16801), .C(n16800), .D(n16799), 
        .Z(n1518) );
  HS65_LH_AOI22X1 U17791 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][15] ), .B(n17384), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][15] ), .D(n17130), 
        .Z(n16804) );
  HS65_LH_AOI22X1 U17792 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][15] ), .B(n17380), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][15] ), .D(n17382), 
        .Z(n16803) );
  HS65_LH_NAND2X2 U17793 ( .A(n16804), .B(n16803), .Z(n16812) );
  HS65_LH_AO22X4 U17794 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][15] ), .B(n17192), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][15] ), .D(n17381), 
        .Z(n16808) );
  HS65_LH_AO22X4 U17795 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][15] ), .B(n17140), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[16][15] ), .D(n17516), 
        .Z(n16807) );
  HS65_LH_AOI22X1 U17796 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][15] ), .B(n17383), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][15] ), .D(n17100), 
        .Z(n16806) );
  HS65_LH_AOI22X1 U17797 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][15] ), .B(n17390), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][15] ), .D(n17073), 
        .Z(n16805) );
  HS65_LH_NAND4ABX3 U17798 ( .A(n16808), .B(n16807), .C(n16806), .D(n16805), 
        .Z(n16811) );
  HS65_LH_AOI22X1 U17799 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][15] ), .B(n17388), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][15] ), .D(n17189), 
        .Z(n16810) );
  HS65_LH_AOI22X1 U17800 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][15] ), .B(n17190), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[17][15] ), .D(n17562), 
        .Z(n16809) );
  HS65_LH_AOI22X1 U17802 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][16] ), .B(n17394), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][16] ), .D(
        n17404), .Z(n16814) );
  HS65_LH_AOI22X1 U17803 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][16] ), .B(n17148), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][16] ), .D(
        n17154), .Z(n16813) );
  HS65_LH_AO22X4 U17805 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][16] ), .B(n17065), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][16] ), .D(n18124), 
        .Z(n16818) );
  HS65_LH_AO22X4 U17806 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][16] ), .B(n17040), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][16] ), .D(n17397), 
        .Z(n16817) );
  HS65_LH_AOI22X1 U17807 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][16] ), .B(n17121), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][16] ), .D(n17120), 
        .Z(n16816) );
  HS65_LH_AOI22X1 U17808 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][16] ), .B(n17152), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[9][16] ), .D(n17396), 
        .Z(n16815) );
  HS65_LH_NAND4ABX3 U17809 ( .A(n16818), .B(n16817), .C(n16816), .D(n16815), 
        .Z(n16821) );
  HS65_LH_AOI22X1 U17810 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][16] ), .B(n17157), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][16] ), .D(n17565), 
        .Z(n16820) );
  HS65_LH_AOI22X1 U17811 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][16] ), .B(n17166), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][16] ), .D(
        n17165), .Z(n16819) );
  HS65_LH_AOI22X1 U17813 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][16] ), .B(n17380), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][16] ), .D(n17189), 
        .Z(n16824) );
  HS65_LH_AOI22X1 U17814 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][16] ), .B(n17177), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][16] ), .D(n17190), 
        .Z(n16823) );
  HS65_LH_NAND2X2 U17815 ( .A(n16824), .B(n16823), .Z(n16832) );
  HS65_LH_AO22X4 U17816 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][16] ), .B(n17387), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][16] ), .D(n17073), 
        .Z(n16828) );
  HS65_LH_AO22X4 U17817 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][16] ), .B(n17379), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][16] ), .D(n17383), 
        .Z(n16827) );
  HS65_LH_AOI22X1 U17818 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][16] ), .B(n17388), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[17][16] ), .D(n17562), 
        .Z(n16826) );
  HS65_LH_AOI22X1 U17819 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][16] ), .B(n17384), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[16][16] ), .D(n17564), 
        .Z(n16825) );
  HS65_LH_NAND4ABX3 U17820 ( .A(n16828), .B(n16827), .C(n16826), .D(n16825), 
        .Z(n16831) );
  HS65_LH_AOI22X1 U17821 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][16] ), .B(n17140), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][16] ), .D(n17192), 
        .Z(n16830) );
  HS65_LH_AOI22X1 U17822 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][16] ), .B(n17180), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][16] ), .D(n17179), 
        .Z(n16829) );
  HS65_LH_NAND4ABX3 U17823 ( .A(n16832), .B(n16831), .C(n16830), .D(n16829), 
        .Z(n1496) );
  HS65_LH_AOI22X1 U17824 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][17] ), .B(n17565), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[8][17] ), .D(
        n17394), .Z(n16834) );
  HS65_LH_AOI22X1 U17825 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][17] ), .B(n17398), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[9][17] ), .D(n21638), 
        .Z(n16833) );
  HS65_LH_NAND2X2 U17826 ( .A(n16834), .B(n16833), .Z(n16842) );
  HS65_LH_AO22X4 U17827 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][17] ), .B(n17166), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][17] ), .D(
        n17154), .Z(n16838) );
  HS65_LH_AO22X4 U17828 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][17] ), .B(n17120), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][17] ), .D(
        n17148), .Z(n16837) );
  HS65_LH_AOI22X1 U17829 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][17] ), .B(n17157), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][17] ), .D(n29623), 
        .Z(n16836) );
  HS65_LH_AOI22X1 U17830 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][17] ), .B(n17400), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][17] ), .D(n17401), 
        .Z(n16835) );
  HS65_LH_NAND4ABX3 U17831 ( .A(n16838), .B(n16837), .C(n16836), .D(n16835), 
        .Z(n16841) );
  HS65_LH_AOI22X1 U17833 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][17] ), .B(n17155), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][17] ), .D(n17149), 
        .Z(n16839) );
  HS65_LH_NAND4ABX3 U17834 ( .A(n16842), .B(n16841), .C(n37115), .D(n16839), 
        .Z(n1472) );
  HS65_LH_AOI22X1 U17835 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][17] ), .B(n17384), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][17] ), .D(n17073), 
        .Z(n16844) );
  HS65_LH_AOI22X1 U17836 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][17] ), .B(n17385), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][17] ), .D(n17130), 
        .Z(n16843) );
  HS65_LH_NAND2X2 U17837 ( .A(n16844), .B(n16843), .Z(n16852) );
  HS65_LH_AO22X4 U17838 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][17] ), .B(n17190), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][17] ), .D(n17189), 
        .Z(n16848) );
  HS65_LH_AO22X4 U17839 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][17] ), .B(n17180), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][17] ), .D(n17100), 
        .Z(n16847) );
  HS65_LH_AOI22X1 U17840 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][17] ), .B(n17177), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][17] ), .D(n17382), 
        .Z(n16846) );
  HS65_LH_AOI22X1 U17841 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][17] ), .B(n17516), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[17][17] ), .D(n17562), 
        .Z(n16845) );
  HS65_LH_NAND4ABX3 U17842 ( .A(n16848), .B(n16847), .C(n16846), .D(n16845), 
        .Z(n16851) );
  HS65_LH_AOI22X1 U17843 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][17] ), .B(n17388), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][17] ), .D(n17192), 
        .Z(n16850) );
  HS65_LH_AOI22X1 U17844 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][17] ), .B(n17191), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][17] ), .D(n17074), 
        .Z(n16849) );
  HS65_LH_NAND4ABX3 U17845 ( .A(n16852), .B(n16851), .C(n16850), .D(n16849), 
        .Z(n1473) );
  HS65_LH_AOI22X1 U17846 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][18] ), .B(n17402), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][18] ), .D(
        n17121), .Z(n16854) );
  HS65_LH_AOI22X1 U17847 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][18] ), .B(n17396), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][18] ), .D(
        n17404), .Z(n16853) );
  HS65_LH_NAND2X2 U17848 ( .A(n16854), .B(n16853), .Z(n16862) );
  HS65_LH_AO22X4 U17849 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][18] ), .B(n17394), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][18] ), .D(
        n17152), .Z(n16858) );
  HS65_LH_AO22X4 U17850 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][18] ), .B(n17065), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][18] ), .D(n17392), 
        .Z(n16857) );
  HS65_LH_AOI22X1 U17851 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][18] ), .B(n17155), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][18] ), .D(n17397), 
        .Z(n16856) );
  HS65_LH_AOI22X1 U17852 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][18] ), .B(n17565), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][18] ), .D(
        n17040), .Z(n16855) );
  HS65_LH_NAND4ABX3 U17853 ( .A(n16858), .B(n16857), .C(n16856), .D(n16855), 
        .Z(n16861) );
  HS65_LH_AOI22X1 U17854 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][18] ), .B(n17401), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][18] ), .D(
        n17166), .Z(n16860) );
  HS65_LH_AOI22X1 U17855 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][18] ), .B(n17120), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][18] ), .D(
        n17148), .Z(n16859) );
  HS65_LH_NAND4ABX3 U17856 ( .A(n16862), .B(n16861), .C(n16860), .D(n16859), 
        .Z(n1449) );
  HS65_LH_AOI22X1 U17857 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][18] ), .B(n17190), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[31][18] ), .D(n17385), 
        .Z(n16864) );
  HS65_LH_AOI22X1 U17858 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][18] ), .B(n17180), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][18] ), .D(n17100), 
        .Z(n16863) );
  HS65_LH_NAND2X2 U17859 ( .A(n16864), .B(n16863), .Z(n16872) );
  HS65_LH_AO22X4 U17860 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][18] ), .B(n17564), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][18] ), .D(n17179), 
        .Z(n16868) );
  HS65_LH_AO22X4 U17861 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][18] ), .B(n17562), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][18] ), .D(n17073), 
        .Z(n16867) );
  HS65_LH_AOI22X1 U17862 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][18] ), .B(n17181), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][18] ), .D(n17378), 
        .Z(n16866) );
  HS65_LH_AOI22X1 U17863 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][18] ), .B(n17390), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][18] ), .D(n17384), 
        .Z(n16865) );
  HS65_LH_NAND4ABX3 U17864 ( .A(n16868), .B(n16867), .C(n16866), .D(n16865), 
        .Z(n16871) );
  HS65_LH_AOI22X1 U17865 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][18] ), .B(n17377), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][18] ), .D(n17074), 
        .Z(n16870) );
  HS65_LH_AOI22X1 U17866 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][18] ), .B(n17191), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][18] ), .D(n17130), 
        .Z(n16869) );
  HS65_LH_NAND4ABX3 U17867 ( .A(n16872), .B(n16871), .C(n16870), .D(n16869), 
        .Z(n1450) );
  HS65_LH_AOI22X1 U17868 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][19] ), .B(n17057), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][19] ), .D(
        n17399), .Z(n16874) );
  HS65_LH_AOI22X1 U17869 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][19] ), .B(n17152), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][19] ), .D(n17154), 
        .Z(n16873) );
  HS65_LH_NAND2X2 U17870 ( .A(n16874), .B(n16873), .Z(n16882) );
  HS65_LH_AO22X4 U17871 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][19] ), .B(n17400), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][19] ), .D(n17392), 
        .Z(n16878) );
  HS65_LH_AO22X4 U17872 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][19] ), .B(n17120), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][19] ), .D(
        n17148), .Z(n16877) );
  HS65_LH_AOI22X1 U17873 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][19] ), .B(n17404), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][19] ), .D(
        n17397), .Z(n16876) );
  HS65_LH_AOI22X1 U17874 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][19] ), .B(n17396), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][19] ), .D(
        n17166), .Z(n16875) );
  HS65_LH_NAND4ABX3 U17875 ( .A(n16878), .B(n16877), .C(n16876), .D(n16875), 
        .Z(n16881) );
  HS65_LH_AOI22X1 U17876 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][19] ), .B(n17401), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][19] ), .D(
        n17155), .Z(n16880) );
  HS65_LH_AOI22X1 U17877 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][19] ), .B(n17065), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][19] ), .D(n17565), 
        .Z(n16879) );
  HS65_LH_NAND4ABX3 U17878 ( .A(n16882), .B(n16881), .C(n16880), .D(n16879), 
        .Z(n1426) );
  HS65_LH_AOI22X1 U17879 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][19] ), .B(n17380), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][19] ), .D(n17074), 
        .Z(n16884) );
  HS65_LH_AOI22X1 U17880 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][19] ), .B(n17190), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][19] ), .D(n17189), 
        .Z(n16883) );
  HS65_LH_NAND2X2 U17881 ( .A(n16884), .B(n16883), .Z(n16892) );
  HS65_LH_AO22X4 U17882 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][19] ), .B(n17516), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][19] ), .D(n17073), 
        .Z(n16888) );
  HS65_LH_AO22X4 U17883 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][19] ), .B(n17388), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][19] ), .D(n17381), 
        .Z(n16887) );
  HS65_LH_AOI22X1 U17884 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][19] ), .B(n17562), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][19] ), .D(n17382), 
        .Z(n16886) );
  HS65_LH_AOI22X1 U17885 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][19] ), .B(n17390), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[31][19] ), .D(n17385), 
        .Z(n16885) );
  HS65_LH_NAND4ABX3 U17886 ( .A(n16888), .B(n16887), .C(n16886), .D(n16885), 
        .Z(n16891) );
  HS65_LH_AOI22X1 U17887 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][19] ), .B(n17379), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][19] ), .D(n17384), 
        .Z(n16890) );
  HS65_LH_AOI22X1 U17888 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][19] ), .B(n17378), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][19] ), .D(n17130), 
        .Z(n16889) );
  HS65_LH_NAND4ABX3 U17889 ( .A(n16892), .B(n16891), .C(n16890), .D(n16889), 
        .Z(n1427) );
  HS65_LH_AOI22X1 U17890 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][20] ), .B(n29623), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][20] ), .D(
        n17399), .Z(n16894) );
  HS65_LH_AOI22X1 U17891 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][20] ), .B(n17040), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][20] ), .D(n17154), 
        .Z(n16893) );
  HS65_LH_AO22X4 U17893 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][20] ), .B(n17065), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][20] ), .D(n17148), 
        .Z(n16898) );
  HS65_LH_AO22X4 U17894 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][20] ), .B(n17120), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][20] ), .D(
        n17149), .Z(n16897) );
  HS65_LH_AOI22X1 U17895 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][20] ), .B(n17057), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][20] ), .D(
        n17401), .Z(n16896) );
  HS65_LH_AOI22X1 U17896 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][20] ), .B(n18124), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[9][20] ), .D(n21638), 
        .Z(n16895) );
  HS65_LH_NAND4ABX3 U17897 ( .A(n16898), .B(n16897), .C(n16896), .D(n16895), 
        .Z(n16901) );
  HS65_LH_AOI22X1 U17898 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][20] ), .B(n17565), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][20] ), .D(
        n17403), .Z(n16900) );
  HS65_LH_AOI22X1 U17899 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][20] ), .B(n17157), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][20] ), .D(n17166), 
        .Z(n16899) );
  HS65_LH_AOI22X1 U17901 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][20] ), .B(n17180), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][20] ), .D(n17387), 
        .Z(n16904) );
  HS65_LH_AOI22X1 U17902 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][20] ), .B(n17179), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[27][20] ), .D(n17177), 
        .Z(n16903) );
  HS65_LH_NAND2X2 U17903 ( .A(n16904), .B(n16903), .Z(n16912) );
  HS65_LH_AO22X4 U17904 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][20] ), .B(n17389), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][20] ), .D(n17100), 
        .Z(n16908) );
  HS65_LH_AO22X4 U17905 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][20] ), .B(n17181), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][20] ), .D(n17377), 
        .Z(n16907) );
  HS65_LH_AOI22X1 U17906 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][20] ), .B(n17516), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[17][20] ), .D(n17562), 
        .Z(n16906) );
  HS65_LH_AOI22X1 U17907 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][20] ), .B(n17386), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[31][20] ), .D(n17385), 
        .Z(n16905) );
  HS65_LH_NAND4ABX3 U17908 ( .A(n16908), .B(n16907), .C(n16906), .D(n16905), 
        .Z(n16911) );
  HS65_LH_AOI22X1 U17909 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][20] ), .B(n17191), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][20] ), .D(n17192), 
        .Z(n16910) );
  HS65_LH_AOI22X1 U17910 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][20] ), .B(n17141), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][20] ), .D(n17074), 
        .Z(n16909) );
  HS65_LH_NAND4ABX3 U17911 ( .A(n16912), .B(n16911), .C(n16910), .D(n16909), 
        .Z(n1404) );
  HS65_LH_AOI22X1 U17912 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][21] ), .B(n17152), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[9][21] ), .D(n17396), 
        .Z(n16914) );
  HS65_LH_AOI22X1 U17913 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][21] ), .B(n17120), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][21] ), .D(
        n17040), .Z(n16913) );
  HS65_LH_NAND2X2 U17914 ( .A(n16914), .B(n16913), .Z(n16922) );
  HS65_LH_AO22X4 U17915 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][21] ), .B(n17121), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][21] ), .D(n18124), 
        .Z(n16918) );
  HS65_LH_AO22X4 U17916 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][21] ), .B(n17404), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][21] ), .D(
        n17165), .Z(n16917) );
  HS65_LH_AOI22X1 U17917 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][21] ), .B(n17065), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][21] ), .D(n17166), 
        .Z(n16916) );
  HS65_LH_AOI22X1 U17918 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][21] ), .B(n17392), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][21] ), .D(n17149), 
        .Z(n16915) );
  HS65_LH_NAND4ABX3 U17919 ( .A(n16918), .B(n16917), .C(n16916), .D(n16915), 
        .Z(n16921) );
  HS65_LH_AOI22X1 U17920 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][21] ), .B(n17563), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][21] ), .D(
        n17148), .Z(n16920) );
  HS65_LH_AOI22X1 U17921 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][21] ), .B(n17057), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][21] ), .D(
        n17154), .Z(n16919) );
  HS65_LH_NAND4ABX3 U17922 ( .A(n16922), .B(n16921), .C(n16920), .D(n16919), 
        .Z(n1380) );
  HS65_LH_AOI22X1 U17923 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][21] ), .B(n17388), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][21] ), .D(n17379), 
        .Z(n16924) );
  HS65_LH_AOI22X1 U17924 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][21] ), .B(n17179), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][21] ), .D(n17378), 
        .Z(n16923) );
  HS65_LH_NAND2X2 U17925 ( .A(n16924), .B(n16923), .Z(n16932) );
  HS65_LH_AO22X4 U17926 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][21] ), .B(n17073), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[27][21] ), .D(n17177), 
        .Z(n16928) );
  HS65_LH_AO22X4 U17927 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][21] ), .B(n17516), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[31][21] ), .D(n17140), 
        .Z(n16927) );
  HS65_LH_AOI22X1 U17928 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][21] ), .B(n17130), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][21] ), .D(n17180), 
        .Z(n16926) );
  HS65_LH_AOI22X1 U17929 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][21] ), .B(n17517), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][21] ), .D(n17191), 
        .Z(n16925) );
  HS65_LH_NAND4ABX3 U17930 ( .A(n16928), .B(n16927), .C(n16926), .D(n16925), 
        .Z(n16931) );
  HS65_LH_AOI22X1 U17931 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][21] ), .B(n17190), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][21] ), .D(n17074), 
        .Z(n16930) );
  HS65_LH_AOI22X1 U17932 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][21] ), .B(n17141), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][21] ), .D(n17377), 
        .Z(n16929) );
  HS65_LH_NAND4ABX3 U17933 ( .A(n16932), .B(n16931), .C(n16930), .D(n16929), 
        .Z(n1381) );
  HS65_LH_AOI22X1 U17934 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][22] ), .B(n18124), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[8][22] ), .D(n17394), 
        .Z(n16934) );
  HS65_LH_AOI22X1 U17935 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][22] ), .B(n17391), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][22] ), .D(
        n17154), .Z(n16933) );
  HS65_LH_AO22X4 U17937 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][22] ), .B(n17393), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][22] ), .D(
        n17565), .Z(n16938) );
  HS65_LH_AO22X4 U17938 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][22] ), .B(n17404), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][22] ), .D(
        n18121), .Z(n16937) );
  HS65_LH_AOI22X1 U17939 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][22] ), .B(n17403), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][22] ), .D(n17165), 
        .Z(n16936) );
  HS65_LH_AOI22X1 U17940 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][22] ), .B(n17399), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][22] ), .D(n17397), 
        .Z(n16935) );
  HS65_LH_NAND4ABX3 U17941 ( .A(n16938), .B(n16937), .C(n16936), .D(n16935), 
        .Z(n16941) );
  HS65_LH_AOI22X1 U17942 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][22] ), .B(n17040), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][22] ), .D(n17157), 
        .Z(n16940) );
  HS65_LH_AOI22X1 U17943 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][22] ), .B(n21638), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][22] ), .D(
        n17065), .Z(n16939) );
  HS65_LH_NAND4ABX3 U17944 ( .A(n37583), .B(n37652), .C(n16940), .D(n16939), 
        .Z(n1357) );
  HS65_LH_AOI22X1 U17945 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][22] ), .B(n17389), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[31][22] ), .D(n17385), 
        .Z(n16944) );
  HS65_LH_AOI22X1 U17946 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][22] ), .B(n17141), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[27][22] ), .D(n17177), 
        .Z(n16943) );
  HS65_LH_NAND2X2 U17947 ( .A(n16944), .B(n16943), .Z(n16952) );
  HS65_LH_AO22X4 U17948 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][22] ), .B(n17074), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][22] ), .D(n17130), 
        .Z(n16948) );
  HS65_LH_AO22X4 U17949 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][22] ), .B(n17191), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][22] ), .D(n17388), 
        .Z(n16947) );
  HS65_LH_AOI22X1 U17950 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][22] ), .B(n17386), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][22] ), .D(n17189), 
        .Z(n16946) );
  HS65_LH_AOI22X1 U17951 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][22] ), .B(n17381), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][22] ), .D(n17382), 
        .Z(n16945) );
  HS65_LH_NAND4ABX3 U17952 ( .A(n16948), .B(n16947), .C(n16946), .D(n16945), 
        .Z(n16951) );
  HS65_LH_AOI22X1 U17953 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][22] ), .B(n17379), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][22] ), .D(n17378), 
        .Z(n16950) );
  HS65_LH_AOI22X1 U17954 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][22] ), .B(n17564), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[17][22] ), .D(n17562), 
        .Z(n16949) );
  HS65_LH_NAND4ABX3 U17955 ( .A(n16952), .B(n16951), .C(n16950), .D(n16949), 
        .Z(n1358) );
  HS65_LH_AOI22X1 U17956 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][23] ), .B(n17399), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][23] ), .D(n17403), 
        .Z(n16954) );
  HS65_LH_AOI22X1 U17957 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][23] ), .B(n17149), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][23] ), .D(
        n18124), .Z(n16953) );
  HS65_LH_NAND2X2 U17958 ( .A(n16954), .B(n16953), .Z(n16962) );
  HS65_LH_AO22X4 U17959 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][23] ), .B(n17057), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][23] ), .D(
        n18121), .Z(n16958) );
  HS65_LH_AO22X4 U17960 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][23] ), .B(n17402), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][23] ), .D(
        n17563), .Z(n16957) );
  HS65_LH_AOI22X1 U17961 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][23] ), .B(n17400), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][23] ), .D(n17398), 
        .Z(n16956) );
  HS65_LH_AOI22X1 U17962 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][23] ), .B(n17391), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][23] ), .D(
        n17404), .Z(n16955) );
  HS65_LH_NAND4ABX3 U17963 ( .A(n16958), .B(n16957), .C(n16956), .D(n16955), 
        .Z(n16961) );
  HS65_LH_AOI22X1 U17964 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][23] ), .B(n17393), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][23] ), .D(
        n17401), .Z(n16960) );
  HS65_LH_AOI22X1 U17965 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][23] ), .B(n17392), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[9][23] ), .D(n21638), 
        .Z(n16959) );
  HS65_LH_NAND4ABX3 U17966 ( .A(n16962), .B(n16961), .C(n16960), .D(n16959), 
        .Z(n1334) );
  HS65_LH_AOI22X1 U17967 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][23] ), .B(n17516), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][23] ), .D(n17074), 
        .Z(n16964) );
  HS65_LH_AOI22X1 U17968 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][23] ), .B(n17380), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][23] ), .D(n17377), 
        .Z(n16963) );
  HS65_LH_NAND2X2 U17969 ( .A(n16964), .B(n16963), .Z(n16972) );
  HS65_LH_AO22X4 U17970 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][23] ), .B(n17140), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][23] ), .D(n17100), 
        .Z(n16968) );
  HS65_LH_AO22X4 U17971 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][23] ), .B(n17387), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][23] ), .D(n17141), 
        .Z(n16967) );
  HS65_LH_AOI22X1 U17972 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][23] ), .B(n17073), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][23] ), .D(n17378), 
        .Z(n16966) );
  HS65_LH_AOI22X1 U17973 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][23] ), .B(n17388), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][23] ), .D(n17180), 
        .Z(n16965) );
  HS65_LH_NAND4ABX3 U17974 ( .A(n16968), .B(n16967), .C(n16966), .D(n16965), 
        .Z(n16971) );
  HS65_LH_AOI22X1 U17975 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][23] ), .B(n17177), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][23] ), .D(n17190), 
        .Z(n16970) );
  HS65_LH_AOI22X1 U17976 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][23] ), .B(n17179), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[17][23] ), .D(n17562), 
        .Z(n16969) );
  HS65_LH_NAND4ABX3 U17977 ( .A(n16972), .B(n16971), .C(n16970), .D(n16969), 
        .Z(n1335) );
  HS65_LH_AOI22X1 U17978 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][24] ), .B(n17394), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[9][24] ), .D(
        n17396), .Z(n16974) );
  HS65_LH_AOI22X1 U17979 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][24] ), .B(n17397), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][24] ), .D(
        n17121), .Z(n16973) );
  HS65_LH_NAND2X2 U17980 ( .A(n16974), .B(n16973), .Z(n16982) );
  HS65_LH_AO22X4 U17981 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][24] ), .B(n17391), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][24] ), .D(
        n17154), .Z(n16978) );
  HS65_LH_AO22X4 U17982 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][24] ), .B(n17403), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][24] ), .D(n17165), 
        .Z(n16977) );
  HS65_LH_AOI22X1 U17983 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][24] ), .B(n17393), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][24] ), .D(
        n17040), .Z(n16976) );
  HS65_LH_AOI22X1 U17984 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][24] ), .B(n17404), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][24] ), .D(
        n17398), .Z(n16975) );
  HS65_LH_AOI22X1 U17986 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][24] ), .B(n17157), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][24] ), .D(n17565), 
        .Z(n16980) );
  HS65_LH_AOI22X1 U17987 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][24] ), .B(n17155), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][24] ), .D(n17120), 
        .Z(n16979) );
  HS65_LH_AOI22X1 U17989 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][24] ), .B(n17380), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][24] ), .D(n17179), 
        .Z(n16984) );
  HS65_LH_AOI22X1 U17990 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][24] ), .B(n17386), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][24] ), .D(n17180), 
        .Z(n16983) );
  HS65_LH_NAND2X2 U17991 ( .A(n16984), .B(n16983), .Z(n16992) );
  HS65_LH_AO22X4 U17992 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][24] ), .B(n17141), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][24] ), .D(n17074), 
        .Z(n16988) );
  HS65_LH_AO22X4 U17993 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][24] ), .B(n17564), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][24] ), .D(n17073), 
        .Z(n16987) );
  HS65_LH_AOI22X1 U17994 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][24] ), .B(n17140), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][24] ), .D(n17189), 
        .Z(n16986) );
  HS65_LH_AOI22X1 U17995 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][24] ), .B(n17130), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][24] ), .D(n17378), 
        .Z(n16985) );
  HS65_LH_NAND4ABX3 U17996 ( .A(n16988), .B(n16987), .C(n16986), .D(n16985), 
        .Z(n16991) );
  HS65_LH_AOI22X1 U17997 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][24] ), .B(n17517), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][24] ), .D(n17379), 
        .Z(n16990) );
  HS65_LH_AOI22X1 U17998 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][24] ), .B(n17177), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][24] ), .D(n17181), 
        .Z(n16989) );
  HS65_LH_AOI22X1 U18000 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][25] ), .B(n17393), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][25] ), .D(
        n29623), .Z(n16994) );
  HS65_LH_AOI22X1 U18001 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][25] ), .B(n17402), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][25] ), .D(
        n17398), .Z(n16993) );
  HS65_LH_NAND2X2 U18002 ( .A(n16994), .B(n16993), .Z(n17002) );
  HS65_LH_AO22X4 U18003 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][25] ), .B(n17149), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[8][25] ), .D(
        n17057), .Z(n16998) );
  HS65_LH_AO22X4 U18004 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][25] ), .B(n17157), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[9][25] ), .D(n17396), 
        .Z(n16997) );
  HS65_LH_AOI22X1 U18005 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][25] ), .B(n17400), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][25] ), .D(n17399), 
        .Z(n16996) );
  HS65_LH_AOI22X1 U18006 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][25] ), .B(n18121), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][25] ), .D(
        n17401), .Z(n16995) );
  HS65_LH_NAND4ABX3 U18007 ( .A(n16998), .B(n16997), .C(n16996), .D(n16995), 
        .Z(n17001) );
  HS65_LH_AOI22X1 U18008 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][25] ), .B(n18124), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][25] ), .D(n17403), 
        .Z(n17000) );
  HS65_LH_AOI22X1 U18009 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][25] ), .B(n17563), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][25] ), .D(
        n17148), .Z(n16999) );
  HS65_LH_AOI22X1 U18011 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][25] ), .B(n17384), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][25] ), .D(n17377), 
        .Z(n17004) );
  HS65_LH_AOI22X1 U18012 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][25] ), .B(n17389), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][25] ), .D(n17179), 
        .Z(n17003) );
  HS65_LH_NAND2X2 U18013 ( .A(n17004), .B(n17003), .Z(n17012) );
  HS65_LH_AO22X4 U18014 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][25] ), .B(n17100), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][25] ), .D(n17130), 
        .Z(n17008) );
  HS65_LH_AO22X4 U18015 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][25] ), .B(n17388), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][25] ), .D(n17386), 
        .Z(n17007) );
  HS65_LH_AOI22X1 U18016 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][25] ), .B(n17516), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][25] ), .D(n17378), 
        .Z(n17006) );
  HS65_LH_AOI22X1 U18017 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][25] ), .B(n17385), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[17][25] ), .D(n17562), 
        .Z(n17005) );
  HS65_LH_NAND4ABX3 U18018 ( .A(n17008), .B(n17007), .C(n17006), .D(n17005), 
        .Z(n17011) );
  HS65_LH_AOI22X1 U18019 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][25] ), .B(n17180), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][25] ), .D(n17074), 
        .Z(n17010) );
  HS65_LH_AOI22X1 U18020 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][25] ), .B(n17177), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][25] ), .D(n17191), 
        .Z(n17009) );
  HS65_LH_NAND4ABX3 U18021 ( .A(n17012), .B(n17011), .C(n17010), .D(n17009), 
        .Z(n1289) );
  HS65_LH_AOI22X1 U18022 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][26] ), .B(n17391), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][26] ), .D(
        n17399), .Z(n17014) );
  HS65_LH_AOI22X1 U18023 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][26] ), .B(n17152), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][26] ), .D(n17166), 
        .Z(n17013) );
  HS65_LH_NAND2X2 U18024 ( .A(n17014), .B(n17013), .Z(n17022) );
  HS65_LH_AO22X4 U18025 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][26] ), .B(n17157), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[8][26] ), .D(n17057), 
        .Z(n17018) );
  HS65_LH_AO22X4 U18026 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][26] ), .B(n17165), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[9][26] ), .D(
        n17396), .Z(n17017) );
  HS65_LH_AOI22X1 U18027 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][26] ), .B(n18121), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][26] ), .D(
        n17155), .Z(n17016) );
  HS65_LH_AOI22X1 U18028 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][26] ), .B(n17563), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][26] ), .D(
        n17149), .Z(n17015) );
  HS65_LH_NAND4ABX3 U18029 ( .A(n17018), .B(n17017), .C(n17016), .D(n17015), 
        .Z(n17021) );
  HS65_LH_AOI22X1 U18030 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][26] ), .B(n17065), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][26] ), .D(n17040), 
        .Z(n17020) );
  HS65_LH_AOI22X1 U18031 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][26] ), .B(n29623), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][26] ), .D(
        n17402), .Z(n17019) );
  HS65_LH_NAND4ABX3 U18032 ( .A(n17022), .B(n17021), .C(n17020), .D(n38228), 
        .Z(n1265) );
  HS65_LH_AOI22X1 U18033 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][26] ), .B(n17383), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[27][26] ), .D(n17390), 
        .Z(n17024) );
  HS65_LH_AOI22X1 U18034 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][26] ), .B(n17384), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][26] ), .D(n17073), 
        .Z(n17023) );
  HS65_LH_NAND2X2 U18035 ( .A(n17024), .B(n17023), .Z(n17032) );
  HS65_LH_AO22X4 U18036 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][26] ), .B(n17517), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[26][26] ), .D(n17381), 
        .Z(n17028) );
  HS65_LH_AO22X4 U18037 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][26] ), .B(n17516), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[31][26] ), .D(n17140), 
        .Z(n17027) );
  HS65_LH_AOI22X1 U18038 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][26] ), .B(n17386), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][26] ), .D(n17100), 
        .Z(n17026) );
  HS65_LH_AOI22X1 U18039 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][26] ), .B(n17387), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][26] ), .D(n17382), 
        .Z(n17025) );
  HS65_LH_NAND4ABX3 U18040 ( .A(n17028), .B(n17027), .C(n17026), .D(n17025), 
        .Z(n17031) );
  HS65_LH_AOI22X1 U18041 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][26] ), .B(n17191), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][26] ), .D(n17377), 
        .Z(n17030) );
  HS65_LH_AOI22X1 U18042 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][26] ), .B(n17181), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][26] ), .D(n17192), 
        .Z(n17029) );
  HS65_LH_AOI22X1 U18044 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][27] ), .B(n17404), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][27] ), .D(
        n17157), .Z(n17034) );
  HS65_LH_AOI22X1 U18045 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][27] ), .B(n17401), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][27] ), .D(
        n17166), .Z(n17033) );
  HS65_LH_NAND2X2 U18046 ( .A(n17034), .B(n17033), .Z(n17044) );
  HS65_LH_AO22X4 U18047 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][27] ), .B(n17396), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][27] ), .D(
        n17154), .Z(n17039) );
  HS65_LH_AO22X4 U18048 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][27] ), .B(n17152), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][27] ), .D(n17149), 
        .Z(n17038) );
  HS65_LH_AOI22X1 U18049 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][27] ), .B(n18124), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[8][27] ), .D(n17394), 
        .Z(n17037) );
  HS65_LH_AOI22X1 U18050 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][27] ), .B(n17391), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][27] ), .D(
        n17565), .Z(n17036) );
  HS65_LH_NAND4ABX3 U18051 ( .A(n17039), .B(n17038), .C(n17037), .D(n17036), 
        .Z(n17043) );
  HS65_LH_AOI22X1 U18053 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][27] ), .B(n17040), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][27] ), .D(n17121), 
        .Z(n17041) );
  HS65_LH_NAND4ABX3 U18054 ( .A(n17044), .B(n17043), .C(n37922), .D(n17041), 
        .Z(n1242) );
  HS65_LH_AOI22X1 U18055 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][27] ), .B(n17381), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][27] ), .D(n17382), 
        .Z(n17047) );
  HS65_LH_AOI22X1 U18056 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][27] ), .B(n17390), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][27] ), .D(n17130), 
        .Z(n17046) );
  HS65_LH_NAND2X2 U18057 ( .A(n17047), .B(n17046), .Z(n17056) );
  HS65_LH_AO22X4 U18058 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][27] ), .B(n17386), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][27] ), .D(n17189), 
        .Z(n17052) );
  HS65_LH_AO22X4 U18059 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][27] ), .B(n17191), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][27] ), .D(n17383), 
        .Z(n17051) );
  HS65_LH_AOI22X1 U18060 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][27] ), .B(n17073), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[17][27] ), .D(n17562), 
        .Z(n17050) );
  HS65_LH_AOI22X1 U18061 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][27] ), .B(n17388), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][27] ), .D(n17378), 
        .Z(n17049) );
  HS65_LH_NAND4ABX3 U18062 ( .A(n17052), .B(n17051), .C(n17050), .D(n17049), 
        .Z(n17055) );
  HS65_LH_AOI22X1 U18063 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][27] ), .B(n17140), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[16][27] ), .D(n17564), 
        .Z(n17054) );
  HS65_LH_AOI22X1 U18064 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][27] ), .B(n17141), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][27] ), .D(n17100), 
        .Z(n17053) );
  HS65_LH_NAND4ABX3 U18065 ( .A(n17056), .B(n17055), .C(n17054), .D(n17053), 
        .Z(n1243) );
  HS65_LH_AOI22X1 U18066 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][28] ), .B(n17400), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][28] ), .D(n17401), 
        .Z(n17059) );
  HS65_LH_AOI22X1 U18067 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][28] ), .B(n17057), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][28] ), .D(
        n17404), .Z(n17058) );
  HS65_LH_AO22X4 U18069 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][28] ), .B(n17393), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][28] ), .D(
        n17563), .Z(n17064) );
  HS65_LH_AO22X4 U18070 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][28] ), .B(n18124), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][28] ), .D(n17392), 
        .Z(n17063) );
  HS65_LH_AOI22X1 U18071 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][28] ), .B(n17397), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][28] ), .D(
        n17154), .Z(n17062) );
  HS65_LH_AOI22X1 U18072 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][28] ), .B(n18121), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[9][28] ), .D(
        n17396), .Z(n17061) );
  HS65_LH_NAND4ABX3 U18073 ( .A(n17064), .B(n17063), .C(n17062), .D(n17061), 
        .Z(n17069) );
  HS65_LH_AOI22X1 U18074 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][28] ), .B(n17391), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][28] ), .D(
        n17065), .Z(n17068) );
  HS65_LH_AOI22X1 U18075 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][28] ), .B(n17121), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][28] ), .D(n17403), 
        .Z(n17067) );
  HS65_LH_AOI22X1 U18077 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][28] ), .B(n17381), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][28] ), .D(n17378), 
        .Z(n17072) );
  HS65_LH_AOI22X1 U18078 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][28] ), .B(n17386), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][28] ), .D(n17181), 
        .Z(n17071) );
  HS65_LH_AO22X4 U18080 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][28] ), .B(n17073), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][28] ), .D(n17179), 
        .Z(n17078) );
  HS65_LH_AO22X4 U18081 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][28] ), .B(n17074), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[27][28] ), .D(n17177), 
        .Z(n17077) );
  HS65_LH_AOI22X1 U18082 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][28] ), .B(n17516), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][28] ), .D(n17189), 
        .Z(n17076) );
  HS65_LH_AOI22X1 U18083 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][28] ), .B(n17517), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][28] ), .D(n17379), 
        .Z(n17075) );
  HS65_LH_NAND4ABX3 U18084 ( .A(n17078), .B(n17077), .C(n17076), .D(n17075), 
        .Z(n17081) );
  HS65_LH_AOI22X1 U18085 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][28] ), .B(n17191), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][28] ), .D(n17130), 
        .Z(n17080) );
  HS65_LH_AOI22X1 U18086 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][28] ), .B(n17141), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[31][28] ), .D(n17140), 
        .Z(n17079) );
  HS65_LH_NAND4ABX3 U18087 ( .A(n17082), .B(n17081), .C(n17080), .D(n17079), 
        .Z(n1220) );
  HS65_LH_AOI22X1 U18088 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][29] ), .B(n17393), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[8][29] ), .D(
        n17394), .Z(n17085) );
  HS65_LH_AOI22X1 U18089 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][29] ), .B(n17563), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][29] ), .D(
        n17404), .Z(n17084) );
  HS65_LH_NAND2X2 U18090 ( .A(n17085), .B(n17084), .Z(n17096) );
  HS65_LH_AO22X4 U18091 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][29] ), .B(n17149), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][29] ), .D(
        n17152), .Z(n17089) );
  HS65_LH_AO22X4 U18092 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][29] ), .B(n17396), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][29] ), .D(
        n17400), .Z(n17088) );
  HS65_LH_AOI22X1 U18093 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][29] ), .B(n17398), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][29] ), .D(n17401), 
        .Z(n17087) );
  HS65_LH_AOI22X1 U18094 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][29] ), .B(n18121), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][29] ), .D(
        n17157), .Z(n17086) );
  HS65_LH_NAND4ABX3 U18095 ( .A(n17089), .B(n17088), .C(n17087), .D(n17086), 
        .Z(n17095) );
  HS65_LH_AOI22X1 U18096 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][29] ), .B(n18124), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][29] ), .D(n17402), 
        .Z(n17094) );
  HS65_LH_AOI22X1 U18097 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][29] ), .B(n17391), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][29] ), .D(
        n17121), .Z(n17093) );
  HS65_LH_AOI22X1 U18099 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][29] ), .B(n17564), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][29] ), .D(n17380), 
        .Z(n17099) );
  HS65_LH_AOI22X1 U18100 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][29] ), .B(n17141), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[17][29] ), .D(n17517), 
        .Z(n17098) );
  HS65_LH_NAND2X2 U18101 ( .A(n17099), .B(n17098), .Z(n17109) );
  HS65_LH_AO22X4 U18102 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][29] ), .B(n17100), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][29] ), .D(n17189), 
        .Z(n17105) );
  HS65_LH_AO22X4 U18103 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][29] ), .B(n17181), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][29] ), .D(n17130), 
        .Z(n17104) );
  HS65_LH_AOI22X1 U18104 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][29] ), .B(n17180), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][29] ), .D(n17382), 
        .Z(n17103) );
  HS65_LH_AOI22X1 U18105 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][29] ), .B(n17383), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[31][29] ), .D(n17385), 
        .Z(n17102) );
  HS65_LH_NAND4ABX3 U18106 ( .A(n17105), .B(n17104), .C(n17103), .D(n17102), 
        .Z(n17108) );
  HS65_LH_AOI22X1 U18107 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][29] ), .B(n17389), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[27][29] ), .D(n17177), 
        .Z(n17107) );
  HS65_LH_AOI22X1 U18108 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][29] ), .B(n17190), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][29] ), .D(n17192), 
        .Z(n17106) );
  HS65_LH_AOI22X1 U18110 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][30] ), .B(n21638), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][30] ), .D(
        n17148), .Z(n17113) );
  HS65_LH_AOI22X1 U18111 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][30] ), .B(n17392), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][30] ), .D(n17155), 
        .Z(n17112) );
  HS65_LH_NAND2X2 U18112 ( .A(n17113), .B(n17112), .Z(n17126) );
  HS65_LH_AO22X4 U18113 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][30] ), .B(n17401), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][30] ), .D(
        n17154), .Z(n17119) );
  HS65_LH_AO22X4 U18114 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][30] ), .B(n17400), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][30] ), .D(n17152), 
        .Z(n17118) );
  HS65_LH_AOI22X1 U18115 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][30] ), .B(n17398), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[8][30] ), .D(n17394), 
        .Z(n17117) );
  HS65_LH_AOI22X1 U18116 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][30] ), .B(n17404), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][30] ), .D(
        n17166), .Z(n17116) );
  HS65_LH_NAND4ABX3 U18117 ( .A(n17119), .B(n17118), .C(n17117), .D(n17116), 
        .Z(n17125) );
  HS65_LH_AOI22X1 U18118 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][30] ), .B(n17120), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[3][30] ), .D(
        n17149), .Z(n17124) );
  HS65_LH_AOI22X1 U18119 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][30] ), .B(n17563), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][30] ), .D(
        n17121), .Z(n17123) );
  HS65_LH_NAND4ABX3 U18120 ( .A(n17126), .B(n17125), .C(n17124), .D(n17123), 
        .Z(n1173) );
  HS65_LH_AOI22X1 U18121 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][30] ), .B(n17516), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][30] ), .D(n17181), 
        .Z(n17129) );
  HS65_LH_AOI22X1 U18122 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][30] ), .B(n17377), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[27][30] ), .D(n17177), 
        .Z(n17128) );
  HS65_LH_NAND2X2 U18123 ( .A(n17129), .B(n17128), .Z(n17145) );
  HS65_LH_AO22X4 U18124 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][30] ), .B(n17517), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[24][30] ), .D(n17130), 
        .Z(n17138) );
  HS65_LH_AO22X4 U18125 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][30] ), .B(n17179), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[18][30] ), .D(n17386), 
        .Z(n17137) );
  HS65_LH_AOI22X1 U18126 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][30] ), .B(n17389), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][30] ), .D(n17383), 
        .Z(n17136) );
  HS65_LH_AOI22X1 U18127 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][30] ), .B(n17381), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][30] ), .D(n17380), 
        .Z(n17135) );
  HS65_LH_NAND4ABX3 U18128 ( .A(n17138), .B(n17137), .C(n17136), .D(n17135), 
        .Z(n17144) );
  HS65_LH_AOI22X1 U18129 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][30] ), .B(n17378), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][30] ), .D(n17379), 
        .Z(n17143) );
  HS65_LH_AOI22X1 U18130 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][30] ), .B(n17141), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[31][30] ), .D(n17140), 
        .Z(n17142) );
  HS65_LH_NAND4ABX3 U18131 ( .A(n17145), .B(n17144), .C(n17143), .D(n17142), 
        .Z(n1174) );
  HS65_LH_AOI22X1 U18132 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][31] ), .B(n17400), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[8][31] ), .D(n17394), 
        .Z(n17151) );
  HS65_LH_AOI22X1 U18133 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][31] ), .B(n17149), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][31] ), .D(
        n17148), .Z(n17150) );
  HS65_LH_NAND2X2 U18134 ( .A(n17151), .B(n17150), .Z(n17170) );
  HS65_LH_AO22X4 U18135 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][31] ), .B(n29623), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][31] ), .D(
        n17152), .Z(n17162) );
  HS65_LH_AO22X4 U18136 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][31] ), .B(n17565), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][31] ), .D(
        n17154), .Z(n17161) );
  HS65_LH_AOI22X1 U18137 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][31] ), .B(n17398), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][31] ), .D(n17155), 
        .Z(n17160) );
  HS65_LH_AOI22X1 U18138 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][31] ), .B(n17399), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][31] ), .D(n17157), 
        .Z(n17159) );
  HS65_LH_AOI22X1 U18140 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][31] ), .B(n18121), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[9][31] ), .D(
        n21638), .Z(n17168) );
  HS65_LH_AOI22X1 U18141 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][31] ), .B(n17166), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][31] ), .D(
        n17165), .Z(n17167) );
  HS65_LH_NAND4ABX3 U18142 ( .A(n17170), .B(n17169), .C(n40976), .D(n17167), 
        .Z(n1150) );
  HS65_LH_AOI22X1 U18143 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][31] ), .B(n17379), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[31][31] ), .D(n17385), 
        .Z(n17176) );
  HS65_LH_AOI22X1 U18144 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][31] ), .B(n17387), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][31] ), .D(n17384), 
        .Z(n17175) );
  HS65_LH_NAND2X2 U18145 ( .A(n17176), .B(n17175), .Z(n17196) );
  HS65_LH_AO22X4 U18146 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][31] ), .B(n17389), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[27][31] ), .D(n17177), 
        .Z(n17188) );
  HS65_LH_AO22X4 U18147 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][31] ), .B(n17180), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][31] ), .D(n17179), 
        .Z(n17187) );
  HS65_LH_AOI22X1 U18148 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][31] ), .B(n17516), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][31] ), .D(n17181), 
        .Z(n17186) );
  HS65_LH_AOI22X1 U18149 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][31] ), .B(n17383), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[17][31] ), .D(n17562), 
        .Z(n17185) );
  HS65_LH_NAND4ABX3 U18150 ( .A(n17188), .B(n17187), .C(n17186), .D(n17185), 
        .Z(n17195) );
  HS65_LH_AOI22X1 U18151 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][31] ), .B(n17190), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][31] ), .D(n17189), 
        .Z(n17194) );
  HS65_LH_AOI22X1 U18152 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][31] ), .B(n17192), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][31] ), .D(n17191), 
        .Z(n17193) );
  HS65_LH_NAND4ABX3 U18153 ( .A(n17196), .B(n17195), .C(n17194), .D(n17193), 
        .Z(n1151) );
  HS65_LH_NOR2X2 U18154 ( .A(n9284), .B(n13893), .Z(n17199) );
  HS65_LH_MX41X4 U18155 ( .D0(n17313), .S0(Data_out_fromRAM[8]), .D1(
        Data_out_fromRAM[24]), .S1(n17505), .D2(Data_out_fromRAM[16]), .S2(
        n17376), .D3(n17454), .S3(Data_out_fromRAM[0]), .Z(n338) );
  HS65_LH_MX41X4 U18156 ( .D0(n17313), .S0(Data_out_fromRAM[9]), .D1(n17376), 
        .S1(Data_out_fromRAM[17]), .D2(Data_out_fromRAM[25]), .S2(n17505), 
        .D3(Data_out_fromRAM[1]), .S3(n17454), .Z(n330) );
  HS65_LH_MX41X4 U18157 ( .D0(n17313), .S0(Data_out_fromRAM[10]), .D1(n17376), 
        .S1(Data_out_fromRAM[18]), .D2(Data_out_fromRAM[26]), .S2(n17505), 
        .D3(n17454), .S3(Data_out_fromRAM[2]), .Z(n329) );
  HS65_LH_MX41X4 U18158 ( .D0(n17313), .S0(Data_out_fromRAM[11]), .D1(n17376), 
        .S1(Data_out_fromRAM[19]), .D2(Data_out_fromRAM[27]), .S2(n17505), 
        .D3(Data_out_fromRAM[3]), .S3(n17454), .Z(n328) );
  HS65_LH_MX41X4 U18159 ( .D0(n17313), .S0(Data_out_fromRAM[12]), .D1(n17376), 
        .S1(Data_out_fromRAM[20]), .D2(Data_out_fromRAM[4]), .S2(n17454), .D3(
        Data_out_fromRAM[28]), .S3(n17505), .Z(n327) );
  HS65_LH_MX41X4 U18160 ( .D0(n17313), .S0(Data_out_fromRAM[13]), .D1(n17376), 
        .S1(Data_out_fromRAM[21]), .D2(Data_out_fromRAM[5]), .S2(n17454), .D3(
        Data_out_fromRAM[29]), .S3(n17505), .Z(n326) );
  HS65_LH_MX41X4 U18161 ( .D0(n17313), .S0(Data_out_fromRAM[14]), .D1(n17376), 
        .S1(Data_out_fromRAM[22]), .D2(Data_out_fromRAM[30]), .S2(n17505), 
        .D3(Data_out_fromRAM[6]), .S3(n17454), .Z(n325) );
  HS65_LH_MX41X4 U18162 ( .D0(n17313), .S0(Data_out_fromRAM[15]), .D1(n17376), 
        .S1(Data_out_fromRAM[23]), .D2(n17454), .S2(Data_out_fromRAM[7]), .D3(
        Data_out_fromRAM[31]), .S3(n17505), .Z(n324) );
  HS65_LH_NAND2X2 U18163 ( .A(n11649), .B(n11644), .Z(n17200) );
  HS65_LH_NAND4ABX3 U18164 ( .A(n11651), .B(n17200), .C(n274), .D(n1103), .Z(
        n276) );
  HS65_LH_NAND2X2 U18165 ( .A(n17203), .B(n15470), .Z(n17201) );
  HS65_LH_OAI21X2 U18166 ( .A(n17446), .B(n17304), .C(n17375), .Z(n17206) );
  HS65_LH_NOR2AX3 U18167 ( .A(n17210), .B(n17209), .Z(n218) );
  HS65_LH_NOR2AX3 U18168 ( .A(n15749), .B(n258), .Z(n179) );
  HS65_LL_DFPHQX4 clk_r_REG261_S1 ( .D(n3901), .E(\u_DataPath/u_fetch/pc1/N3 ), 
        .CP(clk), .Q(n18039) );
  HS65_LL_DFPHQX4 clk_r_REG225_S1 ( .D(n4107), .E(\u_DataPath/u_fetch/pc1/N3 ), 
        .CP(clk), .Q(n18029) );
  HS65_LL_DFPHQX4 clk_r_REG451_S1 ( .D(n4217), .E(\u_DataPath/u_fetch/pc1/N3 ), 
        .CP(clk), .Q(n18021) );
  HS65_LL_DFPHQX4 clk_r_REG198_S1 ( .D(n12672), .E(\u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n17685) );
  HS65_LL_DFPHQX4 clk_r_REG425_S1 ( .D(n12764), .E(\u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n17680) );
  HS65_LL_DFPHQX4 clk_r_REG406_S1 ( .D(n12851), .E(\u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n17677) );
  HS65_LL_DFPHQX4 clk_r_REG385_S1 ( .D(n12941), .E(\u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n17673) );
  HS65_LL_DFPHQX4 clk_r_REG345_S1 ( .D(n13121), .E(\u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n17665) );
  HS65_LL_DFPHQX4 clk_r_REG327_S1 ( .D(n13211), .E(\u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n17661) );
  HS65_LL_DFPHQX4 clk_r_REG224_S1 ( .D(n14104), .E(\u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n17635) );
  HS65_LL_DFPHQX4 clk_r_REG242_S1 ( .D(n14102), .E(\u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n17634) );
  HS65_LL_DFPHQX4 clk_r_REG201_S1 ( .D(n15458), .E(\u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n17482) );
  HS65_LH_DFPRQX4 clk_r_REG794_S3 ( .D(n12336), .CP(clk), .RN(n29651), .Q(
        n17705) );
  HS65_LH_DFPRQX4 clk_r_REG855_S3 ( .D(n12446), .CP(clk), .RN(n29648), .Q(
        n17696) );
  HS65_LH_DFPRQX4 clk_r_REG851_S3 ( .D(n12426), .CP(clk), .RN(n29652), .Q(
        n17698) );
  HS65_LH_DFPRQX4 clk_r_REG847_S3 ( .D(n13578), .CP(clk), .RN(n29648), .Q(
        n17648) );
  HS65_LH_DFPRQX4 clk_r_REG795_S3 ( .D(n12338), .CP(clk), .RN(n29647), .Q(
        n17704) );
  HS65_LH_DFPRQX4 clk_r_REG907_S3 ( .D(n11878), .CP(clk), .RN(n29647), .Q(
        n17728) );
  HS65_LH_DFPRQX4 clk_r_REG749_S3 ( .D(n12291), .CP(clk), .RN(n29697), .Q(
        n17709) );
  HS65_LH_DFPRQX4 clk_r_REG788_S3 ( .D(n12324), .CP(clk), .RN(n29650), .Q(
        n17707) );
  HS65_LH_DFPRQX4 clk_r_REG667_S3 ( .D(n9480), .CP(clk), .RN(n29647), .Q(
        n17847) );
  HS65_LH_DFPRQX4 clk_r_REG859_S3 ( .D(n12471), .CP(clk), .RN(n29697), .Q(
        n17694) );
  HS65_LH_DFPRQX4 clk_r_REG873_S3 ( .D(n15470), .CP(clk), .RN(n18160), .Q(
        n17577) );
  HS65_LH_DFPRQX4 clk_r_REG741_S3 ( .D(n11890), .CP(clk), .RN(n29644), .Q(
        n17726) );
  HS65_LH_DFPRQX4 clk_r_REG802_S3 ( .D(n12370), .CP(clk), .RN(n29644), .Q(
        n17702) );
  HS65_LH_DFPRQX4 clk_r_REG644_S3 ( .D(n13887), .CP(clk), .RN(n29698), .Q(
        n17641) );
  HS65_LH_DFPRQX4 clk_r_REG808_S3 ( .D(n12382), .CP(clk), .RN(n29651), .Q(
        n17701) );
  HS65_LH_DFPRQX4 clk_r_REG673_S3 ( .D(n13890), .CP(clk), .RN(n18160), .Q(
        n17640) );
  HS65_LH_DFPRQX4 clk_r_REG678_S3 ( .D(n11644), .CP(clk), .RN(n29697), .Q(
        n17740) );
  HS65_LH_DFPRQX4 clk_r_REG793_S3 ( .D(n12302), .CP(clk), .RN(n40997), .Q(
        n17708) );
  HS65_LH_DFPRQX4 clk_r_REG912_S3 ( .D(n11867), .CP(clk), .RN(n40998), .Q(
        n17729) );
  HS65_LH_DFPRQX4 clk_r_REG733_S3 ( .D(n11819), .CP(clk), .RN(n29650), .Q(
        n17731) );
  HS65_LH_DFPRQX4 clk_r_REG725_S3 ( .D(n11843), .CP(clk), .RN(n41000), .Q(
        n17730) );
  HS65_LH_DFPRQX4 clk_r_REG718_S3 ( .D(n11795), .CP(clk), .RN(n29643), .Q(
        n17732) );
  HS65_LH_DFPRQX4 clk_r_REG703_S3 ( .D(n11771), .CP(clk), .RN(n29652), .Q(
        n17733) );
  HS65_LH_DFPRQX4 clk_r_REG787_S3 ( .D(n12280), .CP(clk), .RN(n29644), .Q(
        n17710) );
  HS65_LH_DFPRQX4 clk_r_REG672_S3 ( .D(n2972), .CP(clk), .RN(n29698), .Q(
        n18082) );
  HS65_LH_DFPRQX4 clk_r_REG685_S3 ( .D(n11651), .CP(clk), .RN(n29698), .Q(
        n17738) );
  HS65_LH_DFPRQX4 clk_r_REG692_S3 ( .D(n11699), .CP(clk), .RN(n40997), .Q(
        n17736) );
  HS65_LH_DFPRQX4 clk_r_REG891_S3 ( .D(n13650), .CP(clk), .RN(n29698), .Q(
        n17643) );
  HS65_LH_DFPRQX4 clk_r_REG696_S3 ( .D(n11723), .CP(clk), .RN(n29652), .Q(
        n17735) );
  HS65_LH_DFPRQX4 clk_r_REG688_S3 ( .D(n11675), .CP(clk), .RN(n29646), .Q(
        n17737) );
  HS65_LH_DFPRQX4 clk_r_REG510_S2 ( .D(n12552), .CP(clk), .RN(n29698), .Q(
        n17688) );
  HS65_LH_DFPRQX4 clk_r_REG502_S2 ( .D(n12505), .CP(clk), .RN(n29650), .Q(
        n17690) );
  HS65_LH_DFPRQX4 clk_r_REG462_S2 ( .D(n12599), .CP(clk), .RN(n40998), .Q(
        n17686) );
  HS65_LH_DFPRQX4 clk_r_REG454_S2 ( .D(n9953), .CP(clk), .RN(n29697), .Q(
        n17822) );
  HS65_LH_DFPRQX4 clk_r_REG444_S2 ( .D(n12673), .CP(clk), .RN(n29643), .Q(
        n17684) );
  HS65_LH_DFPRQX4 clk_r_REG436_S2 ( .D(n12718), .CP(clk), .RN(n29645), .Q(
        n17683) );
  HS65_LH_DFPRQX4 clk_r_REG428_S2 ( .D(n12763), .CP(clk), .RN(n29643), .Q(
        n17681) );
  HS65_LH_DFPRQX4 clk_r_REG417_S2 ( .D(n12807), .CP(clk), .RN(n29648), .Q(
        n17679) );
  HS65_LH_DFPRQX4 clk_r_REG409_S2 ( .D(n12852), .CP(clk), .RN(n29651), .Q(
        n17676) );
  HS65_LH_DFPRQX4 clk_r_REG396_S2 ( .D(n12897), .CP(clk), .RN(n29646), .Q(
        n17675) );
  HS65_LH_DFPRQX4 clk_r_REG388_S2 ( .D(n12942), .CP(clk), .RN(n29645), .Q(
        n17672) );
  HS65_LH_DFPRQX4 clk_r_REG378_S2 ( .D(n12987), .CP(clk), .RN(n29643), .Q(
        n17671) );
  HS65_LH_DFPRQX4 clk_r_REG371_S2 ( .D(n13032), .CP(clk), .RN(n29652), .Q(
        n17668) );
  HS65_LH_DFPRQX4 clk_r_REG361_S2 ( .D(n13077), .CP(clk), .RN(n29650), .Q(
        n17667) );
  HS65_LH_DFPRQX4 clk_r_REG348_S2 ( .D(n13122), .CP(clk), .RN(n29646), .Q(
        n17664) );
  HS65_LH_DFPRQX4 clk_r_REG338_S2 ( .D(n13167), .CP(clk), .RN(n29644), .Q(
        n17663) );
  HS65_LH_DFPRQX4 clk_r_REG330_S2 ( .D(n13212), .CP(clk), .RN(n29648), .Q(
        n17660) );
  HS65_LH_DFPRQX4 clk_r_REG319_S2 ( .D(n13257), .CP(clk), .RN(n29647), .Q(
        n17659) );
  HS65_LH_DFPRQX4 clk_r_REG311_S2 ( .D(n13302), .CP(clk), .RN(n29647), .Q(
        n17657) );
  HS65_LH_DFPRQX4 clk_r_REG303_S2 ( .D(n11921), .CP(clk), .RN(n29643), .Q(
        n17723) );
  HS65_LH_DFPRQX4 clk_r_REG295_S2 ( .D(n11966), .CP(clk), .RN(n29697), .Q(
        n17721) );
  HS65_LH_DFPRQX4 clk_r_REG287_S2 ( .D(n12011), .CP(clk), .RN(n29698), .Q(
        n17719) );
  HS65_LH_DFPRQX4 clk_r_REG279_S2 ( .D(n12056), .CP(clk), .RN(n29644), .Q(
        n17717) );
  HS65_LH_DFPRQX4 clk_r_REG271_S2 ( .D(n12101), .CP(clk), .RN(n29698), .Q(
        n17715) );
  HS65_LH_DFPRQX4 clk_r_REG263_S2 ( .D(n12146), .CP(clk), .RN(n29646), .Q(
        n17713) );
  HS65_LH_DFPRQX4 clk_r_REG253_S2 ( .D(n12191), .CP(clk), .RN(n29650), .Q(
        n17712) );
  HS65_LH_DFPRQX4 clk_r_REG245_S2 ( .D(n12236), .CP(clk), .RN(n29697), .Q(
        n17711) );
  HS65_LH_DFPRQX4 clk_r_REG235_S2 ( .D(n13347), .CP(clk), .RN(n17245), .Q(
        n17655) );
  HS65_LH_DFPRQX4 clk_r_REG227_S2 ( .D(n13392), .CP(clk), .RN(n29649), .Q(
        n17654) );
  HS65_LH_DFPRQX4 clk_r_REG217_S2 ( .D(n13437), .CP(clk), .RN(n29645), .Q(
        n17653) );
  HS65_LH_DFPRQX4 clk_r_REG212_S2 ( .D(n13540), .CP(clk), .RN(n18160), .Q(
        n17649) );
  HS65_LH_DFPRQX4 clk_r_REG203_S2 ( .D(n13482), .CP(clk), .RN(n29652), .Q(
        n17652) );
  HS65_LH_DFPRQX4 clk_r_REG699_S3 ( .D(n11747), .CP(clk), .RN(n29651), .Q(
        n17734) );
  HS65_LH_DFPRQX4 clk_r_REG742_S3 ( .D(n11889), .CP(clk), .RN(n29652), .Q(
        n17727) );
  HS65_LH_DFPRQX4 clk_r_REG858_S3 ( .D(n12436), .CP(clk), .RN(n29649), .Q(
        n17697) );
  HS65_LH_DFPRQX4 clk_r_REG854_S3 ( .D(n12414), .CP(clk), .RN(n17245), .Q(
        n17699) );
  HS65_LH_DFPRQX4 clk_r_REG864_S3 ( .D(n12458), .CP(clk), .RN(n29646), .Q(
        n17695) );
  HS65_LH_DFPRQX4 clk_r_REG850_S3 ( .D(n12393), .CP(clk), .RN(n29650), .Q(
        n17700) );
  HS65_LH_DFPRQX4 clk_r_REG903_S3 ( .D(n12480), .CP(clk), .RN(n29645), .Q(
        n17693) );
  HS65_LH_DFPRQX4 clk_r_REG801_S3 ( .D(n12325), .CP(clk), .RN(n29645), .Q(
        n17706) );
  HS65_LH_DFPRQX4 clk_r_REG807_S3 ( .D(n12347), .CP(clk), .RN(n29648), .Q(
        n17703) );
  HS65_LH_DFPRQX4 clk_r_REG666_S3 ( .D(n11913), .CP(clk), .RN(n29697), .Q(
        n17725) );
  HS65_LH_DFPRQX4 clk_r_REG684_S3 ( .D(n11645), .CP(clk), .RN(n29697), .Q(
        n17739) );
  HS65_LH_DFPRQX4 clk_r_REG662_S3 ( .D(n11916), .CP(clk), .RN(n29649), .Q(
        n17724) );
  HS65_LH_DFPRQX4 clk_r_REG677_S3 ( .D(n2973), .CP(clk), .RN(n29645), .Q(
        n18081) );
  HS65_LH_DFPRQX4 clk_r_REG9_S1 ( .D(n12490), .CP(clk), .RN(n29650), .Q(n17692) );
  HS65_LH_DFPRQX4 clk_r_REG511_S2 ( .D(n9950), .CP(clk), .RN(n29651), .Q(
        n17825) );
  HS65_LH_DFPRQX4 clk_r_REG503_S2 ( .D(n9949), .CP(clk), .RN(n29650), .Q(
        n17826) );
  HS65_LH_DFPRQX4 clk_r_REG463_S2 ( .D(n9951), .CP(clk), .RN(n29649), .Q(
        n17824) );
  HS65_LH_DFPRQX4 clk_r_REG455_S2 ( .D(n9952), .CP(clk), .RN(n29698), .Q(
        n17823) );
  HS65_LH_DFPRQX4 clk_r_REG445_S2 ( .D(n9962), .CP(clk), .RN(n18160), .Q(
        n17821) );
  HS65_LH_DFPRQX4 clk_r_REG437_S2 ( .D(n9963), .CP(clk), .RN(n41000), .Q(
        n17820) );
  HS65_LH_DFPRQX4 clk_r_REG429_S2 ( .D(n9964), .CP(clk), .RN(n29647), .Q(
        n17819) );
  HS65_LH_DFPRQX4 clk_r_REG418_S2 ( .D(n9965), .CP(clk), .RN(n29649), .Q(
        n17818) );
  HS65_LH_DFPRQX4 clk_r_REG410_S2 ( .D(n9966), .CP(clk), .RN(n17245), .Q(
        n17817) );
  HS65_LH_DFPRQX4 clk_r_REG397_S2 ( .D(n9967), .CP(clk), .RN(n29649), .Q(
        n17816) );
  HS65_LH_DFPRQX4 clk_r_REG389_S2 ( .D(n9968), .CP(clk), .RN(n29646), .Q(
        n17815) );
  HS65_LH_DFPRQX4 clk_r_REG379_S2 ( .D(n9969), .CP(clk), .RN(n29698), .Q(
        n17814) );
  HS65_LH_DFPRQX4 clk_r_REG372_S2 ( .D(n9970), .CP(clk), .RN(n29646), .Q(
        n17813) );
  HS65_LH_DFPRQX4 clk_r_REG362_S2 ( .D(n9971), .CP(clk), .RN(n29652), .Q(
        n17812) );
  HS65_LH_DFPRQX4 clk_r_REG349_S2 ( .D(n9972), .CP(clk), .RN(n29652), .Q(
        n17811) );
  HS65_LH_DFPRQX4 clk_r_REG339_S2 ( .D(n9973), .CP(clk), .RN(n29650), .Q(
        n17810) );
  HS65_LH_DFPRQX4 clk_r_REG331_S2 ( .D(n9974), .CP(clk), .RN(n40997), .Q(
        n17809) );
  HS65_LH_DFPRQX4 clk_r_REG320_S2 ( .D(n9975), .CP(clk), .RN(n29697), .Q(
        n17808) );
  HS65_LH_DFPRQX4 clk_r_REG312_S2 ( .D(n9976), .CP(clk), .RN(n40998), .Q(
        n17807) );
  HS65_LH_DFPRQX4 clk_r_REG304_S2 ( .D(n9977), .CP(clk), .RN(n17245), .Q(
        n17806) );
  HS65_LH_DFPRQX4 clk_r_REG296_S2 ( .D(n9978), .CP(clk), .RN(n29644), .Q(
        n17805) );
  HS65_LH_DFPRQX4 clk_r_REG288_S2 ( .D(n9979), .CP(clk), .RN(n29697), .Q(
        n17804) );
  HS65_LH_DFPRQX4 clk_r_REG280_S2 ( .D(n9980), .CP(clk), .RN(n29646), .Q(
        n17803) );
  HS65_LH_DFPRQX4 clk_r_REG272_S2 ( .D(n9981), .CP(clk), .RN(n29650), .Q(
        n17802) );
  HS65_LH_DFPRQX4 clk_r_REG264_S2 ( .D(n9982), .CP(clk), .RN(n29652), .Q(
        n17801) );
  HS65_LH_DFPRQX4 clk_r_REG254_S2 ( .D(n9983), .CP(clk), .RN(n29647), .Q(
        n17800) );
  HS65_LH_DFPRQX4 clk_r_REG246_S2 ( .D(n9984), .CP(clk), .RN(n18160), .Q(
        n17799) );
  HS65_LH_DFPRQX4 clk_r_REG236_S2 ( .D(n9985), .CP(clk), .RN(n29646), .Q(
        n17798) );
  HS65_LH_DFPRQX4 clk_r_REG228_S2 ( .D(n9986), .CP(clk), .RN(n29651), .Q(
        n17797) );
  HS65_LH_DFPRQX4 clk_r_REG218_S2 ( .D(n9987), .CP(clk), .RN(n29651), .Q(
        n17796) );
  HS65_LH_DFPRQX4 clk_r_REG213_S2 ( .D(n9989), .CP(clk), .RN(n17245), .Q(
        n17794) );
  HS65_LH_DFPRQX4 clk_r_REG204_S2 ( .D(n9988), .CP(clk), .RN(n29644), .Q(
        n17795) );
  HS65_LH_DFPRQX4 clk_r_REG904_S3 ( .D(n10102), .CP(clk), .RN(n29645), .Q(
        n17788) );
  HS65_LH_DFPRQX4 clk_r_REG871_S3 ( .D(n278), .CP(clk), .RN(n29647), .Q(n17446) );
  HS65_LH_DFPRQX4 clk_r_REG689_S3 ( .D(n9477), .CP(clk), .RN(n29643), .Q(
        n17848) );
  HS65_LH_DFPRQX4 clk_r_REG867_S3 ( .D(n15748), .CP(clk), .RN(n29650), .Q(
        n17514) );
  HS65_LH_DFPRQX4 clk_r_REG669_S3 ( .D(n242), .CP(clk), .RN(n29645), .Q(n17438) );
  HS65_LH_DFPRQX4 clk_r_REG679_S3 ( .D(n196), .CP(clk), .RN(n29648), .Q(n17511) );
  HS65_LH_DFPRQX4 clk_r_REG893_S3 ( .D(n15475), .CP(clk), .RN(n29651), .Q(
        n17630) );
  HS65_LH_DFPRQX4 clk_r_REG874_S3 ( .D(n17204), .CP(clk), .RN(n18160), .Q(
        n17444) );
  HS65_LH_DFPRQX4 clk_r_REG621_S1 ( .D(n192), .CP(clk), .RN(n40998), .Q(n17436) );
  HS65_LH_DFPRQX4 clk_r_REG894_S3 ( .D(n178), .CP(clk), .RN(n29651), .Q(n17316) );
  HS65_LH_DFPRQX4 clk_r_REG759_S3 ( .D(n16464), .CP(clk), .RN(n29646), .Q(
        n17409) );
  HS65_LH_DFPRQX4 clk_r_REG751_S3 ( .D(n16417), .CP(clk), .RN(n29644), .Q(
        n17410) );
  HS65_LH_DFPRQX4 clk_r_REG837_S3 ( .D(n17184), .CP(clk), .RN(n18160), .Q(
        n17383) );
  HS65_LH_DFPRQX4 clk_r_REG830_S3 ( .D(n17101), .CP(clk), .RN(n41000), .Q(
        n17382) );
  HS65_LH_DFPRQX4 clk_r_REG818_S3 ( .D(n17133), .CP(clk), .RN(n29646), .Q(
        n17380) );
  HS65_LH_DFPRQX4 clk_r_REG647_S3 ( .D(n274), .CP(clk), .RN(n29650), .Q(n17512) );
  HS65_LH_DFPRQX4 clk_r_REG844_S3 ( .D(n17182), .CP(clk), .RN(n29646), .Q(
        n17516) );
  HS65_LH_DFPRQX4 clk_r_REG826_S3 ( .D(n17131), .CP(clk), .RN(n29645), .Q(
        n17517) );
  HS65_LH_DFPRQX4 clk_r_REG612_S1 ( .D(n282), .CP(clk), .RN(n29646), .Q(n17445) );
  HS65_LH_DFPRQX4 clk_r_REG832_S3 ( .D(n17092), .CP(clk), .RN(n29644), .Q(
        n17391) );
  HS65_LH_DFPRQX4 clk_r_REG809_S3 ( .D(n17171), .CP(clk), .RN(n29648), .Q(
        n17385) );
  HS65_LH_DFPRQX4 clk_r_REG840_S3 ( .D(n17083), .CP(clk), .RN(n29645), .Q(
        n17393) );
  HS65_LH_DFPRQX4 clk_r_REG758_S3 ( .D(n16412), .CP(clk), .RN(n29649), .Q(
        n17407) );
  HS65_LH_DFPRQX4 clk_r_REG752_S3 ( .D(n16461), .CP(clk), .RN(n17245), .Q(
        n17414) );
  HS65_LH_DFPRQX4 clk_r_REG876_S3 ( .D(n209), .CP(clk), .RN(n29652), .Q(n17569) );
  HS65_LH_DFPRQX4 clk_r_REG841_S3 ( .D(n17146), .CP(clk), .RN(n29652), .Q(
        n17394) );
  HS65_LH_DFPRQX4 clk_r_REG834_S3 ( .D(n17158), .CP(clk), .RN(n29651), .Q(
        n17399) );
  HS65_LH_DFPRQX4 clk_r_REG833_S3 ( .D(n17111), .CP(clk), .RN(n29650), .Q(
        n17392) );
  HS65_LH_DFPRQX4 clk_r_REG839_S3 ( .D(n17048), .CP(clk), .RN(n40997), .Q(
        n17388) );
  HS65_LH_DFPRQX4 clk_r_REG836_S3 ( .D(n17172), .CP(clk), .RN(n29651), .Q(
        n17379) );
  HS65_LH_DFPRQX4 clk_r_REG819_S3 ( .D(n17173), .CP(clk), .RN(n29698), .Q(
        n17384) );
  HS65_LH_DFPRQX4 clk_r_REG813_S3 ( .D(n17178), .CP(clk), .RN(n29645), .Q(
        n17389) );
  HS65_LH_DFPRQX4 clk_r_REG823_S3 ( .D(n17110), .CP(clk), .RN(n29652), .Q(
        n17396) );
  HS65_LH_DFPRQX4 clk_r_REG760_S3 ( .D(n16387), .CP(clk), .RN(n29651), .Q(
        n17412) );
  HS65_LH_DFPRQX4 clk_r_REG838_S3 ( .D(n17174), .CP(clk), .RN(n29643), .Q(
        n17387) );
  HS65_LH_DFPRQX4 clk_r_REG829_S3 ( .D(n17134), .CP(clk), .RN(n18160), .Q(
        n17381) );
  HS65_LH_DFPRQX4 clk_r_REG817_S3 ( .D(n17139), .CP(clk), .RN(n29648), .Q(
        n17378) );
  HS65_LH_DFPRQX4 clk_r_REG810_S3 ( .D(n17045), .CP(clk), .RN(n29698), .Q(
        n17390) );
  HS65_LH_DFPRQX4 clk_r_REG835_S3 ( .D(n17114), .CP(clk), .RN(n29647), .Q(
        n17401) );
  HS65_LH_DFPRQX4 clk_r_REG825_S3 ( .D(n17090), .CP(clk), .RN(n29643), .Q(
        n17402) );
  HS65_LH_DFPRQX4 clk_r_REG842_S3 ( .D(n17066), .CP(clk), .RN(n29647), .Q(
        n17403) );
  HS65_LH_DFPRQX4 clk_r_REG824_S3 ( .D(n17147), .CP(clk), .RN(n29645), .Q(
        n17400) );
  HS65_LH_DFPRQX4 clk_r_REG761_S3 ( .D(n16456), .CP(clk), .RN(n29643), .Q(
        n17415) );
  HS65_LH_DFPRQX4 clk_r_REG750_S3 ( .D(n16466), .CP(clk), .RN(n29645), .Q(
        n17408) );
  HS65_LH_DFPRQX4 clk_r_REG768_S3 ( .D(n16352), .CP(clk), .RN(n29648), .Q(
        n17411) );
  HS65_LH_DFPRQX4 clk_r_REG769_S3 ( .D(n16455), .CP(clk), .RN(n29645), .Q(
        n17416) );
  HS65_LH_DFPRQX4 clk_r_REG767_S3 ( .D(n16457), .CP(clk), .RN(n40998), .Q(
        n17406) );
  HS65_LH_DFPRQX4 clk_r_REG762_S3 ( .D(n16429), .CP(clk), .RN(n29649), .Q(
        n17421) );
  HS65_LH_DFPRQX4 clk_r_REG845_S3 ( .D(n17097), .CP(clk), .RN(n29643), .Q(
        n17564) );
  HS65_LH_DFPRQX4 clk_r_REG827_S3 ( .D(n17183), .CP(clk), .RN(n29652), .Q(
        n17562) );
  HS65_LH_DFPRQX4 clk_r_REG812_S3 ( .D(n17156), .CP(clk), .RN(n18160), .Q(
        n17398) );
  HS65_LH_DFPRQX4 clk_r_REG629_S1 ( .D(n179), .CP(clk), .RN(n29651), .Q(n17373) );
  HS65_LH_DFPRQX4 clk_r_REG811_S3 ( .D(n17060), .CP(clk), .RN(n40997), .Q(
        n17397) );
  HS65_LH_DFPRQX4 clk_r_REG831_S3 ( .D(n17132), .CP(clk), .RN(n29646), .Q(
        n17386) );
  HS65_LH_DFPRQX4 clk_r_REG814_S3 ( .D(n17127), .CP(clk), .RN(n29649), .Q(
        n17377) );
  HS65_LH_DFPRQX4 clk_r_REG12_S1 ( .D(n17207), .CP(clk), .RN(n29645), .Q(
        n17573) );
  HS65_LH_DFPRQX4 clk_r_REG772_S3 ( .D(n16317), .CP(clk), .RN(n29651), .Q(
        n17428) );
  HS65_LH_DFPRQX4 clk_r_REG764_S3 ( .D(n16436), .CP(clk), .RN(n29644), .Q(
        n17425) );
  HS65_LH_DFPRQX4 clk_r_REG753_S3 ( .D(n16405), .CP(clk), .RN(n29698), .Q(
        n17423) );
  HS65_LH_DFPRQX4 clk_r_REG770_S3 ( .D(n16439), .CP(clk), .RN(n41000), .Q(
        n17419) );
  HS65_LH_DFPRQX4 clk_r_REG778_S3 ( .D(n16411), .CP(clk), .RN(n29652), .Q(
        n17418) );
  HS65_LH_DFPRQX4 clk_r_REG776_S3 ( .D(n16351), .CP(clk), .RN(n29649), .Q(
        n17413) );
  HS65_LH_DFPRQX4 clk_r_REG781_S3 ( .D(n16393), .CP(clk), .RN(n29651), .Q(
        n17429) );
  HS65_LH_DFPRQX4 clk_r_REG775_S3 ( .D(n16473), .CP(clk), .RN(n18160), .Q(
        n17405) );
  HS65_LH_DFPRQX4 clk_r_REG782_S3 ( .D(n16367), .CP(clk), .RN(n29646), .Q(
        n17431) );
  HS65_LH_DFPRQX4 clk_r_REG777_S3 ( .D(n16377), .CP(clk), .RN(n29652), .Q(
        n17417) );
  HS65_LH_DFPRQX4 clk_r_REG780_S3 ( .D(n16392), .CP(clk), .RN(n29698), .Q(
        n17422) );
  HS65_LH_DFPRQX4 clk_r_REG771_S3 ( .D(n16394), .CP(clk), .RN(n40997), .Q(
        n17426) );
  HS65_LH_DFPRQX4 clk_r_REG763_S3 ( .D(n16400), .CP(clk), .RN(n40998), .Q(
        n17424) );
  HS65_LH_DFPRQX4 clk_r_REG755_S3 ( .D(n16395), .CP(clk), .RN(n29698), .Q(
        n17432) );
  HS65_LH_DFPRQX4 clk_r_REG765_S3 ( .D(n16368), .CP(clk), .RN(n29698), .Q(
        n17430) );
  HS65_LH_DFPRQX4 clk_r_REG754_S3 ( .D(n16437), .CP(clk), .RN(n29649), .Q(
        n17427) );
  HS65_LH_DFPRQX4 clk_r_REG614_S1 ( .D(n17205), .CP(clk), .RN(n29649), .Q(
        n17305) );
  HS65_LH_DFPRQX4 clk_r_REG820_S3 ( .D(n16483), .CP(clk), .RN(n29652), .Q(
        n17395) );
  HS65_LH_DFPRQX4 clk_r_REG816_S3 ( .D(n13904), .CP(clk), .RN(n29651), .Q(
        n18121) );
  HS65_LH_DFPRQX4 clk_r_REG757_S3 ( .D(n13898), .CP(clk), .RN(n29647), .Q(
        n18126) );
  HS65_LH_DFPRQX4 clk_r_REG815_S3 ( .D(n13944), .CP(clk), .RN(n29644), .Q(
        n18124) );
  HS65_LH_DFPRQX4 clk_r_REG774_S3 ( .D(n13896), .CP(clk), .RN(n29645), .Q(
        n18123) );
  HS65_LH_DFPRQX4 clk_r_REG773_S3 ( .D(n13902), .CP(clk), .RN(n29646), .Q(
        n18125) );
  HS65_LH_DFPRQX4 clk_r_REG756_S3 ( .D(n13900), .CP(clk), .RN(n29649), .Q(
        n18122) );
  HS65_LH_DFPRQX4 clk_r_REG822_S3 ( .D(n17035), .CP(clk), .RN(n29648), .Q(
        n17565) );
  HS65_LH_DFPRQX4 clk_r_REG821_S3 ( .D(n17122), .CP(clk), .RN(n17245), .Q(
        n17563) );
  HS65_LH_DFPRQX4 clk_r_REG603_S1 ( .D(n280), .CP(clk), .RN(n17245), .Q(n17440) );
  HS65_LH_DFPRQX4 clk_r_REG645_S3 ( .D(n198), .CP(clk), .RN(n29649), .Q(n17300) );
  HS65_LH_DFPRQX4 clk_r_REG599_S1 ( .D(n15759), .CP(clk), .RN(n29649), .Q(
        n17296) );
  HS65_LH_DFPRQX4 clk_r_REG653_S3 ( .D(n225), .CP(clk), .RN(n29648), .Q(n17435) );
  HS65_LH_DFPRQX4 clk_r_REG601_S1 ( .D(n15761), .CP(clk), .RN(n18160), .Q(
        n17434) );
  HS65_LH_DFPRQX4 clk_r_REG613_S1 ( .D(n15760), .CP(clk), .RN(n29649), .Q(
        n17566) );
  HS65_LH_DFPRQX4 clk_r_REG610_S1 ( .D(n15708), .CP(clk), .RN(n29698), .Q(
        n17267) );
  HS65_LL_DFPHQX27 clk_r_REG197_S1 ( .D(addr_to_iram_0), .E(
        \u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n17639) );
  HS65_LH_DFPQX4 clk_r_REG574_S2 ( .D(\u_DataPath/u_idexreg/N184 ), .CP(clk), 
        .Q(n17527) );
  HS65_LH_DFPQX4 clk_r_REG575_S2 ( .D(n5958), .CP(clk), .Q(n17991) );
  HS65_LH_DFPQX4 clk_r_REG639_S1 ( .D(n13591), .CP(clk), .Q(n17647) );
  HS65_LH_DFPQX4 clk_r_REG609_S3 ( .D(n1065), .CP(clk), .Q(n17326) );
  HS65_LH_DFPQX4 clk_r_REG529_S11 ( .D(\u_DataPath/data_read_ex_2_i [31]), 
        .CP(clk), .Q(n17342) );
  HS65_LH_DFPQX4 clk_r_REG544_S2 ( .D(\u_DataPath/data_read_ex_2_i [18]), .CP(
        clk), .Q(n17343) );
  HS65_LH_DFPQX4 clk_r_REG543_S2 ( .D(\u_DataPath/data_read_ex_2_i [25]), .CP(
        clk), .Q(n17329) );
  HS65_LH_DFPQX4 clk_r_REG494_S2 ( .D(\u_DataPath/data_read_ex_2_i [10]), .CP(
        clk), .Q(n17351) );
  HS65_LH_DFPQX4 clk_r_REG492_S2 ( .D(\u_DataPath/data_read_ex_2_i [8]), .CP(
        clk), .Q(n17350) );
  HS65_LH_DFPQX4 clk_r_REG490_S2 ( .D(\u_DataPath/data_read_ex_2_i [7]), .CP(
        clk), .Q(n17348) );
  HS65_LH_DFPQX4 clk_r_REG482_S2 ( .D(\u_DataPath/data_read_ex_2_i [13]), .CP(
        clk), .Q(n17355) );
  HS65_LH_DFPQX4 clk_r_REG476_S2 ( .D(\u_DataPath/data_read_ex_2_i [11]), .CP(
        clk), .Q(n17349) );
  HS65_LH_DFPQX4 clk_r_REG474_S2 ( .D(\u_DataPath/data_read_ex_2_i [12]), .CP(
        clk), .Q(n17352) );
  HS65_LH_DFPQX4 clk_r_REG472_S2 ( .D(\u_DataPath/data_read_ex_2_i [22]), .CP(
        clk), .Q(n17344) );
  HS65_LH_DFPQX4 clk_r_REG471_S2 ( .D(\u_DataPath/data_read_ex_2_i [15]), .CP(
        clk), .Q(n17353) );
  HS65_LH_DFPQX4 clk_r_REG595_S2 ( .D(\u_DataPath/data_read_ex_2_i [20]), .CP(
        clk), .Q(n17334) );
  HS65_LH_DFPQX4 clk_r_REG545_S2 ( .D(\u_DataPath/data_read_ex_2_i [17]), .CP(
        clk), .Q(n17335) );
  HS65_LH_DFPQX4 clk_r_REG542_S2 ( .D(\u_DataPath/data_read_ex_2_i [26]), .CP(
        clk), .Q(n17332) );
  HS65_LH_DFPQX4 clk_r_REG541_S2 ( .D(\u_DataPath/data_read_ex_2_i [30]), .CP(
        clk), .Q(n17341) );
  HS65_LH_DFPQX4 clk_r_REG497_S2 ( .D(\u_DataPath/data_read_ex_2_i [5]), .CP(
        clk), .Q(n17345) );
  HS65_LH_DFPQX4 clk_r_REG496_S2 ( .D(\u_DataPath/data_read_ex_2_i [9]), .CP(
        clk), .Q(n17346) );
  HS65_LH_DFPQX4 clk_r_REG491_S2 ( .D(\u_DataPath/data_read_ex_2_i [23]), .CP(
        clk), .Q(n17333) );
  HS65_LH_DFPQX4 clk_r_REG487_S2 ( .D(\u_DataPath/data_read_ex_2_i [28]), .CP(
        clk), .Q(n17336) );
  HS65_LH_DFPQX4 clk_r_REG486_S2 ( .D(\u_DataPath/data_read_ex_2_i [21]), .CP(
        clk), .Q(n17337) );
  HS65_LH_DFPQX4 clk_r_REG485_S2 ( .D(\u_DataPath/data_read_ex_2_i [24]), .CP(
        clk), .Q(n17340) );
  HS65_LH_DFPQX4 clk_r_REG484_S2 ( .D(\u_DataPath/data_read_ex_2_i [29]), .CP(
        clk), .Q(n17331) );
  HS65_LH_DFPQX4 clk_r_REG483_S2 ( .D(\u_DataPath/data_read_ex_2_i [19]), .CP(
        clk), .Q(n17339) );
  HS65_LH_DFPQX4 clk_r_REG480_S2 ( .D(\u_DataPath/data_read_ex_2_i [16]), .CP(
        clk), .Q(n17330) );
  HS65_LH_DFPQX4 clk_r_REG478_S2 ( .D(\u_DataPath/data_read_ex_2_i [6]), .CP(
        clk), .Q(n17347) );
  HS65_LH_DFPQX4 clk_r_REG469_S2 ( .D(\u_DataPath/data_read_ex_2_i [27]), .CP(
        clk), .Q(n17338) );
  HS65_LH_DFPQX4 clk_r_REG468_S2 ( .D(\u_DataPath/data_read_ex_2_i [2]), .CP(
        clk), .Q(n17354) );
  HS65_LH_DFPQX4 clk_r_REG597_S2 ( .D(n15212), .CP(clk), .Q(n17608) );
  HS65_LH_DFPQX4 clk_r_REG37_S5 ( .D(n35544), .CP(clk), .Q(n17280) );
  HS65_LH_DFPQX4 clk_r_REG571_S2 ( .D(\u_DataPath/cw_to_ex_i [0]), .CP(clk), 
        .Q(n17246) );
  HS65_LH_DFPQX4 clk_r_REG41_S6 ( .D(n35195), .CP(clk), .Q(n17272) );
  HS65_LH_DFPQX4 clk_r_REG266_S4 ( .D(n1029), .CP(clk), .Q(n17284) );
  HS65_LH_DFPQX4 clk_r_REG257_S4 ( .D(n1027), .CP(clk), .Q(n17285) );
  HS65_LH_DFPQX4 clk_r_REG206_S4 ( .D(n1020), .CP(clk), .Q(n17286) );
  HS65_LH_DFPQX4 clk_r_REG568_S2 ( .D(\u_DataPath/cw_to_ex_i [1]), .CP(clk), 
        .Q(n17283) );
  HS65_LH_DFPQX4 clk_r_REG640_S1 ( .D(n11622), .CP(clk), .Q(n17741) );
  HS65_LH_DFPQX4 clk_r_REG572_S2 ( .D(n14225), .CP(clk), .Q(n17607) );
  HS65_LH_DFPQX4 clk_r_REG13_S2 ( .D(\u_DataPath/cw_to_ex_i [4]), .CP(clk), 
        .Q(n17266) );
  HS65_LH_DFPQX4 clk_r_REG611_S2 ( .D(\u_DataPath/cw_to_ex_i [3]), .CP(clk), 
        .Q(n17328) );
  HS65_LH_DFPQX4 clk_r_REG573_S2 ( .D(n14244), .CP(clk), .Q(n17606) );
  HS65_LH_DFPQX4 clk_r_REG636_S1 ( .D(n10721), .CP(clk), .Q(n17760) );
  HS65_LH_DFPQX4 clk_r_REG499_S11 ( .D(n9234), .CP(clk), .Q(n17862) );
  HS65_LH_DFPQX4 clk_r_REG800_S1 ( .D(n15488), .CP(clk), .Q(n17620) );
  HS65_LH_DFPQX4 clk_r_REG642_S1 ( .D(n13613), .CP(clk), .Q(n17646) );
  HS65_LH_DFPQX4 clk_r_REG898_S5 ( .D(n10158), .CP(clk), .Q(n17782) );
  HS65_LH_DFPQX4 clk_r_REG600_S2 ( .D(n15319), .CP(clk), .Q(n17605) );
  HS65_LH_DFPQX4 clk_r_REG899_S5 ( .D(n15477), .CP(clk), .Q(n17629) );
  HS65_LH_DFPQX4 clk_r_REG791_S1 ( .D(n15485), .CP(clk), .Q(n17623) );
  HS65_LH_DFPQX4 clk_r_REG631_S3 ( .D(n9290), .CP(clk), .Q(n17855) );
  HS65_LH_DFPQX4 clk_r_REG628_S3 ( .D(n9289), .CP(clk), .Q(n17856) );
  HS65_LH_DFPQX4 clk_r_REG900_S5 ( .D(n10228), .CP(clk), .Q(n17781) );
  HS65_LH_DFPQX4 clk_r_REG569_S2 ( .D(n15374), .CP(clk), .Q(n17473) );
  HS65_LH_DFPQX4 clk_r_REG546_S2 ( .D(n15385), .CP(clk), .Q(n17472) );
  HS65_LH_DFPQX4 clk_r_REG556_S2 ( .D(n15709), .CP(clk), .Q(n17469) );
  HS65_LH_DFPQX4 clk_r_REG524_S10 ( .D(n15210), .CP(clk), .Q(n17311) );
  HS65_LH_DFPQX4 clk_r_REG570_S2 ( .D(n15380), .CP(clk), .Q(n17475) );
  HS65_LH_DFPQX4 clk_r_REG523_S11 ( .D(n9112), .CP(clk), .Q(n17867) );
  HS65_LH_DFPQX4 clk_r_REG549_S2 ( .D(n15501), .CP(clk), .Q(n17314) );
  HS65_LH_DFPQX4 clk_r_REG879_S5 ( .D(n10678), .CP(clk), .Q(n17762) );
  HS65_LH_DFPQX4 clk_r_REG561_S2 ( .D(n15149), .CP(clk), .Q(n17468) );
  HS65_LH_DFPQX4 clk_r_REG557_S2 ( .D(n15720), .CP(clk), .Q(n17467) );
  HS65_LH_DFPQX4 clk_r_REG604_S2 ( .D(n10755), .CP(clk), .Q(n17755) );
  HS65_LH_DFPQX4 clk_r_REG508_S4 ( .D(n2821), .CP(clk), .Q(n18090) );
  HS65_LH_DFPQX4 clk_r_REG506_S4 ( .D(n2774), .CP(clk), .Q(n18091) );
  HS65_LH_DFPQX4 clk_r_REG514_S3 ( .D(n10754), .CP(clk), .Q(n17756) );
  HS65_LH_DFPQX4 clk_r_REG466_S3 ( .D(n8838), .CP(clk), .Q(n17876) );
  HS65_LH_DFPQX4 clk_r_REG552_S2 ( .D(n15411), .CP(clk), .Q(n17523) );
  HS65_LH_DFPQX4 clk_r_REG504_S3 ( .D(n9374), .CP(clk), .Q(n17850) );
  HS65_LH_DFPQX4 clk_r_REG547_S2 ( .D(n15151), .CP(clk), .Q(n17315) );
  HS65_LH_DFPQX4 clk_r_REG550_S2 ( .D(n15408), .CP(clk), .Q(n17471) );
  HS65_LH_DFPQX4 clk_r_REG799_S1 ( .D(n9822), .CP(clk), .Q(n17831) );
  HS65_LH_DFPQX4 clk_r_REG553_S2 ( .D(n15342), .CP(clk), .Q(n17587) );
  HS65_LH_DFPQX4 clk_r_REG532_S1 ( .D(n9319), .CP(clk), .Q(n17851) );
  HS65_LH_DFPQX4 clk_r_REG14_S2 ( .D(n15407), .CP(clk), .Q(n17310) );
  HS65_LH_DFPQX4 clk_r_REG605_S2 ( .D(n8837), .CP(clk), .Q(n17877) );
  HS65_LH_DFPQX4 clk_r_REG660_S1 ( .D(n8558), .CP(clk), .Q(n17887) );
  HS65_LH_DFPQX4 clk_r_REG548_S2 ( .D(n15522), .CP(clk), .Q(n17638) );
  HS65_LH_DFPQX4 clk_r_REG618_S2 ( .D(n10382), .CP(clk), .Q(n17770) );
  HS65_LH_DFPQX4 clk_r_REG551_S2 ( .D(n14821), .CP(clk), .Q(n17604) );
  HS65_LH_DFPQX4 clk_r_REG786_S1 ( .D(n9668), .CP(clk), .Q(n17838) );
  HS65_LH_DFPQX4 clk_r_REG562_S2 ( .D(n15495), .CP(clk), .Q(n17603) );
  HS65_LH_DFPQX4 clk_r_REG558_S2 ( .D(n15393), .CP(clk), .Q(n17602) );
  HS65_LH_DFPQX4 clk_r_REG792_S1 ( .D(n9738), .CP(clk), .Q(n17835) );
  HS65_LH_DFPQX4 clk_r_REG633_S3 ( .D(n10040), .CP(clk), .Q(n17791) );
  HS65_LH_DFPQX4 clk_r_REG465_S4 ( .D(n10154), .CP(clk), .Q(n17784) );
  HS65_LH_DFPQX4 clk_r_REG457_S4 ( .D(n4211), .CP(clk), .Q(n18023) );
  HS65_LH_DFPQX4 clk_r_REG447_S2 ( .D(n2921), .CP(clk), .Q(n18084) );
  HS65_LH_DFPQX4 clk_r_REG439_S4 ( .D(n4323), .CP(clk), .Q(n18018) );
  HS65_LH_DFPQX4 clk_r_REG431_S4 ( .D(n2869), .CP(clk), .Q(n18088) );
  HS65_LH_DFPQX4 clk_r_REG420_S4 ( .D(n2975), .CP(clk), .Q(n18080) );
  HS65_LH_DFPQX4 clk_r_REG412_S4 ( .D(n3025), .CP(clk), .Q(n18078) );
  HS65_LH_DFPQX4 clk_r_REG400_S4 ( .D(n3078), .CP(clk), .Q(n18075) );
  HS65_LH_DFPQX4 clk_r_REG394_S4 ( .D(n3128), .CP(clk), .Q(n18073) );
  HS65_LH_DFPQX4 clk_r_REG384_S4 ( .D(n3181), .CP(clk), .Q(n18070) );
  HS65_LH_DFPQX4 clk_r_REG376_S4 ( .D(n3231), .CP(clk), .Q(n18068) );
  HS65_LH_DFPQX4 clk_r_REG367_S4 ( .D(n3284), .CP(clk), .Q(n18065) );
  HS65_LH_DFPQX4 clk_r_REG359_S4 ( .D(n3334), .CP(clk), .Q(n18063) );
  HS65_LH_DFPQX4 clk_r_REG344_S4 ( .D(n3387), .CP(clk), .Q(n18060) );
  HS65_LH_DFPQX4 clk_r_REG336_S4 ( .D(n3437), .CP(clk), .Q(n18058) );
  HS65_LH_DFPQX4 clk_r_REG326_S4 ( .D(n3490), .CP(clk), .Q(n18055) );
  HS65_LH_DFPQX4 clk_r_REG317_S4 ( .D(n3540), .CP(clk), .Q(n18053) );
  HS65_LH_DFPQX4 clk_r_REG42_S8 ( .D(n10750), .CP(clk), .Q(n17758) );
  HS65_LH_DFPQX4 clk_r_REG698_S4 ( .D(n7689), .CP(clk), .Q(n17925) );
  HS65_LH_DFPQX4 clk_r_REG695_S4 ( .D(n7882), .CP(clk), .Q(n17917) );
  HS65_LH_DFPQX4 clk_r_REG592_S3 ( .D(n9990), .CP(clk), .Q(n17793) );
  HS65_LH_DFPQX4 clk_r_REG882_S5 ( .D(n9483), .CP(clk), .Q(n17846) );
  HS65_LH_DFPQX4 clk_r_REG643_S1 ( .D(n10456), .CP(clk), .Q(n17769) );
  HS65_LH_DFPQX4 clk_r_REG701_S4 ( .D(n6789), .CP(clk), .Q(n17962) );
  HS65_LH_DFPQX4 clk_r_REG748_S4 ( .D(n9417), .CP(clk), .Q(n17849) );
  HS65_LH_DFPQX4 clk_r_REG806_S1 ( .D(n9869), .CP(clk), .Q(n17829) );
  HS65_LH_DFPQX4 clk_r_REG641_S1 ( .D(n10457), .CP(clk), .Q(n17768) );
  HS65_LH_DFPQX4 clk_r_REG739_S4 ( .D(n7008), .CP(clk), .Q(n17952) );
  HS65_LH_DFPQX4 clk_r_REG735_S4 ( .D(n9821), .CP(clk), .Q(n17832) );
  HS65_LH_DFPQX4 clk_r_REG731_S4 ( .D(n7365), .CP(clk), .Q(n17939) );
  HS65_LH_DFPQX4 clk_r_REG727_S4 ( .D(n9739), .CP(clk), .Q(n17834) );
  HS65_LH_DFPQX4 clk_r_REG723_S4 ( .D(n7989), .CP(clk), .Q(n17913) );
  HS65_LH_DFPQX4 clk_r_REG720_S4 ( .D(n9669), .CP(clk), .Q(n17837) );
  HS65_LH_DFPQX4 clk_r_REG716_S4 ( .D(n5950), .CP(clk), .Q(n17994) );
  HS65_LH_DFPQX4 clk_r_REG705_S4 ( .D(n9584), .CP(clk), .Q(n17840) );
  HS65_LH_DFPQX4 clk_r_REG560_S2 ( .D(n15514), .CP(clk), .Q(n17601) );
  HS65_LH_DFPQX4 clk_r_REG559_S2 ( .D(n15493), .CP(clk), .Q(n17591) );
  HS65_LH_DFPQX4 clk_r_REG564_S2 ( .D(n15397), .CP(clk), .Q(n17600) );
  HS65_LH_DFPQX4 clk_r_REG563_S2 ( .D(n15715), .CP(clk), .Q(n17590) );
  HS65_LH_DFPQX4 clk_r_REG309_S4 ( .D(n3593), .CP(clk), .Q(n18051) );
  HS65_LH_DFPQX4 clk_r_REG911_S1 ( .D(n9583), .CP(clk), .Q(n17841) );
  HS65_LH_DFPQX4 clk_r_REG619_S2 ( .D(n10373), .CP(clk), .Q(n17771) );
  HS65_LH_DFPQX4 clk_r_REG877_S4 ( .D(n11620), .CP(clk), .Q(n17742) );
  HS65_LH_DFPQX4 clk_r_REG687_S4 ( .D(n8098), .CP(clk), .Q(n17905) );
  HS65_LH_DFPQX4 clk_r_REG567_S2 ( .D(n14230), .CP(clk), .Q(n17474) );
  HS65_LH_DFPQX4 clk_r_REG691_S4 ( .D(n6898), .CP(clk), .Q(n17956) );
  HS65_LH_DFPQX4 clk_r_REG744_S4 ( .D(n9870), .CP(clk), .Q(n17828) );
  HS65_LH_DFPQX4 clk_r_REG624_S3 ( .D(write_byte_snps_wire), .CP(clk), .Q(
        n17627) );
  HS65_LH_DFPQX4 clk_r_REG1_S1 ( .D(n8449), .CP(clk), .Q(n17891) );
  HS65_LH_DFPQX4 clk_r_REG554_S2 ( .D(n15414), .CP(clk), .Q(n17515) );
  HS65_LH_DFPQX4 clk_r_REG566_S2 ( .D(n14966), .CP(clk), .Q(n17470) );
  HS65_LH_DFPQX4 clk_r_REG683_S1 ( .D(n7499), .CP(clk), .Q(n17932) );
  HS65_LH_DFPQX4 clk_r_REG676_S1 ( .D(n6446), .CP(clk), .Q(n17975) );
  HS65_LH_DFPQX4 clk_r_REG634_S2 ( .D(n14046), .CP(clk), .Q(n17636) );
  HS65_LH_DFPQX4 clk_r_REG555_S2 ( .D(n15506), .CP(clk), .Q(n17592) );
  HS65_LH_DFPQX4 clk_r_REG665_S1 ( .D(n8665), .CP(clk), .Q(n17882) );
  HS65_LH_DFPQX4 clk_r_REG671_S1 ( .D(n8926), .CP(clk), .Q(n17871) );
  HS65_LH_DFPQX4 clk_r_REG301_S4 ( .D(n3643), .CP(clk), .Q(n18049) );
  HS65_LH_DFPQX4 clk_r_REG638_S1 ( .D(n9292), .CP(clk), .Q(n17854) );
  HS65_LH_DFPQX4 clk_r_REG869_S2 ( .D(n9871), .CP(clk), .Q(n17827) );
  HS65_LH_DFPQX4 clk_r_REG880_S4 ( .D(n10244), .CP(clk), .Q(n17779) );
  HS65_LH_DFPQX4 clk_r_REG622_S2 ( .D(n10245), .CP(clk), .Q(n17778) );
  HS65_LH_DFPQX4 clk_r_REG870_S2 ( .D(n9868), .CP(clk), .Q(n17830) );
  HS65_LH_DFPQX4 clk_r_REG736_S5 ( .D(n9798), .CP(clk), .Q(n17833) );
  HS65_LH_DFPQX4 clk_r_REG728_S5 ( .D(n9715), .CP(clk), .Q(n17836) );
  HS65_LH_DFPQX4 clk_r_REG721_S5 ( .D(n9645), .CP(clk), .Q(n17839) );
  HS65_LH_DFPQX4 clk_r_REG706_S5 ( .D(n9560), .CP(clk), .Q(n17842) );
  HS65_LH_DFPQX4 clk_r_REG745_S5 ( .D(n10889), .CP(clk), .Q(n17753) );
  HS65_LH_DFPQX4 clk_r_REG637_S1 ( .D(n9285), .CP(clk), .Q(n17858) );
  HS65_LH_DFPQX4 clk_r_REG193_S1 ( .D(n8796), .CP(clk), .Q(n17879) );
  HS65_LH_DFPQX4 clk_r_REG158_S1 ( .D(n6576), .CP(clk), .Q(n17972) );
  HS65_LH_DFPQX4 clk_r_REG649_S4 ( .D(n10769), .CP(clk), .Q(n17754) );
  HS65_LH_DFPQX4 clk_r_REG897_S4 ( .D(n10346), .CP(clk), .Q(n17772) );
  HS65_LH_DFPQX4 clk_r_REG626_S3 ( .D(n15702), .CP(clk), .Q(n17509) );
  HS65_LH_DFPQX4 clk_r_REG627_S3 ( .D(n9286), .CP(clk), .Q(n17857) );
  HS65_LH_DFPQX4 clk_r_REG625_S3 ( .D(n10565), .CP(clk), .Q(n17763) );
  HS65_LH_DFPQX4 clk_r_REG293_S4 ( .D(n3696), .CP(clk), .Q(n18047) );
  HS65_LH_DFPQX4 clk_r_REG520_S10 ( .D(n9166), .CP(clk), .Q(n17864) );
  HS65_LH_DFPQX4 clk_r_REG111_S1 ( .D(n8229), .CP(clk), .Q(n17901) );
  HS65_LH_DFPQX4 clk_r_REG83_S1 ( .D(n7562), .CP(clk), .Q(n17930) );
  HS65_LH_DFPQX4 clk_r_REG881_S4 ( .D(n10241), .CP(clk), .Q(n17780) );
  HS65_LH_DFPQX4 clk_r_REG635_S2 ( .D(n10090), .CP(clk), .Q(n17789) );
  HS65_LH_DFPQX4 clk_r_REG630_S2 ( .D(n10103), .CP(clk), .Q(n17787) );
  HS65_LH_DFPQX4 clk_r_REG78_S10 ( .D(n9256), .CP(clk), .Q(n17860) );
  HS65_LH_DFPQX4 clk_r_REG190_S5 ( .D(\u_DataPath/dataOut_exe_i [2]), .CP(clk), 
        .Q(n17287) );
  HS65_LH_DFPQX4 clk_r_REG886_S4 ( .D(n10293), .CP(clk), .Q(n17776) );
  HS65_LH_DFPQX4 clk_r_REG883_S4 ( .D(n10270), .CP(clk), .Q(n17777) );
  HS65_LH_DFPQX4 clk_r_REG878_S4 ( .D(n10128), .CP(clk), .Q(n17786) );
  HS65_LH_DFPQX4 clk_r_REG650_S4 ( .D(n10751), .CP(clk), .Q(n17757) );
  HS65_LH_DFPQX4 clk_r_REG285_S4 ( .D(n3746), .CP(clk), .Q(n18045) );
  HS65_LH_DFPQX4 clk_r_REG895_S4 ( .D(n10321), .CP(clk), .Q(n17773) );
  HS65_LH_DFPQX4 clk_r_REG623_S3 ( .D(n14078), .CP(clk), .Q(n17524) );
  HS65_LH_DFPQX4 clk_r_REG525_S10 ( .D(n9543), .CP(clk), .Q(n17843) );
  HS65_LH_DFPQX4 clk_r_REG585_S3 ( .D(n14210), .CP(clk), .Q(n17278) );
  HS65_LH_DFPQX4 clk_r_REG489_S1 ( .D(n7154), .CP(clk), .Q(n17947) );
  HS65_LH_DFPQX4 clk_r_REG477_S1 ( .D(n9077), .CP(clk), .Q(n17868) );
  HS65_LH_DFPQX4 clk_r_REG521_S10 ( .D(n9163), .CP(clk), .Q(n17865) );
  HS65_LH_DFPQX4 clk_r_REG194_S1 ( .D(n8792), .CP(clk), .Q(n17880) );
  HS65_LH_DFPQX4 clk_r_REG84_S1 ( .D(n7559), .CP(clk), .Q(n17931) );
  HS65_LH_DFPQX4 clk_r_REG513_S4 ( .D(n2822), .CP(clk), .Q(n18089) );
  HS65_LH_DFPQX4 clk_r_REG500_S12 ( .D(n2773), .CP(clk), .Q(n18092) );
  HS65_LH_DFPQX4 clk_r_REG79_S10 ( .D(n9252), .CP(clk), .Q(n17861) );
  HS65_LH_DFPQX4 clk_r_REG159_S1 ( .D(n6572), .CP(clk), .Q(n17973) );
  HS65_LH_DFPQX4 clk_r_REG112_S1 ( .D(n8226), .CP(clk), .Q(n17902) );
  HS65_LH_DFPQX4 clk_r_REG887_S4 ( .D(n10488), .CP(clk), .Q(n17765) );
  HS65_LH_DFPQX4 clk_r_REG632_S2 ( .D(n10065), .CP(clk), .Q(n17790) );
  HS65_LH_DFPQX4 clk_r_REG460_S4 ( .D(n4212), .CP(clk), .Q(n18022) );
  HS65_LH_DFPQX4 clk_r_REG450_S2 ( .D(n2922), .CP(clk), .Q(n18083) );
  HS65_LH_DFPQX4 clk_r_REG443_S4 ( .D(n4324), .CP(clk), .Q(n18017) );
  HS65_LH_DFPQX4 clk_r_REG434_S4 ( .D(n2870), .CP(clk), .Q(n18087) );
  HS65_LH_DFPQX4 clk_r_REG424_S4 ( .D(n2976), .CP(clk), .Q(n18079) );
  HS65_LH_DFPQX4 clk_r_REG415_S4 ( .D(n3027), .CP(clk), .Q(n18076) );
  HS65_LH_DFPQX4 clk_r_REG405_S4 ( .D(n3079), .CP(clk), .Q(n18074) );
  HS65_LH_DFPQX4 clk_r_REG393_S4 ( .D(n3130), .CP(clk), .Q(n18071) );
  HS65_LH_DFPQX4 clk_r_REG382_S4 ( .D(n3182), .CP(clk), .Q(n18069) );
  HS65_LH_DFPQX4 clk_r_REG375_S6 ( .D(n3233), .CP(clk), .Q(n18066) );
  HS65_LH_DFPQX4 clk_r_REG365_S4 ( .D(n3285), .CP(clk), .Q(n18064) );
  HS65_LH_DFPQX4 clk_r_REG354_S5 ( .D(n3336), .CP(clk), .Q(n18061) );
  HS65_LH_DFPQX4 clk_r_REG342_S4 ( .D(n3388), .CP(clk), .Q(n18059) );
  HS65_LH_DFPQX4 clk_r_REG335_S4 ( .D(n3439), .CP(clk), .Q(n18057) );
  HS65_LH_DFPQX4 clk_r_REG324_S4 ( .D(n3491), .CP(clk), .Q(n18054) );
  HS65_LH_DFPQX4 clk_r_REG315_S4 ( .D(n3542), .CP(clk), .Q(n18052) );
  HS65_LH_DFPQX4 clk_r_REG307_S4 ( .D(n3594), .CP(clk), .Q(n18050) );
  HS65_LH_DFPQX4 clk_r_REG299_S4 ( .D(n3645), .CP(clk), .Q(n18048) );
  HS65_LH_DFPQX4 clk_r_REG291_S4 ( .D(n3697), .CP(clk), .Q(n18046) );
  HS65_LH_DFPQX4 clk_r_REG283_S4 ( .D(n3748), .CP(clk), .Q(n18044) );
  HS65_LH_DFPQX4 clk_r_REG196_S3 ( .D(n10155), .CP(clk), .Q(n17783) );
  HS65_LH_DFPQX4 clk_r_REG586_S3 ( .D(n14034), .CP(clk), .Q(n17631) );
  HS65_LH_DFPQX4 clk_r_REG277_S4 ( .D(n3799), .CP(clk), .Q(n18043) );
  HS65_LH_DFPQX4 clk_r_REG155_S4 ( .D(\u_DataPath/dataOut_exe_i [3]), .CP(clk), 
        .Q(n17288) );
  HS65_LH_DFPQX4 clk_r_REG888_S4 ( .D(n10485), .CP(clk), .Q(n17767) );
  HS65_LH_DFPQX4 clk_r_REG275_S4 ( .D(n3800), .CP(clk), .Q(n18042) );
  HS65_LH_DFPQX4 clk_r_REG576_S2 ( .D(n10015), .CP(clk), .Q(n17792) );
  HS65_LH_DFPQX4 clk_r_REG116_S1 ( .D(n7946), .CP(clk), .Q(n17915) );
  HS65_LH_DFPQX4 clk_r_REG5_S1 ( .D(n8406), .CP(clk), .Q(n17894) );
  HS65_LH_DFPQX4 clk_r_REG577_S3 ( .D(n15207), .CP(clk), .Q(n17312) );
  HS65_LH_DFPQX4 clk_r_REG34_S1 ( .D(n6745), .CP(clk), .Q(n17964) );
  HS65_LH_DFPQX4 clk_r_REG29_S1 ( .D(n7645), .CP(clk), .Q(n17926) );
  HS65_LH_DFPQX4 clk_r_REG187_S1 ( .D(n5908), .CP(clk), .Q(n17995) );
  HS65_LH_DFPQX4 clk_r_REG177_S1 ( .D(n8054), .CP(clk), .Q(n17908) );
  HS65_LH_DFPQX4 clk_r_REG142_S1 ( .D(n6402), .CP(clk), .Q(n17977) );
  HS65_LH_DFPQX4 clk_r_REG126_S1 ( .D(n7838), .CP(clk), .Q(n17919) );
  HS65_LH_DFPQX4 clk_r_REG122_S1 ( .D(n7455), .CP(clk), .Q(n17934) );
  HS65_LH_DFPQX4 clk_r_REG101_S1 ( .D(n6856), .CP(clk), .Q(n17957) );
  HS65_LH_DFPQX4 clk_r_REG24_S1 ( .D(n8881), .CP(clk), .Q(n17874) );
  HS65_LH_DFPQX4 clk_r_REG18_S1 ( .D(n8622), .CP(clk), .Q(n17884) );
  HS65_LH_DFPQX4 clk_r_REG269_S4 ( .D(n3849), .CP(clk), .Q(n18041) );
  HS65_LH_DFPQX4 clk_r_REG108_S8 ( .D(\u_DataPath/dataOut_exe_i [4]), .CP(clk), 
        .Q(n17289) );
  HS65_LH_DFPQX4 clk_r_REG587_S3 ( .D(n14239), .CP(clk), .Q(n17612) );
  HS65_LH_DFPQX4 clk_r_REG191_S5 ( .D(Address_toRAM_0), .CP(clk), .Q(n17459)
         );
  HS65_LH_DFPQX4 clk_r_REG156_S4 ( .D(Address_toRAM_1), .CP(clk), .Q(n17483)
         );
  HS65_LH_DFPQX4 clk_r_REG94_S5 ( .D(\u_DataPath/dataOut_exe_i [8]), .CP(clk), 
        .Q(n17290) );
  HS65_LH_DFPQX4 clk_r_REG131_S1 ( .D(n7322), .CP(clk), .Q(n17940) );
  HS65_LH_DFPQX4 clk_r_REG38_S1 ( .D(n6964), .CP(clk), .Q(n17954) );
  HS65_LH_DFPQX4 clk_r_REG152_S1 ( .D(n8513), .CP(clk), .Q(n17889) );
  HS65_LH_DFPQX4 clk_r_REG267_S4 ( .D(n3851), .CP(clk), .Q(n18040) );
  HS65_LH_DFPQX4 clk_r_REG448_S3 ( .D(n8272), .CP(clk), .Q(n17899) );
  HS65_LH_DFPQX4 clk_r_REG104_S7 ( .D(\u_DataPath/dataOut_exe_i [7]), .CP(clk), 
        .Q(n17366) );
  HS65_LH_DFPQX4 clk_r_REG578_S3 ( .D(n14256), .CP(clk), .Q(n17616) );
  HS65_LH_DFPQX4 clk_r_REG262_S4 ( .D(n3902), .CP(clk), .Q(n18038) );
  HS65_LH_DFPQX4 clk_r_REG97_S1 ( .D(n8311), .CP(clk), .Q(n17898) );
  HS65_LH_DFPQX4 clk_r_REG495_S1 ( .D(n7750), .CP(clk), .Q(n17923) );
  HS65_LH_DFPQX4 clk_r_REG493_S1 ( .D(n6657), .CP(clk), .Q(n17969) );
  HS65_LH_DFPQX4 clk_r_REG481_S1 ( .D(n7237), .CP(clk), .Q(n17944) );
  HS65_LH_DFPQX4 clk_r_REG475_S1 ( .D(n6314), .CP(clk), .Q(n17981) );
  HS65_LH_DFPQX4 clk_r_REG473_S1 ( .D(n7071), .CP(clk), .Q(n17950) );
  HS65_LH_DFPQX4 clk_r_REG470_S1 ( .D(n6230), .CP(clk), .Q(n17984) );
  HS65_LH_DFPQX4 clk_r_REG81_S11 ( .D(\u_DataPath/dataOut_exe_i [5]), .CP(clk), 
        .Q(n17364) );
  HS65_LH_DFPQX4 clk_r_REG132_S1 ( .D(n7320), .CP(clk), .Q(n17941) );
  HS65_LH_DFPQX4 clk_r_REG39_S1 ( .D(n6962), .CP(clk), .Q(n17955) );
  HS65_LH_DFPQX4 clk_r_REG117_S1 ( .D(n7942), .CP(clk), .Q(n17916) );
  HS65_LH_DFPQX4 clk_r_REG35_S1 ( .D(n6742), .CP(clk), .Q(n17965) );
  HS65_LH_DFPQX4 clk_r_REG30_S1 ( .D(n7642), .CP(clk), .Q(n17927) );
  HS65_LH_DFPQX4 clk_r_REG153_S1 ( .D(n8511), .CP(clk), .Q(n17890) );
  HS65_LH_DFPQX4 clk_r_REG188_S1 ( .D(n5905), .CP(clk), .Q(n17996) );
  HS65_LH_DFPQX4 clk_r_REG178_S1 ( .D(n8051), .CP(clk), .Q(n17909) );
  HS65_LH_DFPQX4 clk_r_REG143_S1 ( .D(n6399), .CP(clk), .Q(n17978) );
  HS65_LH_DFPQX4 clk_r_REG127_S1 ( .D(n7835), .CP(clk), .Q(n17920) );
  HS65_LH_DFPQX4 clk_r_REG123_S1 ( .D(n7452), .CP(clk), .Q(n17935) );
  HS65_LH_DFPQX4 clk_r_REG102_S1 ( .D(n6853), .CP(clk), .Q(n17958) );
  HS65_LH_DFPQX4 clk_r_REG25_S1 ( .D(n8878), .CP(clk), .Q(n17875) );
  HS65_LH_DFPQX4 clk_r_REG19_S1 ( .D(n8619), .CP(clk), .Q(n17885) );
  HS65_LH_DFPQX4 clk_r_REG6_S1 ( .D(n8402), .CP(clk), .Q(n17895) );
  HS65_LH_DFPQX4 clk_r_REG357_S1 ( .D(n6145), .CP(clk), .Q(n17988) );
  HS65_LH_DFPQX4 clk_r_REG109_S8 ( .D(\Address_toRAM[2]_snps_wire ), .CP(clk), 
        .Q(n18148) );
  HS65_LH_DFPQX4 clk_r_REG526_S10 ( .D(n9524), .CP(clk), .Q(n17845) );
  HS65_LH_DFPQX4 clk_r_REG95_S5 ( .D(\Address_toRAM[6]_snps_wire ), .CP(clk), 
        .Q(n18149) );
  HS65_LH_DFPQX4 clk_r_REG579_S3 ( .D(n14272), .CP(clk), .Q(n17615) );
  HS65_LH_DFPQX4 clk_r_REG258_S4 ( .D(n3903), .CP(clk), .Q(n18037) );
  HS65_LH_DFPQX4 clk_r_REG441_S3 ( .D(n7604), .CP(clk), .Q(n17928) );
  HS65_LH_DFPQX4 clk_r_REG590_S3 ( .D(n14238), .CP(clk), .Q(n17476) );
  HS65_LH_DFPQX4 clk_r_REG582_S3 ( .D(n15209), .CP(clk), .Q(n17479) );
  HS65_LH_DFPQX4 clk_r_REG161_S3 ( .D(\u_DataPath/dataOut_exe_i [6]), .CP(clk), 
        .Q(n17365) );
  HS65_LH_DFPQX4 clk_r_REG588_S3 ( .D(n14141), .CP(clk), .Q(n17477) );
  HS65_LH_DFPQX4 clk_r_REG105_S7 ( .D(\Address_toRAM[5]_snps_wire ), .CP(clk), 
        .Q(n18147) );
  HS65_LH_DFPQX4 clk_r_REG432_S3 ( .D(n9014), .CP(clk), .Q(n17869) );
  HS65_LH_DFPQX4 clk_r_REG583_S3 ( .D(n14257), .CP(clk), .Q(n17618) );
  HS65_LH_DFPQX4 clk_r_REG252_S4 ( .D(n3952), .CP(clk), .Q(n18036) );
  HS65_LH_DFPQX4 clk_r_REG86_S3 ( .D(\u_DataPath/dataOut_exe_i [9]), .CP(clk), 
        .Q(n17291) );
  HS65_LH_DFPQX4 clk_r_REG580_S3 ( .D(n15208), .CP(clk), .Q(n17478) );
  HS65_LH_DFPQX4 clk_r_REG458_S3 ( .D(n6618), .CP(clk), .Q(n17970) );
  HS65_LH_DFPQX4 clk_r_REG591_S3 ( .D(n14242), .CP(clk), .Q(n17610) );
  HS65_LH_DFPQX4 clk_r_REG581_S3 ( .D(n14206), .CP(clk), .Q(n17614) );
  HS65_LH_DFPQX4 clk_r_REG498_S11 ( .D(\Address_toRAM[3]_snps_wire ), .CP(clk), 
        .Q(n18137) );
  HS65_LH_DFPQX4 clk_r_REG250_S4 ( .D(n3954), .CP(clk), .Q(n18035) );
  HS65_LH_DFPQX4 clk_r_REG584_S3 ( .D(n14274), .CP(clk), .Q(n17617) );
  HS65_LH_DFPQX4 clk_r_REG589_S3 ( .D(n14240), .CP(clk), .Q(n17611) );
  HS65_LH_DFPQX4 clk_r_REG107_S7 ( .D(n14613), .CP(clk), .Q(n17254) );
  HS65_LH_DFPQX4 clk_r_REG98_S5 ( .D(n15240), .CP(clk), .Q(n17260) );
  HS65_LH_DFPQX4 clk_r_REG89_S3 ( .D(n14785), .CP(clk), .Q(n17256) );
  HS65_LH_DFPQX4 clk_r_REG162_S3 ( .D(\Address_toRAM[4]_snps_wire ), .CP(clk), 
        .Q(n18150) );
  HS65_LH_DFPQX4 clk_r_REG160_S4 ( .D(n14220), .CP(clk), .Q(n17257) );
  HS65_LH_DFPQX4 clk_r_REG113_S8 ( .D(n14224), .CP(clk), .Q(n17259) );
  HS65_LH_DFPQX4 clk_r_REG244_S4 ( .D(n4005), .CP(clk), .Q(n18033) );
  HS65_LH_DFPQX4 clk_r_REG164_S3 ( .D(n15136), .CP(clk), .Q(n17251) );
  HS65_LH_DFPQX4 clk_r_REG87_S3 ( .D(\Address_toRAM[7]_snps_wire ), .CP(clk), 
        .Q(n18153) );
  HS65_LH_DFPQX4 clk_r_REG240_S4 ( .D(n4006), .CP(clk), .Q(n18032) );
  HS65_LH_DFPQX4 clk_r_REG90_S4 ( .D(\u_DataPath/dataOut_exe_i [10]), .CP(clk), 
        .Q(n17292) );
  HS65_LH_DFPQX4 clk_r_REG422_S3 ( .D(n7199), .CP(clk), .Q(n17945) );
  HS65_LH_DFPQX4 clk_r_REG137_S4 ( .D(n33213), .CP(clk), .Q(n17462) );
  HS65_LH_DFPQX4 clk_r_REG165_S3 ( .D(n4376), .CP(clk), .Q(n18016) );
  HS65_LH_DFPQX4 clk_r_REG234_S4 ( .D(n4055), .CP(clk), .Q(n18031) );
  HS65_LH_DFPQX4 clk_r_REG91_S4 ( .D(\Address_toRAM[8]_snps_wire ), .CP(clk), 
        .Q(n17520) );
  HS65_LH_DFPQX4 clk_r_REG93_S4 ( .D(n14409), .CP(clk), .Q(n17253) );
  HS65_LH_DFPQX4 clk_r_REG232_S4 ( .D(n4057), .CP(clk), .Q(n18030) );
  HS65_LH_DFPQX4 clk_r_REG398_S3 ( .D(n15621), .CP(clk), .Q(n17270) );
  HS65_LH_DFPQX4 clk_r_REG403_S3 ( .D(n14200), .CP(clk), .Q(n17277) );
  HS65_LH_DFPQX4 clk_r_REG413_S3 ( .D(n8366), .CP(clk), .Q(n17896) );
  HS65_LH_DFPQX4 clk_r_REG138_S4 ( .D(n33052), .CP(clk), .Q(n17308) );
  HS65_LH_DFPQX4 clk_r_REG166_S4 ( .D(\u_DataPath/dataOut_exe_i [11]), .CP(clk), .Q(n17293) );
  HS65_LH_DFPQX4 clk_r_REG505_S3 ( .D(n11595), .CP(clk), .Q(n17743) );
  HS65_LH_DFPQX4 clk_r_REG515_S3 ( .D(n9208), .CP(clk), .Q(n17863) );
  HS65_LH_DFPQX4 clk_r_REG222_S4 ( .D(n4109), .CP(clk), .Q(n18027) );
  HS65_LH_DFPQX4 clk_r_REG538_S9 ( .D(n9284), .CP(clk), .Q(n17859) );
  HS65_LH_DFPQX4 clk_r_REG226_S4 ( .D(n4108), .CP(clk), .Q(n18028) );
  HS65_LH_DFPQX4 clk_r_REG334_S3 ( .D(n15053), .CP(clk), .Q(n17466) );
  HS65_LH_DFPQX4 clk_r_REG438_S3 ( .D(n11495), .CP(clk), .Q(n17748) );
  HS65_LH_DFPQX4 clk_r_REG169_S4 ( .D(n14616), .CP(clk), .Q(n17252) );
  HS65_LH_DFPQX4 clk_r_REG419_S3 ( .D(n11456), .CP(clk), .Q(n17750) );
  HS65_LH_DFPQX4 clk_r_REG442_S3 ( .D(n5116), .CP(clk), .Q(n18005) );
  HS65_LH_DFPQX4 clk_r_REG423_S3 ( .D(n5367), .CP(clk), .Q(n18001) );
  HS65_LH_DFPQX4 clk_r_REG399_S3 ( .D(n11417), .CP(clk), .Q(n17752) );
  HS65_LH_DFPQX4 clk_r_REG404_S3 ( .D(n5003), .CP(clk), .Q(n18007) );
  HS65_LH_DFPQX4 clk_r_REG456_S3 ( .D(n11534), .CP(clk), .Q(n17746) );
  HS65_LH_DFPQX4 clk_r_REG459_S3 ( .D(n6543), .CP(clk), .Q(n17974) );
  HS65_LH_DFPQX4 clk_r_REG323_S3 ( .D(n15123), .CP(clk), .Q(n17465) );
  HS65_LH_DFPQX4 clk_r_REG446_S1 ( .D(n11514), .CP(clk), .Q(n17747) );
  HS65_LH_DFPQX4 clk_r_REG430_S3 ( .D(n11475), .CP(clk), .Q(n17749) );
  HS65_LH_DFPQX4 clk_r_REG433_S3 ( .D(n4393), .CP(clk), .Q(n18015) );
  HS65_LH_DFPQX4 clk_r_REG411_S3 ( .D(n11436), .CP(clk), .Q(n17751) );
  HS65_LH_DFPQX4 clk_r_REG449_S1 ( .D(n8198), .CP(clk), .Q(n17904) );
  HS65_LH_DFPQX4 clk_r_REG414_S3 ( .D(n4736), .CP(clk), .Q(n18011) );
  HS65_LH_DFPQX4 clk_r_REG507_S3 ( .D(n11573), .CP(clk), .Q(n17744) );
  HS65_LH_DFPQX4 clk_r_REG512_S3 ( .D(n9122), .CP(clk), .Q(n17866) );
  HS65_LH_DFPQX4 clk_r_REG464_S3 ( .D(n11553), .CP(clk), .Q(n17745) );
  HS65_LH_DFPQX4 clk_r_REG208_S4 ( .D(n4160), .CP(clk), .Q(n18025) );
  HS65_LH_DFPQX4 clk_r_REG467_S3 ( .D(n8756), .CP(clk), .Q(n17881) );
  HS65_LH_DFPQX4 clk_r_REG167_S4 ( .D(\Address_toRAM[9]_snps_wire ), .CP(clk), 
        .Q(n18151) );
  HS65_LH_DFPQX4 clk_r_REG216_S4 ( .D(n4158), .CP(clk), .Q(n18026) );
  HS65_LH_DFPQX4 clk_r_REG402_S3 ( .D(n7796), .CP(clk), .Q(n17921) );
  HS65_LH_DFPQX4 clk_r_REG352_S3 ( .D(n6217), .CP(clk), .Q(n17985) );
  HS65_LH_DFPQX4 clk_r_REG381_S3 ( .D(n6369), .CP(clk), .Q(n17979) );
  HS65_LH_DFPQX4 clk_r_REG374_S3 ( .D(n7132), .CP(clk), .Q(n17948) );
  HS65_LH_DFPQX4 clk_r_REG392_S3 ( .D(n6708), .CP(clk), .Q(n17966) );
  HS65_LH_DFPQX4 clk_r_REG341_S3 ( .D(n6305), .CP(clk), .Q(n17982) );
  HS65_LH_DFPQX4 clk_r_REG364_S3 ( .D(n7302), .CP(clk), .Q(n17942) );
  HS65_LH_DFPQX4 clk_r_REG333_S3 ( .D(n8612), .CP(clk), .Q(n17886) );
  HS65_LH_DFPQX4 clk_r_REG170_S5 ( .D(\u_DataPath/dataOut_exe_i [12]), .CP(clk), .Q(n17367) );
  HS65_LH_DFPQX4 clk_r_REG210_S4 ( .D(n4272), .CP(clk), .Q(n18019) );
  HS65_LH_DFPQX4 clk_r_REG192_S5 ( .D(n8812), .CP(clk), .Q(n17878) );
  HS65_LH_DFPQX4 clk_r_REG215_S4 ( .D(n4271), .CP(clk), .Q(n18020) );
  HS65_LH_DFPQX4 clk_r_REG173_S5 ( .D(n15238), .CP(clk), .Q(n17250) );
  HS65_LH_DFPQX4 clk_r_REG145_S10 ( .D(\u_DataPath/dataOut_exe_i [13]), .CP(
        clk), .Q(n17368) );
  HS65_LH_DFPQX4 clk_r_REG171_S5 ( .D(\Address_toRAM[10]_snps_wire ), .CP(clk), 
        .Q(n18154) );
  HS65_LH_DFPQX4 clk_r_REG148_S10 ( .D(n14631), .CP(clk), .Q(n17255) );
  HS65_LH_DFPQX4 clk_r_REG146_S10 ( .D(\Address_toRAM[11]_snps_wire ), .CP(clk), .Q(n18152) );
  HS65_LH_DFPQX4 clk_r_REG537_S9 ( .D(n10726), .CP(clk), .Q(n17759) );
  HS65_LH_DFPQX4 clk_r_REG157_S4 ( .D(n6592), .CP(clk), .Q(n17971) );
  HS65_LH_DFPQX4 clk_r_REG96_S5 ( .D(n8337), .CP(clk), .Q(n17897) );
  HS65_LH_DFPQX4 clk_r_REG110_S8 ( .D(n8246), .CP(clk), .Q(n17900) );
  HS65_LH_DFPQX4 clk_r_REG106_S7 ( .D(n7174), .CP(clk), .Q(n17946) );
  HS65_LH_DFPQX4 clk_r_REG82_S11 ( .D(n7579), .CP(clk), .Q(n17929) );
  HS65_LH_DFPQX4 clk_r_REG180_S3 ( .D(\u_DataPath/dataOut_exe_i [15]), .CP(clk), .Q(n17369) );
  HS65_LH_DFPQX4 clk_r_REG15_S3 ( .D(\u_DataPath/dataOut_exe_i [17]), .CP(clk), 
        .Q(n17261) );
  HS65_LH_DFPQX4 clk_r_REG149_S3 ( .D(\u_DataPath/dataOut_exe_i [16]), .CP(clk), .Q(n17370) );
  HS65_LH_DFPQX4 clk_r_REG88_S3 ( .D(n7770), .CP(clk), .Q(n17922) );
  HS65_LH_DFPQX4 clk_r_REG163_S3 ( .D(n8988), .CP(clk), .Q(n17870) );
  HS65_LH_DFPQX4 clk_r_REG99_S6 ( .D(n32607), .CP(clk), .Q(n17318) );
  HS65_LH_DFPQX4 clk_r_REG181_S3 ( .D(Address_toRAM_13), .CP(clk), .Q(n17488)
         );
  HS65_LH_DFPQX4 clk_r_REG16_S3 ( .D(Address_toRAM_15), .CP(clk), .Q(n17487)
         );
  HS65_LH_DFPQX4 clk_r_REG150_S3 ( .D(Address_toRAM_14), .CP(clk), .Q(n17485)
         );
  HS65_LH_DFPQX4 clk_r_REG183_S3 ( .D(n14338), .CP(clk), .Q(n17248) );
  HS65_LH_DFPQX4 clk_r_REG184_S3 ( .D(n6041), .CP(clk), .Q(n17989) );
  HS65_LH_DFPQX4 clk_r_REG92_S4 ( .D(n6677), .CP(clk), .Q(n17968) );
  HS65_LH_DFPQX4 clk_r_REG21_S3 ( .D(\u_DataPath/dataOut_exe_i [18]), .CP(clk), 
        .Q(n17262) );
  HS65_LH_DFPQX4 clk_r_REG516_S4 ( .D(n10704), .CP(clk), .Q(n17761) );
  HS65_LH_DFPQX4 clk_r_REG8_S3 ( .D(n32487), .CP(clk), .Q(n17271) );
  HS65_LH_DFPQX4 clk_r_REG22_S3 ( .D(Address_toRAM_16), .CP(clk), .Q(n17486)
         );
  HS65_LH_DFPQX4 clk_r_REG168_S4 ( .D(n6334), .CP(clk), .Q(n17980) );
  HS65_LH_DFPQX4 clk_r_REG27_S3 ( .D(n32469), .CP(clk), .Q(n17273) );
  HS65_LH_DFPQX4 clk_r_REG80_S10 ( .D(n14217), .CP(clk), .Q(n17258) );
  HS65_LH_DFPQX4 clk_r_REG517_S9 ( .D(n15750), .CP(clk), .Q(n17313) );
  HS65_LH_DFPQX4 clk_r_REG73_S9 ( .D(\Data_in[28]_snps_wire ), .CP(clk), .Q(
        n17522) );
  HS65_LH_DFPQX4 clk_r_REG72_S9 ( .D(\Data_in[31]_snps_wire ), .CP(clk), .Q(
        n17521) );
  HS65_LH_DFPQX4 clk_r_REG71_S9 ( .D(\Data_in[27]_snps_wire ), .CP(clk), .Q(
        n17519) );
  HS65_LH_DFPQX4 clk_r_REG70_S9 ( .D(Data_in_23), .CP(clk), .Q(n17455) );
  HS65_LH_DFPQX4 clk_r_REG69_S9 ( .D(Data_in_24), .CP(clk), .Q(n17456) );
  HS65_LH_DFPQX4 clk_r_REG68_S9 ( .D(Data_in_25), .CP(clk), .Q(n17457) );
  HS65_LH_DFPQX4 clk_r_REG67_S9 ( .D(Data_in_26), .CP(clk), .Q(n17458) );
  HS65_LH_DFPQX4 clk_r_REG139_S4 ( .D(\u_DataPath/dataOut_exe_i [19]), .CP(clk), .Q(n17371) );
  HS65_LH_DFPQX4 clk_r_REG534_S4 ( .D(n9314), .CP(clk), .Q(n17852) );
  HS65_LH_DFPQX4 clk_r_REG32_S4 ( .D(n32137), .CP(clk), .Q(n17275) );
  HS65_LH_DFPQX4 clk_r_REG140_S4 ( .D(Address_toRAM_17), .CP(clk), .Q(n17484)
         );
  HS65_LH_DFPQX4 clk_r_REG75_S9 ( .D(\Data_in[30]_snps_wire ), .CP(clk), .Q(
        n18139) );
  HS65_LH_DFPQX4 clk_r_REG74_S9 ( .D(\Data_in[29]_snps_wire ), .CP(clk), .Q(
        n18138) );
  HS65_LH_DFPQX4 clk_r_REG76_S9 ( .D(n17198), .CP(clk), .Q(n17454) );
  HS65_LH_DFPQX4 clk_r_REG536_S4 ( .D(\nibble[0]_snps_wire ), .CP(clk), .Q(
        n18127) );
  HS65_LH_DFPQX4 clk_r_REG530_S4 ( .D(n288), .CP(clk), .Q(n17281) );
  HS65_LH_DFPQX4 clk_r_REG77_S9 ( .D(\nibble[1]_snps_wire ), .CP(clk), .Q(
        n17453) );
  HS65_LH_DFPQX4 clk_r_REG535_S4 ( .D(n17199), .CP(clk), .Q(n17376) );
  HS65_LH_DFPQX4 clk_r_REG518_S9 ( .D(n17197), .CP(clk), .Q(n17505) );
  HS65_LH_DFPQX4 clk_r_REG172_S5 ( .D(n7091), .CP(clk), .Q(n17949) );
  HS65_LH_DFPQX4 clk_r_REG51_S9 ( .D(write_op_snps_wire), .CP(clk), .Q(n17510)
         );
  HS65_LH_DFPQX4 clk_r_REG185_S4 ( .D(n32079), .CP(clk), .Q(n17276) );
  HS65_LH_DFPQX4 clk_r_REG519_S9 ( .D(n312), .CP(clk), .Q(n17568) );
  HS65_LH_DFPQX4 clk_r_REG58_S9 ( .D(Data_in_0), .CP(clk), .Q(n17491) );
  HS65_LH_DFPQX4 clk_r_REG57_S9 ( .D(Data_in_3), .CP(clk), .Q(n17452) );
  HS65_LH_DFPQX4 clk_r_REG56_S9 ( .D(Data_in_4), .CP(clk), .Q(n17451) );
  HS65_LH_DFPQX4 clk_r_REG55_S9 ( .D(Data_in_1), .CP(clk), .Q(n17450) );
  HS65_LH_DFPQX4 clk_r_REG54_S9 ( .D(Data_in_2), .CP(clk), .Q(n17449) );
  HS65_LH_DFPQX4 clk_r_REG53_S9 ( .D(Data_in_5), .CP(clk), .Q(n17448) );
  HS65_LH_DFPQX4 clk_r_REG52_S9 ( .D(Data_in_6), .CP(clk), .Q(n17447) );
  HS65_LH_DFPQX4 clk_r_REG533_S4 ( .D(read_op_snps_wire), .CP(clk), .Q(n18155)
         );
  HS65_LH_DFPQX4 clk_r_REG119_S10 ( .D(\u_DataPath/dataOut_exe_i [21]), .CP(
        clk), .Q(n17372) );
  HS65_LH_DFPQX4 clk_r_REG2_S2 ( .D(\u_DataPath/dataOut_exe_i [20]), .CP(clk), 
        .Q(n17263) );
  HS65_LH_DFPQX4 clk_r_REG531_S4 ( .D(n9307), .CP(clk), .Q(n17853) );
  HS65_LH_DFPQX4 clk_r_REG147_S10 ( .D(n7257), .CP(clk), .Q(n17943) );
  HS65_LH_DFPQX4 clk_r_REG355_S4 ( .D(Address_toRAM_12), .CP(clk), .Q(n17460)
         );
  HS65_LH_DFPQX4 clk_r_REG353_S4 ( .D(n14365), .CP(clk), .Q(n17249) );
  HS65_LH_DFPQX4 clk_r_REG59_S9 ( .D(\Data_in[7]_snps_wire ), .CP(clk), .Q(
        n18136) );
  HS65_LH_DFPQX4 clk_r_REG358_S4 ( .D(n14304), .CP(clk), .Q(n17247) );
  HS65_LH_DFPQX4 clk_r_REG3_S2 ( .D(Address_toRAM_18), .CP(clk), .Q(n17461) );
  HS65_LH_DFPQX4 clk_r_REG120_S10 ( .D(Address_toRAM_19), .CP(clk), .Q(n17489)
         );
  HS65_LH_DFPQX4 clk_r_REG66_S9 ( .D(\Data_in[16]_snps_wire ), .CP(clk), .Q(
        n18140) );
  HS65_LH_DFPQX4 clk_r_REG65_S9 ( .D(\Data_in[17]_snps_wire ), .CP(clk), .Q(
        n18141) );
  HS65_LH_DFPQX4 clk_r_REG64_S9 ( .D(\Data_in[18]_snps_wire ), .CP(clk), .Q(
        n18142) );
  HS65_LH_DFPQX4 clk_r_REG63_S9 ( .D(\Data_in[19]_snps_wire ), .CP(clk), .Q(
        n18143) );
  HS65_LH_DFPQX4 clk_r_REG62_S9 ( .D(\Data_in[20]_snps_wire ), .CP(clk), .Q(
        n18144) );
  HS65_LH_DFPQX4 clk_r_REG61_S9 ( .D(\Data_in[21]_snps_wire ), .CP(clk), .Q(
        n18145) );
  HS65_LH_DFPQX4 clk_r_REG60_S9 ( .D(\Data_in[22]_snps_wire ), .CP(clk), .Q(
        n18146) );
  HS65_LH_DFPQX4 clk_r_REG50_S9 ( .D(\Data_in[11]_snps_wire ), .CP(clk), .Q(
        n18132) );
  HS65_LH_DFPQX4 clk_r_REG49_S9 ( .D(\Data_in[15]_snps_wire ), .CP(clk), .Q(
        n18135) );
  HS65_LH_DFPQX4 clk_r_REG48_S9 ( .D(\Data_in[9]_snps_wire ), .CP(clk), .Q(
        n18133) );
  HS65_LH_DFPQX4 clk_r_REG47_S9 ( .D(\Data_in[12]_snps_wire ), .CP(clk), .Q(
        n18128) );
  HS65_LH_DFPQX4 clk_r_REG46_S9 ( .D(\Data_in[13]_snps_wire ), .CP(clk), .Q(
        n18129) );
  HS65_LH_DFPQX4 clk_r_REG45_S9 ( .D(\Data_in[14]_snps_wire ), .CP(clk), .Q(
        n18134) );
  HS65_LH_DFPQX4 clk_r_REG44_S9 ( .D(\Data_in[8]_snps_wire ), .CP(clk), .Q(
        n18130) );
  HS65_LH_DFPQX4 clk_r_REG43_S9 ( .D(\Data_in[10]_snps_wire ), .CP(clk), .Q(
        n18131) );
  HS65_LH_DFPQX4 clk_r_REG129_S3 ( .D(n31402), .CP(clk), .Q(n17317) );
  HS65_LH_DFPQX4 clk_r_REG134_S4 ( .D(n31384), .CP(clk), .Q(n17274) );
  HS65_LH_DFPQX4 clk_r_REG356_S4 ( .D(n6165), .CP(clk), .Q(n17987) );
  HS65_LH_DFPQX4 clk_r_REG114_S9 ( .D(n31366), .CP(clk), .Q(n17282) );
  HS65_LH_DFPQX4 clk_r_REG136_S6 ( .D(n31350), .CP(clk), .Q(n17307) );
  HS65_LH_DFPQX4 clk_r_REG174_S6 ( .D(\u_DataPath/dataOut_exe_i [22]), .CP(clk), .Q(n17264) );
  HS65_LH_DFPQX4 clk_r_REG135_S4 ( .D(n31277), .CP(clk), .Q(n17309) );
  HS65_LH_DFPQX4 clk_r_REG115_S9 ( .D(n31366), .CP(clk), .Q(n17910) );
  HS65_LH_DFPQX4 clk_r_REG175_S6 ( .D(Address_toRAM_20), .CP(clk), .Q(n17490)
         );
  HS65_LH_DFPQX4 clk_r_REG186_S4 ( .D(n32079), .CP(clk), .Q(n17990) );
  HS65_LH_DFPQX4 clk_r_REG130_S3 ( .D(n31402), .CP(clk), .Q(n17936) );
  HS65_LH_DFPQX4 clk_r_REG33_S4 ( .D(n32137), .CP(clk), .Q(n17959) );
  HS65_LH_DFPQX4 clk_r_REG28_S3 ( .D(n32469), .CP(clk), .Q(n17924) );
  HS65_LH_DFPQX4 clk_r_REG125_S3 ( .D(n31259), .CP(clk), .Q(n17918) );
  HS65_LH_DFPQX4 clk_r_REG100_S6 ( .D(\u_DataPath/dataOut_exe_i [23]), .CP(clk), .Q(n17265) );
  HS65_LH_DFPQX4 clk_r_REG176_S6 ( .D(n8093), .CP(clk), .Q(n17907) );
  HS65_LH_DFPQX4 clk_r_REG4_S2 ( .D(n8439), .CP(clk), .Q(n17893) );
  HS65_LH_DFPQX4 clk_r_REG23_S3 ( .D(n8906), .CP(clk), .Q(n17873) );
  HS65_LH_DFPQX4 clk_r_REG17_S3 ( .D(n8641), .CP(clk), .Q(n17883) );
  HS65_LH_DFPQX4 clk_r_REG141_S4 ( .D(n6430), .CP(clk), .Q(n17976) );
  HS65_LH_DFPQX4 clk_r_REG121_S10 ( .D(n7487), .CP(clk), .Q(n17933) );
  HS65_LH_DFPQX4 clk_r_REG182_S3 ( .D(n6250), .CP(clk), .Q(n17983) );
  HS65_LH_DFPQX4 clk_r_REG151_S3 ( .D(n8531), .CP(clk), .Q(n17888) );
  HS65_LH_DFPQX9 clk_r_REG596_S2 ( .D(\u_DataPath/cw_to_ex_i [14]), .CP(clk), 
        .Q(n17528) );
  HS65_LL_DFPHQX27 clk_r_REG251_S1 ( .D(addr_to_iram_24), .E(
        \u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n18116) );
  HS65_LL_DFPHQX27 clk_r_REG233_S1 ( .D(addr_to_iram_26), .E(
        \u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n18118) );
  HS65_LL_DFPHQX27 clk_r_REG209_S1 ( .D(addr_to_iram_28), .E(
        \u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n18119) );
  HS65_LL_DFPHQX27 clk_r_REG211_S1 ( .D(addr_to_iram_29), .E(
        \u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n18120) );
  HS65_LL_DFPHQX27 clk_r_REG268_S1 ( .D(addr_to_iram_22), .E(
        \u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n18114) );
  HS65_LL_DFPHQX27 clk_r_REG440_S1 ( .D(addr_to_iram_3), .E(
        \u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n18093) );
  HS65_LL_DFPHQX27 clk_r_REG427_S1 ( .D(addr_to_iram_4), .E(
        \u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n18095) );
  HS65_LL_DFPHQX27 clk_r_REG200_S1 ( .D(addr_to_iram_2), .E(
        \u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n18094) );
  HS65_LL_DFPHQX27 clk_r_REG401_S1 ( .D(addr_to_iram_7), .E(
        \u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n18097) );
  HS65_LL_DFPHQX27 clk_r_REG421_S1 ( .D(addr_to_iram_5), .E(
        \u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n18096) );
  HS65_LL_DFPHQX27 clk_r_REG383_S1 ( .D(addr_to_iram_9), .E(
        \u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n18099) );
  HS65_LL_DFPHQX27 clk_r_REG408_S1 ( .D(addr_to_iram_6), .E(
        \u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n18098) );
  HS65_LL_DFPHQX27 clk_r_REG366_S1 ( .D(addr_to_iram_11), .E(
        \u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n18101) );
  HS65_LL_DFPHQX27 clk_r_REG387_S1 ( .D(addr_to_iram_8), .E(
        \u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n18100) );
  HS65_LL_DFPHQX27 clk_r_REG343_S1 ( .D(addr_to_iram_13), .E(
        \u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n18103) );
  HS65_LL_DFPHQX27 clk_r_REG370_S1 ( .D(addr_to_iram_10), .E(
        \u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n18102) );
  HS65_LL_DFPHQX27 clk_r_REG325_S1 ( .D(addr_to_iram_15), .E(
        \u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n18105) );
  HS65_LL_DFPHQX27 clk_r_REG347_S1 ( .D(addr_to_iram_12), .E(
        \u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n18104) );
  HS65_LL_DFPHQX27 clk_r_REG308_S1 ( .D(addr_to_iram_17), .E(
        \u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n18107) );
  HS65_LL_DFPHQX27 clk_r_REG329_S1 ( .D(addr_to_iram_14), .E(
        \u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n18106) );
  HS65_LL_DFPHQX27 clk_r_REG292_S1 ( .D(addr_to_iram_19), .E(
        \u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n18109) );
  HS65_LL_DFPHQX27 clk_r_REG316_S1 ( .D(addr_to_iram_16), .E(
        \u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n18108) );
  HS65_LL_DFPHQX27 clk_r_REG276_S1 ( .D(addr_to_iram_21), .E(
        \u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n18111) );
  HS65_LL_DFPHQX27 clk_r_REG300_S1 ( .D(addr_to_iram_18), .E(
        \u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n18110) );
  HS65_LL_DFPHQX27 clk_r_REG259_S1 ( .D(addr_to_iram_23), .E(
        \u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n18113) );
  HS65_LL_DFPHQX27 clk_r_REG284_S1 ( .D(addr_to_iram_20), .E(
        \u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n18112) );
  HS65_LL_DFPHQX27 clk_r_REG223_S1 ( .D(addr_to_iram_27), .E(
        \u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n18117) );
  HS65_LL_DFPHQX27 clk_r_REG241_S1 ( .D(addr_to_iram_25), .E(
        \u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n18115) );
  HS65_LL_DFPHQX27 clk_r_REG453_S1 ( .D(addr_to_iram_1), .E(
        \u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n18156) );
  HS65_LH_DFPHQX4 clk_r_REG278_S1 ( .D(n12087), .E(\u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n17716) );
  HS65_LH_DFPHQX4 clk_r_REG294_S1 ( .D(n11987), .E(\u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n17720) );
  HS65_LH_DFPHQX4 clk_r_REG318_S1 ( .D(n13260), .E(\u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n17658) );
  HS65_LH_DFPHQX4 clk_r_REG302_S1 ( .D(n11934), .E(\u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n17722) );
  HS65_LH_DFPHQX4 clk_r_REG270_S1 ( .D(n12138), .E(\u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n17714) );
  HS65_LH_DFPHQX4 clk_r_REG395_S1 ( .D(n12898), .E(\u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n17674) );
  HS65_LH_DFPHQX4 clk_r_REG337_S1 ( .D(n13168), .E(\u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n17662) );
  HS65_LH_DFPHQX4 clk_r_REG377_S1 ( .D(n12988), .E(\u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n17670) );
  HS65_LH_DFPHQX4 clk_r_REG360_S1 ( .D(n13078), .E(\u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n17666) );
  HS65_LH_DFPHQX4 clk_r_REG509_S1 ( .D(n12551), .E(\u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n17689) );
  HS65_LH_DFPHQX4 clk_r_REG416_S1 ( .D(n12808), .E(\u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n17678) );
  HS65_LH_DFPHQX4 clk_r_REG435_S1 ( .D(n12719), .E(\u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n17682) );
  HS65_LH_DFPHQX4 clk_r_REG501_S1 ( .D(n12504), .E(\u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n17691) );
  HS65_LH_DFPHQX4 clk_r_REG461_S1 ( .D(n12598), .E(\u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n17687) );
  HS65_LH_DFPHQX4 clk_r_REG369_S1 ( .D(n3232), .E(\u_DataPath/u_fetch/pc1/N3 ), 
        .CP(clk), .Q(n18067) );
  HS65_LH_DFPHQX4 clk_r_REG328_S1 ( .D(n3441), .E(\u_DataPath/u_fetch/pc1/N3 ), 
        .CP(clk), .Q(n18056) );
  HS65_LH_DFPHQX4 clk_r_REG452_S1 ( .D(n4210), .E(\u_DataPath/u_fetch/pc1/N3 ), 
        .CP(clk), .Q(n18024) );
  HS65_LH_DFPHQX4 clk_r_REG386_S1 ( .D(n3129), .E(\u_DataPath/u_fetch/pc1/N3 ), 
        .CP(clk), .Q(n18072) );
  HS65_LH_DFPHQX4 clk_r_REG407_S1 ( .D(n3026), .E(\u_DataPath/u_fetch/pc1/N3 ), 
        .CP(clk), .Q(n18077) );
  HS65_LH_DFPHQX4 clk_r_REG199_S1 ( .D(n2920), .E(\u_DataPath/u_fetch/pc1/N3 ), 
        .CP(clk), .Q(n18085) );
  HS65_LH_DFPHQX4 clk_r_REG346_S1 ( .D(n3335), .E(\u_DataPath/u_fetch/pc1/N3 ), 
        .CP(clk), .Q(n18062) );
  HS65_LH_DFPHQX4 clk_r_REG310_S1 ( .D(n13311), .E(\u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n17656) );
  HS65_LH_DFPHQX4 clk_r_REG286_S1 ( .D(n12036), .E(\u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n17718) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N111 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][18] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N98 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][5] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N96 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][3] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N120 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][27] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N122 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][29] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N96 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][3] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N120 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][27] ) );
  HS65_LH_DFPHQX4 clk_r_REG368_S1 ( .D(n13031), .E(\u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n17669) );
  HS65_LH_DFPSQX9 clk_r_REG902_S3 ( .D(n191), .CP(clk), .SN(n29646), .Q(n17574) );
  HS65_LH_DFPSQX9 clk_r_REG663_S3 ( .D(n15429), .CP(clk), .SN(n29697), .Q(
        n17579) );
  HS65_LH_DFPSQX9 clk_r_REG617_S1 ( .D(n15731), .CP(clk), .SN(n29651), .Q(
        n17441) );
  HS65_LH_DFPSQX9 clk_r_REG655_S3 ( .D(n217), .CP(clk), .SN(n17245), .Q(n17269) );
  HS65_LH_DFPSQX9 clk_r_REG803_S3 ( .D(n15179), .CP(clk), .SN(n29651), .Q(
        n17581) );
  HS65_LH_DFPSQX9 clk_r_REG856_S3 ( .D(n15169), .CP(clk), .SN(n40999), .Q(
        n17584) );
  HS65_LH_DFPSQX9 clk_r_REG848_S3 ( .D(n15168), .CP(clk), .SN(n18160), .Q(
        n17585) );
  HS65_LH_DFPSQX9 clk_r_REG908_S3 ( .D(n1912), .CP(clk), .SN(n29698), .Q(
        n17626) );
  HS65_LH_DFPSQX9 clk_r_REG872_S3 ( .D(n15757), .CP(clk), .SN(n17245), .Q(
        n17567) );
  HS65_LH_DFPSQX9 clk_r_REG789_S3 ( .D(n14053), .CP(clk), .SN(n18160), .Q(
        n17633) );
  HS65_LH_DFPSQX9 clk_r_REG906_S3 ( .D(n10151), .CP(clk), .SN(n29698), .Q(
        n17785) );
  HS65_LH_DFPSQX9 clk_r_REG796_S3 ( .D(n1928), .CP(clk), .SN(n18160), .Q(
        n17582) );
  HS65_LH_DFPSQX9 clk_r_REG657_S3 ( .D(n15428), .CP(clk), .SN(n29649), .Q(
        n17580) );
  HS65_LH_DFPSQX9 clk_r_REG674_S3 ( .D(n15430), .CP(clk), .SN(n40997), .Q(
        n17578) );
  HS65_LH_DFPSQX9 clk_r_REG901_S3 ( .D(n13879), .CP(clk), .SN(n29645), .Q(
        n17642) );
  HS65_LH_DFPSQX9 clk_r_REG680_S3 ( .D(n200), .CP(clk), .SN(n29698), .Q(n17437) );
  HS65_LH_DFPSQX9 clk_r_REG648_S3 ( .D(n276), .CP(clk), .SN(n29645), .Q(n17268) );
  HS65_LH_DFPSQX9 clk_r_REG602_S1 ( .D(n230), .CP(clk), .SN(n29649), .Q(n17294) );
  HS65_LH_DFPSQX9 clk_r_REG654_S3 ( .D(n240), .CP(clk), .SN(n29652), .Q(n17298) );
  HS65_LH_DFPSQX9 clk_r_REG843_S3 ( .D(n17153), .CP(clk), .SN(n29650), .Q(
        n17404) );
  HS65_LH_DFPSQX9 clk_r_REG885_S3 ( .D(n10316), .CP(clk), .SN(n40998), .Q(
        n17775) );
  HS65_LH_DFPSQX9 clk_r_REG646_S3 ( .D(n236), .CP(clk), .SN(n29649), .Q(n17513) );
  HS65_LH_DFPSQX9 clk_r_REG865_S3 ( .D(n13646), .CP(clk), .SN(n29646), .Q(
        n17644) );
  HS65_LH_DFPSQX9 clk_r_REG616_S1 ( .D(n17201), .CP(clk), .SN(n41000), .Q(
        n17375) );
  HS65_LH_DFPSQX9 clk_r_REG598_S1 ( .D(n17202), .CP(clk), .SN(n29645), .Q(
        n17304) );
  HS65_LH_DFPSQX9 clk_r_REG620_S1 ( .D(n15732), .CP(clk), .SN(n29646), .Q(
        n17443) );
  HS65_LH_DFPSQX9 clk_r_REG875_S3 ( .D(n15740), .CP(clk), .SN(n29650), .Q(
        n17442) );
  HS65_LH_DFPSQX9 clk_r_REG658_S3 ( .D(n251), .CP(clk), .SN(n29652), .Q(n17295) );
  HS65_LH_DFPSQX9 clk_r_REG892_S3 ( .D(n15474), .CP(clk), .SN(n41000), .Q(
        n17576) );
  HS65_LH_DFPSQX9 clk_r_REG866_S3 ( .D(n17208), .CP(clk), .SN(n29652), .Q(
        n17433) );
  HS65_LH_BFX35 U4230 ( .A(n17447), .Z(n29596) );
  HS65_LH_BFX35 U4334 ( .A(n18155), .Z(n29597) );
  HS65_LH_BFX35 U4337 ( .A(n17460), .Z(n29598) );
  HS65_LH_BFX35 U4438 ( .A(n18136), .Z(n29599) );
  HS65_LH_BFX35 U4441 ( .A(n17461), .Z(n29600) );
  HS65_LH_AOI21X2 U4542 ( .A(n38566), .B(n33214), .C(n33067), .Z(n15426) );
  HS65_LH_NAND2X2 U4545 ( .A(n16037), .B(n16036), .Z(n29538) );
  HS65_LH_NAND2X2 U4646 ( .A(n16894), .B(n16893), .Z(n16902) );
  HS65_LH_NAND4ABX3 U4649 ( .A(n16798), .B(n16797), .C(n16796), .D(n16795), 
        .Z(n16801) );
  HS65_LH_NAND2X2 U4753 ( .A(n16794), .B(n16793), .Z(n16802) );
  HS65_LH_AOI22X1 U4854 ( .A(n17417), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][22] ), .C(n36561), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][22] ), .Z(n16232)
         );
  HS65_LH_NAND2X2 U4958 ( .A(n16814), .B(n16813), .Z(n16822) );
  HS65_LH_NAND2X2 U4961 ( .A(n17059), .B(n17058), .Z(n17070) );
  HS65_LH_BFX2 U5383 ( .A(n18122), .Z(n18348) );
  HS65_LH_BFX2 U6156 ( .A(n27626), .Z(n19087) );
  HS65_LH_BFX2 U6157 ( .A(n17584), .Z(n19088) );
  HS65_LH_BFX2 U6158 ( .A(n19088), .Z(n19089) );
  HS65_LH_BFX2 U6159 ( .A(n19089), .Z(n19090) );
  HS65_LH_NAND4ABX3 U6163 ( .A(n16518), .B(n16517), .C(n16516), .D(n16515), 
        .Z(n16521) );
  HS65_LH_NAND4ABX3 U7082 ( .A(n16312), .B(n16311), .C(n16310), .D(n16309), 
        .Z(n16315) );
  HS65_LH_NAND4ABX3 U7091 ( .A(n16301), .B(n16300), .C(n16299), .D(n16298), 
        .Z(n16304) );
  HS65_LH_NAND4ABX3 U7691 ( .A(n16241), .B(n16240), .C(n16239), .D(n16238), 
        .Z(n16244) );
  HS65_LH_IVX2 U8219 ( .A(n17423), .Z(n20341) );
  HS65_LH_IVX2 U8221 ( .A(n20341), .Z(n20342) );
  HS65_LH_BFX2 U8427 ( .A(n35786), .Z(n20433) );
  HS65_LH_NAND4ABX3 U8491 ( .A(n16323), .B(n16322), .C(n16321), .D(n16320), 
        .Z(n16327) );
  HS65_LH_BFX2 U9499 ( .A(n17420), .Z(n20916) );
  HS65_LH_NAND4ABX3 U9983 ( .A(n17162), .B(n17161), .C(n17160), .D(n17159), 
        .Z(n17169) );
  HS65_LH_BFX2 U9985 ( .A(n29426), .Z(n21117) );
  HS65_LH_NAND2X2 U11931 ( .A(n16654), .B(n16653), .Z(n16662) );
  HS65_LH_BFX2 U11943 ( .A(n17396), .Z(n21638) );
  HS65_LH_IVX2 U12054 ( .A(n33653), .Z(n21749) );
  HS65_LH_BFX2 U12767 ( .A(n19090), .Z(n21994) );
  HS65_LH_BFX2 U12781 ( .A(n21994), .Z(n22001) );
  HS65_LH_BFX2 U12816 ( .A(n22001), .Z(n22006) );
  HS65_LH_NAND4ABX3 U19258 ( .A(n16752), .B(n16751), .C(n16750), .D(n16749), 
        .Z(n1588) );
  HS65_LH_NAND4ABX3 U19390 ( .A(n15955), .B(n15954), .C(n15953), .D(n15952), 
        .Z(n2502) );
  HS65_LH_IVX2 U20459 ( .A(n15491), .Z(n24656) );
  HS65_LH_AOI21X2 U20581 ( .A(n32748), .B(n14661), .C(n14660), .Z(n14693) );
  HS65_LH_IVX2 U21655 ( .A(n26258), .Z(n25850) );
  HS65_LH_IVX2 U21656 ( .A(n25850), .Z(n25851) );
  HS65_LH_IVX2 U21728 ( .A(n15718), .Z(n25922) );
  HS65_LH_IVX2 U22046 ( .A(n39522), .Z(n26240) );
  HS65_LH_IVX2 U22047 ( .A(n26240), .Z(n26241) );
  HS65_LH_IVX2 U22063 ( .A(n27019), .Z(n26257) );
  HS65_LH_IVX2 U22064 ( .A(n26257), .Z(n26258) );
  HS65_LH_IVX2 U22382 ( .A(n33749), .Z(n26577) );
  HS65_LH_IVX2 U22564 ( .A(n33785), .Z(n26759) );
  HS65_LH_BFX2 U22821 ( .A(n27066), .Z(n27019) );
  HS65_LH_BFX2 U22868 ( .A(n27100), .Z(n27066) );
  HS65_LH_BFX2 U22902 ( .A(n39496), .Z(n27100) );
  HS65_LH_NAND4ABX3 U23230 ( .A(n16792), .B(n16791), .C(n16790), .D(n16789), 
        .Z(n1542) );
  HS65_LH_BFX2 U23244 ( .A(n22006), .Z(n27442) );
  HS65_LH_BFX2 U23264 ( .A(n27442), .Z(n27462) );
  HS65_LH_BFX2 U23283 ( .A(n27462), .Z(n27481) );
  HS65_LH_BFX2 U23300 ( .A(n27481), .Z(n27498) );
  HS65_LH_BFX2 U23318 ( .A(n27498), .Z(n27516) );
  HS65_LH_BFX2 U23336 ( .A(n27516), .Z(n27534) );
  HS65_LH_BFX2 U23357 ( .A(n27534), .Z(n27555) );
  HS65_LH_BFX2 U23375 ( .A(n27555), .Z(n27573) );
  HS65_LH_BFX2 U23393 ( .A(n27573), .Z(n27591) );
  HS65_LH_BFX2 U23411 ( .A(n27591), .Z(n27609) );
  HS65_LH_BFX2 U23428 ( .A(n27639), .Z(n27626) );
  HS65_LH_BFX2 U23441 ( .A(n27652), .Z(n27639) );
  HS65_LH_BFX2 U23454 ( .A(n27665), .Z(n27652) );
  HS65_LH_BFX2 U23467 ( .A(n27609), .Z(n27665) );
  HS65_LH_BFX2 U23589 ( .A(n27790), .Z(n27787) );
  HS65_LH_BFX2 U23592 ( .A(n39488), .Z(n27790) );
  HS65_LH_NAND4ABX3 U24692 ( .A(n16592), .B(n16591), .C(n16590), .D(n16589), 
        .Z(n1772) );
  HS65_LH_NAND4ABX3 U24935 ( .A(n16978), .B(n16977), .C(n16976), .D(n16975), 
        .Z(n16981) );
  HS65_LH_BFX2 U25233 ( .A(n29434), .Z(n29426) );
  HS65_LH_BFX2 U25241 ( .A(n29440), .Z(n29434) );
  HS65_LH_BFX2 U25247 ( .A(n29443), .Z(n29440) );
  HS65_LH_IVX2 U25249 ( .A(n29451), .Z(n29442) );
  HS65_LH_IVX2 U25250 ( .A(n29442), .Z(n29443) );
  HS65_LH_IVX2 U25258 ( .A(n40905), .Z(n29451) );
  HS65_LH_CNIVX3 U25361 ( .A(n9508), .Z(n17214) );
  HS65_LH_IVX2 U25362 ( .A(n29694), .Z(n29647) );
  HS65_LH_IVX2 U25363 ( .A(n29694), .Z(n29697) );
  HS65_LH_NOR2X2 U25364 ( .A(n6651), .B(n15069), .Z(n15075) );
  HS65_LH_IVX2 U25365 ( .A(n29694), .Z(n29648) );
  HS65_LH_IVX4 U25368 ( .A(n29694), .Z(n29649) );
  HS65_LH_AOI22X1 U25369 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][27] ), .B(n17120), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][27] ), .D(
        n17398), .Z(n29534) );
  HS65_LH_AOI22X1 U25370 ( .A(n36264), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][26] ), .C(n29603), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][26] ), .Z(
        n29535) );
  HS65_LH_AOI22X1 U25371 ( .A(n16406), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][30] ), .C(n17423), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[15][30] ), .Z(
        n29536) );
  HS65_LH_AOI21X2 U25374 ( .A(n17567), .B(n17305), .C(n17573), .Z(n29540) );
  HS65_LH_NAND2X2 U25375 ( .A(n16067), .B(n16066), .Z(n16075) );
  HS65_LH_OAI21X2 U25376 ( .A(n14894), .B(n15218), .C(n14893), .Z(n14903) );
  HS65_LH_NAND2X2 U25377 ( .A(n29635), .B(n40560), .Z(n15392) );
  HS65_LH_NAND4ABX3 U25378 ( .A(n16427), .B(n16426), .C(n16425), .D(n16424), 
        .Z(n1974) );
  HS65_LH_BFX2 U25379 ( .A(n18125), .Z(n29542) );
  HS65_LH_NAND4ABX3 U25380 ( .A(n15895), .B(n15894), .C(n15893), .D(n15892), 
        .Z(n2574) );
  HS65_LH_BFX2 U25381 ( .A(n17430), .Z(n29543) );
  HS65_LH_BFX2 U25385 ( .A(n17414), .Z(n29547) );
  HS65_LH_NAND2X2 U25386 ( .A(n16157), .B(n16156), .Z(n16165) );
  HS65_LH_IVX2 U25387 ( .A(n36264), .Z(n29548) );
  HS65_LH_IVX2 U25388 ( .A(n29548), .Z(n29549) );
  HS65_LH_NAND4ABX3 U25389 ( .A(n16115), .B(n16114), .C(n16113), .D(n16112), 
        .Z(n2310) );
  HS65_LH_NAND2X2 U25390 ( .A(n16097), .B(n16096), .Z(n16105) );
  HS65_LH_NAND2X2 U25392 ( .A(n35802), .B(n15906), .Z(n15915) );
  HS65_LH_BFX2 U25393 ( .A(n17426), .Z(n29551) );
  HS65_LH_BFX2 U25394 ( .A(n17418), .Z(n29552) );
  HS65_LH_NAND4ABX3 U25395 ( .A(n16225), .B(n16224), .C(n36423), .D(n16222), 
        .Z(n2165) );
  HS65_LH_BFX2 U25396 ( .A(n17411), .Z(n29553) );
  HS65_LH_NAND2X2 U25397 ( .A(n15977), .B(n15976), .Z(n15985) );
  HS65_LH_AOI22X1 U25398 ( .A(n17425), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][18] ), .C(n29561), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][18] ), .Z(n16139) );
  HS65_LH_NAND2X2 U25399 ( .A(n16147), .B(n16146), .Z(n16155) );
  HS65_LH_BFX2 U25400 ( .A(n35698), .Z(n29554) );
  HS65_LH_NAND2X2 U25401 ( .A(n15765), .B(n15764), .Z(n15777) );
  HS65_LH_NAND4ABX3 U25406 ( .A(n15935), .B(n36695), .C(n36698), .D(n15932), 
        .Z(n2526) );
  HS65_LH_NAND2X2 U25407 ( .A(n15917), .B(n15916), .Z(n15925) );
  HS65_LH_OA222X4 U25408 ( .A(n17611), .B(n17843), .C(n17631), .D(
        \u_DataPath/dataOut_exe_i [31]), .E(n17476), .F(n17363), .Z(n29559) );
  HS65_LH_BFX2 U25409 ( .A(n36571), .Z(n29560) );
  HS65_LH_BFX2 U25410 ( .A(n17424), .Z(n29561) );
  HS65_LH_BFX35 U25411 ( .A(n17486), .Z(n29562) );
  HS65_LH_BFX35 U25412 ( .A(n17485), .Z(n29563) );
  HS65_LH_BFX35 U25413 ( .A(n17487), .Z(n29564) );
  HS65_LH_BFX35 U25414 ( .A(n17488), .Z(n29565) );
  HS65_LH_BFX35 U25415 ( .A(n18152), .Z(n29566) );
  HS65_LH_BFX35 U25416 ( .A(n18154), .Z(n29567) );
  HS65_LH_BFX35 U25417 ( .A(n18151), .Z(n29568) );
  HS65_LH_BFX35 U25418 ( .A(n17520), .Z(n29569) );
  HS65_LH_BFX35 U25419 ( .A(n18153), .Z(n29570) );
  HS65_LH_BFX35 U25420 ( .A(n18150), .Z(n29571) );
  HS65_LH_BFX35 U25421 ( .A(n18137), .Z(n29572) );
  HS65_LH_BFX35 U25422 ( .A(n18147), .Z(n29573) );
  HS65_LH_BFX35 U25423 ( .A(n18149), .Z(n29574) );
  HS65_LH_BFX35 U25424 ( .A(n18148), .Z(n29575) );
  HS65_LH_BFX35 U25425 ( .A(n17483), .Z(n29576) );
  HS65_LH_BFX35 U25426 ( .A(n17522), .Z(n29577) );
  HS65_LH_BFX35 U25427 ( .A(n17521), .Z(n29578) );
  HS65_LH_BFX35 U25428 ( .A(n17519), .Z(n29579) );
  HS65_LH_BFX35 U25429 ( .A(n17455), .Z(n29580) );
  HS65_LH_BFX35 U25430 ( .A(n17456), .Z(n29581) );
  HS65_LH_BFX35 U25431 ( .A(n17457), .Z(n29582) );
  HS65_LH_BFX35 U25432 ( .A(n17458), .Z(n29583) );
  HS65_LH_BFX35 U25433 ( .A(n17484), .Z(n29584) );
  HS65_LH_BFX35 U25434 ( .A(n18139), .Z(n29585) );
  HS65_LH_BFX35 U25435 ( .A(n18138), .Z(n29586) );
  HS65_LH_BFX35 U25436 ( .A(n18127), .Z(n29587) );
  HS65_LH_BFX35 U25437 ( .A(n17453), .Z(n29588) );
  HS65_LH_BFX35 U25438 ( .A(n17510), .Z(n29589) );
  HS65_LH_BFX35 U25439 ( .A(n17491), .Z(n29590) );
  HS65_LH_BFX35 U25440 ( .A(n17452), .Z(n29591) );
  HS65_LH_BFX35 U25441 ( .A(n17451), .Z(n29592) );
  HS65_LH_NAND4ABX3 U25443 ( .A(n16902), .B(n16901), .C(n16900), .D(n16899), 
        .Z(n1403) );
  HS65_LH_BFX2 U25446 ( .A(n18123), .Z(n29602) );
  HS65_LH_NAND2X2 U25447 ( .A(n15877), .B(n15876), .Z(n15885) );
  HS65_LH_NAND2X2 U25448 ( .A(n16247), .B(n16246), .Z(n16255) );
  HS65_LH_BFX2 U25449 ( .A(n17431), .Z(n29603) );
  HS65_LH_BFX2 U25450 ( .A(n17422), .Z(n29604) );
  HS65_LH_NAND2X2 U25451 ( .A(n16047), .B(n16046), .Z(n16055) );
  HS65_LH_NAND2X2 U25452 ( .A(n16381), .B(n16380), .Z(n16391) );
  HS65_LH_NAND2X2 U25453 ( .A(n16107), .B(n16106), .Z(n16115) );
  HS65_LH_IVX2 U25454 ( .A(n36759), .Z(n29605) );
  HS65_LH_IVX2 U25455 ( .A(n29605), .Z(n29606) );
  HS65_LH_NAND2X2 U25456 ( .A(n15897), .B(n15896), .Z(n15905) );
  HS65_LH_IVX2 U25459 ( .A(n17407), .Z(n29609) );
  HS65_LH_IVX2 U25460 ( .A(n29609), .Z(n29610) );
  HS65_LH_AOI22X1 U25465 ( .A(n18123), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][11] ), .C(n40994), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[19][11] ), .Z(n16013)
         );
  HS65_LH_IVX2 U25466 ( .A(n17406), .Z(n29615) );
  HS65_LH_IVX2 U25467 ( .A(n29615), .Z(n29616) );
  HS65_LH_IVX2 U25468 ( .A(n17405), .Z(n29617) );
  HS65_LH_IVX2 U25469 ( .A(n29617), .Z(n29618) );
  HS65_LH_NAND2X2 U25470 ( .A(n15797), .B(n15796), .Z(n15805) );
  HS65_LH_IVX2 U25471 ( .A(n17427), .Z(n29619) );
  HS65_LH_IVX2 U25472 ( .A(n29619), .Z(n29620) );
  HS65_LH_NAND4ABX3 U25474 ( .A(n16612), .B(n16611), .C(n16610), .D(n16609), 
        .Z(n1749) );
  HS65_LH_NAND2X2 U25475 ( .A(n16594), .B(n16593), .Z(n16602) );
  HS65_LH_NAND4ABX3 U25476 ( .A(n16692), .B(n16691), .C(n16690), .D(n16689), 
        .Z(n1657) );
  HS65_LH_BFX2 U25477 ( .A(n17412), .Z(n29622) );
  HS65_LH_NAND4ABX3 U25478 ( .A(n16812), .B(n16811), .C(n16810), .D(n16809), 
        .Z(n1519) );
  HS65_LH_BFX2 U25479 ( .A(n17404), .Z(n29623) );
  HS65_LH_BFX2 U25480 ( .A(n15422), .Z(n29624) );
  HS65_LH_IVX2 U25491 ( .A(n15394), .Z(n29635) );
  HS65_LH_NAND4ABX3 U25498 ( .A(n16822), .B(n16821), .C(n16820), .D(n16819), 
        .Z(n1495) );
  HS65_LH_IVX2 U25500 ( .A(n29694), .Z(n29643) );
  HS65_LH_IVX2 U25501 ( .A(n29694), .Z(n29644) );
  HS65_LH_IVX4 U25502 ( .A(n29694), .Z(n29645) );
  HS65_LH_IVX4 U25503 ( .A(n29694), .Z(n29646) );
  HS65_LH_IVX4 U25504 ( .A(n29694), .Z(n29652) );
  HS65_LH_CNIVX3 U25505 ( .A(n12489), .Z(n29650) );
  HS65_LH_IVX35 U25506 ( .A(n29653), .Z(n29654) );
  HS65_LH_IVX35 U25507 ( .A(n29655), .Z(n29656) );
  HS65_LH_IVX35 U25508 ( .A(n29657), .Z(n29658) );
  HS65_LH_IVX35 U25509 ( .A(n29659), .Z(n29660) );
  HS65_LH_IVX35 U25510 ( .A(n29661), .Z(n29662) );
  HS65_LH_IVX35 U25511 ( .A(n29663), .Z(n29664) );
  HS65_LH_IVX35 U25512 ( .A(n29665), .Z(n29666) );
  HS65_LH_IVX35 U25513 ( .A(n29667), .Z(n29668) );
  HS65_LH_IVX35 U25514 ( .A(n29669), .Z(n29670) );
  HS65_LH_IVX35 U25515 ( .A(n29671), .Z(n29672) );
  HS65_LH_IVX35 U25516 ( .A(n29673), .Z(n29674) );
  HS65_LH_IVX35 U25517 ( .A(n29675), .Z(n29676) );
  HS65_LH_IVX35 U25518 ( .A(n29677), .Z(n29678) );
  HS65_LH_IVX35 U25519 ( .A(n29679), .Z(n29680) );
  HS65_LH_IVX35 U25520 ( .A(n29681), .Z(n29682) );
  HS65_LH_IVX35 U25521 ( .A(n29683), .Z(n29684) );
  HS65_LH_IVX35 U25522 ( .A(n29685), .Z(n29686) );
  HS65_LH_IVX35 U25523 ( .A(n29687), .Z(n29688) );
  HS65_LH_IVX2 U25524 ( .A(n9508), .Z(n17213) );
  HS65_LH_NAND2X4 U25525 ( .A(n15341), .B(n15500), .Z(n14626) );
  HS65_LH_NOR2X2 U25526 ( .A(n14922), .B(n17474), .Z(n15422) );
  HS65_LH_NOR2X3 U25527 ( .A(n14897), .B(n15344), .Z(n15517) );
  HS65_LH_IVX35 U25528 ( .A(n29689), .Z(n29690) );
  HS65_LH_IVX2 U25529 ( .A(n17527), .Z(n29691) );
  HS65_LH_CNIVX3 U25530 ( .A(n29691), .Z(n29692) );
  HS65_LH_CNIVX3 U25531 ( .A(n29691), .Z(n29693) );
  HS65_LH_IVX4 U25534 ( .A(n29694), .Z(n29698) );
  HS65_LH_OR2X4 U25535 ( .A(n14547), .B(n15344), .Z(n29699) );
  HS65_LH_IVX2 U25536 ( .A(n15707), .Z(n17245) );
  HS65_LH_IVX2 U25537 ( .A(n38579), .Z(n10437) );
  HS65_LH_IVX2 U25538 ( .A(n6651), .Z(n14037) );
  HS65_LH_IVX2 U25539 ( .A(n29699), .Z(n13892) );
  HS65_LH_DFPSQX4 clk_r_REG766_S3 ( .D(n1913), .CP(clk), .SN(n40998), .Q(
        n17625) );
  HS65_LH_DFPSQX4 clk_r_REG905_S3 ( .D(n13639), .CP(clk), .SN(n40997), .Q(
        n17645) );
  HS65_LH_DFPSQX4 clk_r_REG884_S3 ( .D(n10317), .CP(clk), .SN(n41000), .Q(
        n17774) );
  HS65_LH_DFPSQX4 clk_r_REG681_S3 ( .D(n1101), .CP(clk), .SN(n40999), .Q(
        n17572) );
  HS65_LH_DFPSQX4 clk_r_REG668_S3 ( .D(n1103), .CP(clk), .SN(n40998), .Q(
        n17571) );
  HS65_LH_DFPSQX4 clk_r_REG852_S3 ( .D(n15167), .CP(clk), .SN(n40997), .Q(
        n17586) );
  HS65_LH_DFPSQX4 clk_r_REG828_S3 ( .D(n1113), .CP(clk), .SN(n41000), .Q(
        n17575) );
  HS65_LH_DFPSQX4 clk_r_REG651_S3 ( .D(n243), .CP(clk), .SN(n40999), .Q(n17439) );
  HS65_LH_DFPSQX4 clk_r_REG693_S3 ( .D(n277), .CP(clk), .SN(n40998), .Q(n17303) );
  HS65_LH_DFPSQX4 clk_r_REG10_S1 ( .D(n258), .CP(clk), .SN(n40997), .Q(n17632)
         );
  HS65_LH_DFPSQX4 clk_r_REG656_S3 ( .D(n224), .CP(clk), .SN(n41000), .Q(n17299) );
  HS65_LH_DFPSQX4 clk_r_REG11_S1 ( .D(n15753), .CP(clk), .SN(n40999), .Q(
        n17301) );
  HS65_LH_DFPSQX4 clk_r_REG779_S3 ( .D(n16447), .CP(clk), .SN(n40998), .Q(
        n17420) );
  HS65_LH_DFPSQX4 clk_r_REG652_S3 ( .D(n218), .CP(clk), .SN(n40997), .Q(n17374) );
  HS65_LL_DFPHQX27 clk_r_REG260_S1 ( .D(n14100), .E(
        \u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n17637) );
  HS65_LH_DFPQX4 clk_r_REG565_S3 ( .D(n40862), .CP(clk), .Q(n17599) );
  HS65_LH_DFPQX4 clk_r_REG890_S5 ( .D(n40270), .CP(clk), .Q(n17764) );
  HS65_LH_DFPQX4 clk_r_REG889_S5 ( .D(n40293), .CP(clk), .Q(n17766) );
  HS65_LH_DFPQX4 clk_r_REG740_S5 ( .D(n40316), .CP(clk), .Q(n17951) );
  HS65_LH_DFPQX4 clk_r_REG732_S5 ( .D(n40339), .CP(clk), .Q(n17938) );
  HS65_LH_DFPQX4 clk_r_REG724_S5 ( .D(n40385), .CP(clk), .Q(n17912) );
  HS65_LH_DFPQX4 clk_r_REG717_S5 ( .D(n40408), .CP(clk), .Q(n17993) );
  HS65_LH_DFPQX4 clk_r_REG702_S5 ( .D(n40362), .CP(clk), .Q(n17961) );
  HS65_LH_DFPQX4 clk_r_REG913_S1 ( .D(n2733), .CP(clk), .Q(n18159) );
  HS65_LH_DFPQX4 clk_r_REG896_S5 ( .D(\u_DataPath/cw_tomem_i [0]), .CP(clk), 
        .Q(n17561) );
  HS65_LH_DFPQX4 clk_r_REG265_S3 ( .D(\u_DataPath/pc_4_to_ex_i [24]), .CP(clk), 
        .Q(n17543) );
  HS65_LH_DFPQX4 clk_r_REG214_S3 ( .D(\u_DataPath/pc_4_to_ex_i [31]), .CP(clk), 
        .Q(n17550) );
  HS65_LH_DFPQX4 clk_r_REG205_S3 ( .D(\u_DataPath/pc_4_to_ex_i [30]), .CP(clk), 
        .Q(n17549) );
  HS65_LH_DFPQX4 clk_r_REG390_S3 ( .D(\u_DataPath/pc_4_to_ex_i [10]), .CP(clk), 
        .Q(n17529) );
  HS65_LH_DFPQX4 clk_r_REG380_S3 ( .D(\u_DataPath/pc_4_to_ex_i [11]), .CP(clk), 
        .Q(n17530) );
  HS65_LH_DFPQX4 clk_r_REG363_S3 ( .D(\u_DataPath/pc_4_to_ex_i [13]), .CP(clk), 
        .Q(n17532) );
  HS65_LH_DFPQX4 clk_r_REG340_S3 ( .D(\u_DataPath/pc_4_to_ex_i [15]), .CP(clk), 
        .Q(n17534) );
  HS65_LH_DFPQX4 clk_r_REG321_S3 ( .D(\u_DataPath/pc_4_to_ex_i [17]), .CP(clk), 
        .Q(n17536) );
  HS65_LH_DFPQX4 clk_r_REG313_S3 ( .D(\u_DataPath/pc_4_to_ex_i [18]), .CP(clk), 
        .Q(n17537) );
  HS65_LH_DFPQX4 clk_r_REG305_S3 ( .D(\u_DataPath/pc_4_to_ex_i [19]), .CP(clk), 
        .Q(n17538) );
  HS65_LH_DFPQX4 clk_r_REG297_S3 ( .D(\u_DataPath/pc_4_to_ex_i [20]), .CP(clk), 
        .Q(n17539) );
  HS65_LH_DFPQX4 clk_r_REG289_S3 ( .D(\u_DataPath/pc_4_to_ex_i [21]), .CP(clk), 
        .Q(n17540) );
  HS65_LH_DFPQX4 clk_r_REG281_S3 ( .D(\u_DataPath/pc_4_to_ex_i [22]), .CP(clk), 
        .Q(n17541) );
  HS65_LH_DFPQX4 clk_r_REG273_S3 ( .D(\u_DataPath/pc_4_to_ex_i [23]), .CP(clk), 
        .Q(n17542) );
  HS65_LH_DFPQX4 clk_r_REG255_S3 ( .D(\u_DataPath/pc_4_to_ex_i [25]), .CP(clk), 
        .Q(n17544) );
  HS65_LH_DFPQX4 clk_r_REG247_S3 ( .D(\u_DataPath/pc_4_to_ex_i [26]), .CP(clk), 
        .Q(n17545) );
  HS65_LH_DFPQX4 clk_r_REG237_S3 ( .D(\u_DataPath/pc_4_to_ex_i [27]), .CP(clk), 
        .Q(n17546) );
  HS65_LH_DFPQX4 clk_r_REG229_S3 ( .D(\u_DataPath/pc_4_to_ex_i [28]), .CP(clk), 
        .Q(n17547) );
  HS65_LH_DFPQX4 clk_r_REG219_S3 ( .D(\u_DataPath/pc_4_to_ex_i [29]), .CP(clk), 
        .Q(n17548) );
  HS65_LH_DFPQX4 clk_r_REG700_S4 ( .D(\u_DataPath/u_idexreg/N35 ), .CP(clk), 
        .Q(n17556) );
  HS65_LH_DFPQX4 clk_r_REG350_S3 ( .D(\u_DataPath/pc_4_to_ex_i [14]), .CP(clk), 
        .Q(n17533) );
  HS65_LH_DFPQX4 clk_r_REG373_S3 ( .D(\u_DataPath/pc_4_to_ex_i [12]), .CP(clk), 
        .Q(n17531) );
  HS65_LH_DFPQX4 clk_r_REG332_S3 ( .D(\u_DataPath/pc_4_to_ex_i [16]), .CP(clk), 
        .Q(n17535) );
  HS65_LH_DFPQX4 clk_r_REG734_S4 ( .D(\u_DataPath/u_idexreg/N39 ), .CP(clk), 
        .Q(n17560) );
  HS65_LH_DFPQX4 clk_r_REG726_S4 ( .D(\u_DataPath/u_idexreg/N38 ), .CP(clk), 
        .Q(n17559) );
  HS65_LH_DFPQX4 clk_r_REG719_S4 ( .D(\u_DataPath/u_idexreg/N37 ), .CP(clk), 
        .Q(n17558) );
  HS65_LH_DFPQX4 clk_r_REG704_S4 ( .D(\u_DataPath/u_idexreg/N36 ), .CP(clk), 
        .Q(n17557) );
  HS65_LH_DFPQX4 clk_r_REG790_S1 ( .D(\u_DataPath/idex_rt_i [2]), .CP(clk), 
        .Q(n17499) );
  HS65_LH_DFPQX4 clk_r_REG797_S1 ( .D(\u_DataPath/u_idexreg/N44 ), .CP(clk), 
        .Q(n17498) );
  HS65_LH_DFPQX4 clk_r_REG783_S1 ( .D(\u_DataPath/u_idexreg/N42 ), .CP(clk), 
        .Q(n17500) );
  HS65_LH_DFPQX4 clk_r_REG249_S4 ( .D(n38676), .CP(clk), .Q(n17960) );
  HS65_LH_DFPQX4 clk_r_REG686_S4 ( .D(\u_DataPath/u_idexreg/N31 ), .CP(clk), 
        .Q(n17552) );
  HS65_LH_DFPQX4 clk_r_REG306_S3 ( .D(n14380), .CP(clk), .Q(n17597) );
  HS65_LH_DFPQX4 clk_r_REG290_S3 ( .D(n14696), .CP(clk), .Q(n17596) );
  HS65_LH_DFPQX4 clk_r_REG274_S3 ( .D(n14484), .CP(clk), .Q(n17595) );
  HS65_LH_DFPQX4 clk_r_REG256_S3 ( .D(n14749), .CP(clk), .Q(n17594) );
  HS65_LH_DFPQX4 clk_r_REG238_S3 ( .D(n14299), .CP(clk), .Q(n17593) );
  HS65_LH_DFPQX4 clk_r_REG220_S3 ( .D(n14655), .CP(clk), .Q(n17589) );
  HS65_LH_DFPQX4 clk_r_REG314_S3 ( .D(n8924), .CP(clk), .Q(n17872) );
  HS65_LH_DFPQX4 clk_r_REG298_S3 ( .D(n8448), .CP(clk), .Q(n17892) );
  HS65_LH_DFPQX4 clk_r_REG282_S3 ( .D(n8097), .CP(clk), .Q(n17906) );
  HS65_LH_DFPQX4 clk_r_REG248_S3 ( .D(n6788), .CP(clk), .Q(n17963) );
  HS65_LH_DFPQX4 clk_r_REG230_S3 ( .D(n7988), .CP(clk), .Q(n17914) );
  HS65_LH_DFPQX4 clk_r_REG861_S1 ( .D(\u_DataPath/u_idexreg/N56 ), .CP(clk), 
        .Q(n17526) );
  HS65_LH_DFPQX4 clk_r_REG743_S4 ( .D(\u_DataPath/u_idexreg/N40 ), .CP(clk), 
        .Q(n18158) );
  HS65_LH_DFPQX4 clk_r_REG697_S4 ( .D(\u_DataPath/u_idexreg/N34 ), .CP(clk), 
        .Q(n17555) );
  HS65_LH_DFPQX4 clk_r_REG694_S4 ( .D(\u_DataPath/u_idexreg/N33 ), .CP(clk), 
        .Q(n17554) );
  HS65_LH_DFPQX4 clk_r_REG690_S4 ( .D(\u_DataPath/u_idexreg/N32 ), .CP(clk), 
        .Q(n17553) );
  HS65_LH_DFPQX4 clk_r_REG322_S3 ( .D(n15052), .CP(clk), .Q(n17598) );
  HS65_LH_DFPQX4 clk_r_REG909_S1 ( .D(\u_DataPath/idex_rt_i [0]), .CP(clk), 
        .Q(n17492) );
  HS65_LH_DFPQX4 clk_r_REG804_S1 ( .D(\u_DataPath/idex_rt_i [4]), .CP(clk), 
        .Q(n17497) );
  HS65_LH_DFPQX4 clk_r_REG351_S3 ( .D(n6189), .CP(clk), .Q(n17986) );
  HS65_LH_DFPQX4 clk_r_REG391_S3 ( .D(n6703), .CP(clk), .Q(n17967) );
  HS65_LH_DFPQX4 clk_r_REG737_S1 ( .D(n1907), .CP(clk), .Q(n17518) );
  HS65_LH_DFPQX4 clk_r_REG593_S4 ( .D(n9538), .CP(clk), .Q(n17844) );
  HS65_LH_DFPQX4 clk_r_REG863_S1 ( .D(n5507), .CP(clk), .Q(n18000) );
  HS65_LH_DFPQX4 clk_r_REG239_S4 ( .D(n40452), .CP(clk), .Q(n17992) );
  HS65_LH_DFPQX4 clk_r_REG862_S1 ( .D(n5234), .CP(clk), .Q(n18002) );
  HS65_LH_DFPQX4 clk_r_REG910_S1 ( .D(n14115), .CP(clk), .Q(n17624) );
  HS65_LH_DFPQX4 clk_r_REG805_S1 ( .D(n14118), .CP(clk), .Q(n17621) );
  HS65_LH_DFPQX4 clk_r_REG746_S1 ( .D(n14124), .CP(clk), .Q(n17507) );
  HS65_LH_DFPQX4 clk_r_REG0_S1 ( .D(\u_DataPath/u_idexreg/N29 ), .CP(clk), .Q(
        n17551) );
  HS65_LH_DFPQX4 clk_r_REG853_S1 ( .D(\u_DataPath/rs_ex_i [2]), .CP(clk), .Q(
        n17494) );
  HS65_LH_DFPQX4 clk_r_REG846_S1 ( .D(\u_DataPath/rs_ex_i [0]), .CP(clk), .Q(
        n17496) );
  HS65_LH_DFPQX4 clk_r_REG857_S1 ( .D(\u_DataPath/rs_ex_i [3]), .CP(clk), .Q(
        n17493) );
  HS65_LH_DFPQX4 clk_r_REG849_S1 ( .D(\u_DataPath/rs_ex_i [1]), .CP(clk), .Q(
        n17495) );
  HS65_LH_DFPQX4 clk_r_REG738_S1 ( .D(n1106), .CP(clk), .Q(n17619) );
  HS65_LH_DFPQX4 clk_r_REG661_S1 ( .D(n15641), .CP(clk), .Q(n17609) );
  HS65_LH_DFPQX4 clk_r_REG528_S7 ( .D(n38566), .CP(clk), .Q(n17463) );
  HS65_LH_DFPQX4 clk_r_REG798_S1 ( .D(n13531), .CP(clk), .Q(n17651) );
  HS65_LH_DFPQX4 clk_r_REG682_S1 ( .D(\u_DataPath/u_idexreg/N30 ), .CP(clk), 
        .Q(n17501) );
  HS65_LH_DFPQX4 clk_r_REG664_S1 ( .D(\u_DataPath/u_idexreg/N26 ), .CP(clk), 
        .Q(n17504) );
  HS65_LH_DFPQX4 clk_r_REG675_S1 ( .D(\u_DataPath/u_idexreg/N28 ), .CP(clk), 
        .Q(n17502) );
  HS65_LH_DFPQX4 clk_r_REG670_S1 ( .D(\u_DataPath/u_idexreg/N27 ), .CP(clk), 
        .Q(n17503) );
  HS65_LH_DFPQX4 clk_r_REG747_S1 ( .D(n17211), .CP(clk), .Q(n17628) );
  HS65_LH_DFPQX4 clk_r_REG539_S6 ( .D(n40544), .CP(clk), .Q(n17464) );
  HS65_LH_DFPQX4 clk_r_REG712_S1 ( .D(n110), .CP(clk), .Q(n17319) );
  HS65_LH_DFPQX4 clk_r_REG722_S1 ( .D(n15714), .CP(clk), .Q(n17508) );
  HS65_LH_DFPQX4 clk_r_REG707_S1 ( .D(n15711), .CP(clk), .Q(n17506) );
  HS65_LH_DFPQX4 clk_r_REG715_S1 ( .D(n105), .CP(clk), .Q(n17324) );
  HS65_LH_DFPQX4 clk_r_REG540_S6 ( .D(n14540), .CP(clk), .Q(n17588) );
  HS65_LH_DFPQX4 clk_r_REG231_S4 ( .D(n40581), .CP(clk), .Q(n17911) );
  HS65_LH_DFPQX4 clk_r_REG608_S3 ( .D(n1040), .CP(clk), .Q(n17525) );
  HS65_LH_DFPQX4 clk_r_REG729_S1 ( .D(n15670), .CP(clk), .Q(n17480) );
  HS65_LH_DFPQX4 clk_r_REG784_S1 ( .D(n13537), .CP(clk), .Q(n17650) );
  HS65_LH_DFPQX4 clk_r_REG710_S1 ( .D(n114), .CP(clk), .Q(n17321) );
  HS65_LH_DFPQX4 clk_r_REG714_S1 ( .D(n108), .CP(clk), .Q(n17323) );
  HS65_LH_DFPQX4 clk_r_REG713_S1 ( .D(n112), .CP(clk), .Q(n17322) );
  HS65_LH_DFPQX4 clk_r_REG711_S1 ( .D(n109), .CP(clk), .Q(n17325) );
  HS65_LH_DFPQX4 clk_r_REG221_S4 ( .D(n40630), .CP(clk), .Q(n17937) );
  HS65_LH_DFPQX4 clk_r_REG785_S1 ( .D(n14117), .CP(clk), .Q(n17622) );
  HS65_LH_DFPQX4 clk_r_REG606_S3 ( .D(n1067), .CP(clk), .Q(n17327) );
  HS65_LH_DFPQX4 clk_r_REG708_S1 ( .D(n111), .CP(clk), .Q(n17306) );
  HS65_LH_DFPQX4 clk_r_REG730_S1 ( .D(n15669), .CP(clk), .Q(n17613) );
  HS65_LH_DFPQX4 clk_r_REG709_S1 ( .D(n107), .CP(clk), .Q(n17320) );
  HS65_LH_DFPQX4 clk_r_REG207_S4 ( .D(n40840), .CP(clk), .Q(n17953) );
  HS65_LH_DFPQX4 clk_r_REG594_S4 ( .D(n102), .CP(clk), .Q(n17279) );
  HS65_LH_DFPQX4 clk_r_REG527_S11 ( .D(\u_DataPath/data_read_ex_1_i [31]), 
        .CP(clk), .Q(n17363) );
  HS65_LH_DFPQX4 clk_r_REG522_S11 ( .D(\u_DataPath/data_read_ex_1_i [1]), .CP(
        clk), .Q(n17356) );
  HS65_LH_DFPQX4 clk_r_REG479_S2 ( .D(\u_DataPath/data_read_ex_1_i [3]), .CP(
        clk), .Q(n17358) );
  HS65_LH_DFPQX4 clk_r_REG195_S2 ( .D(\u_DataPath/data_read_ex_1_i [2]), .CP(
        clk), .Q(n17357) );
  HS65_LH_DFPQX4 clk_r_REG133_S2 ( .D(\u_DataPath/data_read_ex_1_i [29]), .CP(
        clk), .Q(n17361) );
  HS65_LH_DFPQX4 clk_r_REG40_S2 ( .D(\u_DataPath/data_read_ex_1_i [30]), .CP(
        clk), .Q(n17362) );
  HS65_LH_DFPQX4 clk_r_REG36_S2 ( .D(\u_DataPath/data_read_ex_1_i [26]), .CP(
        clk), .Q(n17360) );
  HS65_LH_DFPQX4 clk_r_REG7_S2 ( .D(\u_DataPath/data_read_ex_1_i [20]), .CP(
        clk), .Q(n17359) );
  HS65_LH_DFPQX4 clk_r_REG488_S2 ( .D(n8219), .CP(clk), .Q(n17903) );
  HS65_LH_DFPQX4 clk_r_REG189_S2 ( .D(n5901), .CP(clk), .Q(n17997) );
  HS65_LH_DFPQX4 clk_r_REG179_S2 ( .D(n4804), .CP(clk), .Q(n18010) );
  HS65_LH_DFPQX4 clk_r_REG144_S2 ( .D(n5769), .CP(clk), .Q(n17998) );
  HS65_LH_DFPQX4 clk_r_REG128_S2 ( .D(n4935), .CP(clk), .Q(n18008) );
  HS65_LH_DFPQX4 clk_r_REG124_S2 ( .D(n5175), .CP(clk), .Q(n18003) );
  HS65_LH_DFPQX4 clk_r_REG118_S2 ( .D(n4868), .CP(clk), .Q(n18009) );
  HS65_LH_DFPQX4 clk_r_REG103_S2 ( .D(n5571), .CP(clk), .Q(n17999) );
  HS65_LH_DFPQX4 clk_r_REG31_S2 ( .D(n5067), .CP(clk), .Q(n18006) );
  HS65_LH_DFPQX4 clk_r_REG154_S2 ( .D(n4610), .CP(clk), .Q(n18012) );
  HS65_LH_DFPQX4 clk_r_REG85_S2 ( .D(n5133), .CP(clk), .Q(n18004) );
  HS65_LH_DFPQX4 clk_r_REG26_S2 ( .D(n4477), .CP(clk), .Q(n18014) );
  HS65_LH_DFPQX4 clk_r_REG20_S2 ( .D(n4543), .CP(clk), .Q(n18013) );
  HS65_LH_DFPQX4 clk_r_REG607_S3 ( .D(n1059), .CP(clk), .Q(n18157) );
  HS65_LH_DFPHQX4 clk_r_REG426_S1 ( .D(n2871), .E(\u_DataPath/u_fetch/pc1/N3 ), 
        .CP(clk), .Q(n18086) );
  HS65_LH_DFPSQX4 clk_r_REG868_S1 ( .D(n226), .CP(clk), .SN(n29650), .Q(n17297) );
  HS65_LH_DFPSQX4 clk_r_REG659_S3 ( .D(n239), .CP(clk), .SN(n41000), .Q(n17570) );
  HS65_LH_DFPSQX4 clk_r_REG860_S3 ( .D(n15170), .CP(clk), .SN(n29650), .Q(
        n17583) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N122 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][29] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(
        \u_DataPath/u_decode_unit/reg_file0/N108 ), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][15] ) );
  HS65_LH_DFPHQX4 clk_r_REG243_S1 ( .D(n4004), .E(\u_DataPath/u_fetch/pc1/N3 ), 
        .CP(clk), .Q(n18034) );
  HS65_LH_DFPHQX4 clk_r_REG202_S1 ( .D(n15462), .E(\u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n17481) );
  HS65_LH_DFPSQX4 clk_r_REG615_S1 ( .D(n17203), .CP(clk), .SN(n29643), .Q(
        n17302) );
  HS65_LL_CNBFX14 U3521 ( .A(n17450), .Z(n29593) );
  HS65_LL_CNBFX14 U3542 ( .A(n17449), .Z(n29594) );
  HS65_LL_CNBFX14 U3546 ( .A(n17448), .Z(n29595) );
  HS65_LH_NAND4ABX3 U4750 ( .A(n16281), .B(n16280), .C(n16279), .D(n16278), 
        .Z(n16284) );
  HS65_LHS_XNOR2X3 U4857 ( .A(n17550), .B(n15388), .Z(n15389) );
  HS65_LH_NAND2X2 U5069 ( .A(n16574), .B(n16573), .Z(n16582) );
  HS65_LH_IVX2 U5173 ( .A(n18126), .Z(n36570) );
  HS65_LH_IVX2 U5175 ( .A(n17416), .Z(n36758) );
  HS65_LH_IVX2 U5177 ( .A(n17413), .Z(n36560) );
  HS65_LH_BFX9 U5178 ( .A(n17425), .Z(n35786) );
  HS65_LH_IVX2 U5179 ( .A(n17428), .Z(n36384) );
  HS65_LH_BFX9 U5180 ( .A(n17429), .Z(n36045) );
  HS65_LH_BFX9 U5181 ( .A(n17432), .Z(n36264) );
  HS65_LHS_XNOR2X3 U5182 ( .A(n18120), .B(n14108), .Z(n14109) );
  HS65_LH_NOR2X6 U5183 ( .A(n17634), .B(n15465), .Z(n15464) );
  HS65_LH_NAND3X2 U5184 ( .A(n34000), .B(n17305), .C(n17577), .Z(n40985) );
  HS65_LH_BFX9 U5185 ( .A(n17600), .Z(n32748) );
  HS65_LH_NAND2X7 U5186 ( .A(\u_DataPath/takeBranch_out_i ), .B(n17561), .Z(
        n15476) );
  HS65_LH_IVX9 U5187 ( .A(n29694), .Z(n18160) );
  HS65_LH_BFX2 U5188 ( .A(n29701), .Z(n29700) );
  HS65_LH_BFX2 U5189 ( .A(n33259), .Z(n29701) );
  HS65_LH_BFX2 U5190 ( .A(n38701), .Z(n29702) );
  HS65_LH_BFX2 U5191 ( .A(n18092), .Z(n29703) );
  HS65_LH_BFX2 U5192 ( .A(n18091), .Z(n29704) );
  HS65_LH_BFX2 U5194 ( .A(n29706), .Z(n29705) );
  HS65_LH_BFX2 U5196 ( .A(n29707), .Z(n29706) );
  HS65_LH_BFX2 U5198 ( .A(n29708), .Z(n29707) );
  HS65_LH_BFX2 U5200 ( .A(n29709), .Z(n29708) );
  HS65_LH_BFX2 U5202 ( .A(n29710), .Z(n29709) );
  HS65_LH_BFX2 U5204 ( .A(n29711), .Z(n29710) );
  HS65_LH_BFX2 U5206 ( .A(n29712), .Z(n29711) );
  HS65_LH_BFX2 U5208 ( .A(n29713), .Z(n29712) );
  HS65_LH_BFX2 U5210 ( .A(n29714), .Z(n29713) );
  HS65_LH_BFX2 U5212 ( .A(n29715), .Z(n29714) );
  HS65_LH_BFX2 U5215 ( .A(n29716), .Z(n29715) );
  HS65_LH_BFX2 U5216 ( .A(n29717), .Z(n29716) );
  HS65_LH_BFX2 U5217 ( .A(n29718), .Z(n29717) );
  HS65_LH_BFX2 U5218 ( .A(n29719), .Z(n29718) );
  HS65_LH_BFX2 U5219 ( .A(n29720), .Z(n29719) );
  HS65_LH_BFX2 U5220 ( .A(n29721), .Z(n29720) );
  HS65_LH_BFX2 U5221 ( .A(n34387), .Z(n29721) );
  HS65_LH_BFX2 U5222 ( .A(n29723), .Z(n29722) );
  HS65_LH_BFX2 U5223 ( .A(n29724), .Z(n29723) );
  HS65_LH_BFX2 U5224 ( .A(n29725), .Z(n29724) );
  HS65_LH_BFX2 U5225 ( .A(n29726), .Z(n29725) );
  HS65_LH_BFX2 U5226 ( .A(n29727), .Z(n29726) );
  HS65_LH_BFX2 U5227 ( .A(n29728), .Z(n29727) );
  HS65_LH_BFX2 U5228 ( .A(n29729), .Z(n29728) );
  HS65_LH_BFX2 U5229 ( .A(n29730), .Z(n29729) );
  HS65_LH_BFX2 U5230 ( .A(n29731), .Z(n29730) );
  HS65_LH_BFX2 U5231 ( .A(n29732), .Z(n29731) );
  HS65_LH_BFX2 U5232 ( .A(n29733), .Z(n29732) );
  HS65_LH_BFX2 U5233 ( .A(n29734), .Z(n29733) );
  HS65_LH_BFX2 U5234 ( .A(n29735), .Z(n29734) );
  HS65_LH_BFX2 U5235 ( .A(n29736), .Z(n29735) );
  HS65_LH_BFX2 U5236 ( .A(n29737), .Z(n29736) );
  HS65_LH_BFX2 U5237 ( .A(n29738), .Z(n29737) );
  HS65_LH_BFX2 U5238 ( .A(n29739), .Z(n29738) );
  HS65_LH_BFX2 U5239 ( .A(n29740), .Z(n29739) );
  HS65_LH_BFX2 U5240 ( .A(n29741), .Z(n29740) );
  HS65_LH_BFX2 U5241 ( .A(n29742), .Z(n29741) );
  HS65_LH_BFX2 U5242 ( .A(n29743), .Z(n29742) );
  HS65_LH_BFX2 U5243 ( .A(n17733), .Z(n29743) );
  HS65_LH_BFX2 U5244 ( .A(n29745), .Z(n29744) );
  HS65_LH_BFX2 U5245 ( .A(n29746), .Z(n29745) );
  HS65_LH_BFX2 U5246 ( .A(n29747), .Z(n29746) );
  HS65_LH_BFX2 U5247 ( .A(n29748), .Z(n29747) );
  HS65_LH_BFX2 U5248 ( .A(n29749), .Z(n29748) );
  HS65_LH_BFX2 U5249 ( .A(n29750), .Z(n29749) );
  HS65_LH_BFX2 U5250 ( .A(n29751), .Z(n29750) );
  HS65_LH_BFX2 U5251 ( .A(n29752), .Z(n29751) );
  HS65_LH_BFX2 U5252 ( .A(n29753), .Z(n29752) );
  HS65_LH_BFX2 U5253 ( .A(n29754), .Z(n29753) );
  HS65_LH_BFX2 U5254 ( .A(n29755), .Z(n29754) );
  HS65_LH_BFX2 U5255 ( .A(n29756), .Z(n29755) );
  HS65_LH_BFX2 U5256 ( .A(n29757), .Z(n29756) );
  HS65_LH_BFX2 U5257 ( .A(n29758), .Z(n29757) );
  HS65_LH_BFX2 U5258 ( .A(n29759), .Z(n29758) );
  HS65_LH_BFX2 U5259 ( .A(n29760), .Z(n29759) );
  HS65_LH_BFX2 U5260 ( .A(n29761), .Z(n29760) );
  HS65_LH_BFX2 U5261 ( .A(n29762), .Z(n29761) );
  HS65_LH_BFX2 U5262 ( .A(n29763), .Z(n29762) );
  HS65_LH_BFX2 U5263 ( .A(n29764), .Z(n29763) );
  HS65_LH_BFX2 U5264 ( .A(n17580), .Z(n29764) );
  HS65_LH_BFX2 U5265 ( .A(n34579), .Z(n29765) );
  HS65_LH_BFX2 U5266 ( .A(n17578), .Z(n29766) );
  HS65_LH_BFX2 U5267 ( .A(n29768), .Z(n29767) );
  HS65_LH_BFX2 U5268 ( .A(n29769), .Z(n29768) );
  HS65_LH_BFX2 U5269 ( .A(n33830), .Z(n29769) );
  HS65_LH_BFX2 U5270 ( .A(n18090), .Z(n29770) );
  HS65_LH_BFX2 U5271 ( .A(n18089), .Z(n29771) );
  HS65_LH_BFX2 U5272 ( .A(n29777), .Z(n29772) );
  HS65_LH_BFX2 U5273 ( .A(n29775), .Z(n29773) );
  HS65_LH_IVX2 U5274 ( .A(n29780), .Z(n29774) );
  HS65_LH_IVX2 U5275 ( .A(n29774), .Z(n29775) );
  HS65_LH_IVX2 U5276 ( .A(n29782), .Z(n29776) );
  HS65_LH_IVX2 U5278 ( .A(n29776), .Z(n29777) );
  HS65_LH_BFX2 U5279 ( .A(n18022), .Z(n29778) );
  HS65_LH_IVX2 U5280 ( .A(n29785), .Z(n29779) );
  HS65_LH_IVX2 U5281 ( .A(n29779), .Z(n29780) );
  HS65_LH_IVX2 U5282 ( .A(n29787), .Z(n29781) );
  HS65_LH_IVX2 U5283 ( .A(n29781), .Z(n29782) );
  HS65_LH_BFX2 U5284 ( .A(n29778), .Z(n29783) );
  HS65_LH_IVX2 U5285 ( .A(n29790), .Z(n29784) );
  HS65_LH_IVX2 U5286 ( .A(n29784), .Z(n29785) );
  HS65_LH_IVX2 U5287 ( .A(n29792), .Z(n29786) );
  HS65_LH_IVX2 U5288 ( .A(n29786), .Z(n29787) );
  HS65_LH_BFX2 U5289 ( .A(n29783), .Z(n29788) );
  HS65_LH_IVX2 U5290 ( .A(n29795), .Z(n29789) );
  HS65_LH_IVX2 U5291 ( .A(n29789), .Z(n29790) );
  HS65_LH_IVX2 U5292 ( .A(n29797), .Z(n29791) );
  HS65_LH_IVX2 U5293 ( .A(n29791), .Z(n29792) );
  HS65_LH_BFX2 U5294 ( .A(n29788), .Z(n29793) );
  HS65_LH_IVX2 U5295 ( .A(n29800), .Z(n29794) );
  HS65_LH_IVX2 U5296 ( .A(n29794), .Z(n29795) );
  HS65_LH_IVX2 U5297 ( .A(n29802), .Z(n29796) );
  HS65_LH_IVX2 U5298 ( .A(n29796), .Z(n29797) );
  HS65_LH_BFX2 U5299 ( .A(n29793), .Z(n29798) );
  HS65_LH_IVX2 U5300 ( .A(n29806), .Z(n29799) );
  HS65_LH_IVX2 U5301 ( .A(n29799), .Z(n29800) );
  HS65_LH_IVX2 U5302 ( .A(n29808), .Z(n29801) );
  HS65_LH_IVX2 U5303 ( .A(n29801), .Z(n29802) );
  HS65_LH_BFX2 U5304 ( .A(n29798), .Z(n29803) );
  HS65_LH_BFX2 U5305 ( .A(n29803), .Z(n29804) );
  HS65_LH_IVX2 U5306 ( .A(n29811), .Z(n29805) );
  HS65_LH_IVX2 U5307 ( .A(n29805), .Z(n29806) );
  HS65_LH_IVX2 U5308 ( .A(n29813), .Z(n29807) );
  HS65_LH_IVX2 U5309 ( .A(n29807), .Z(n29808) );
  HS65_LH_BFX2 U5310 ( .A(n29804), .Z(n29809) );
  HS65_LH_IVX2 U5311 ( .A(n29816), .Z(n29810) );
  HS65_LH_IVX2 U5312 ( .A(n29810), .Z(n29811) );
  HS65_LH_IVX2 U5313 ( .A(n29818), .Z(n29812) );
  HS65_LH_IVX2 U5314 ( .A(n29812), .Z(n29813) );
  HS65_LH_BFX2 U5315 ( .A(n29809), .Z(n29814) );
  HS65_LH_IVX2 U5316 ( .A(n29821), .Z(n29815) );
  HS65_LH_IVX2 U5317 ( .A(n29815), .Z(n29816) );
  HS65_LH_IVX2 U5318 ( .A(n29823), .Z(n29817) );
  HS65_LH_IVX2 U5319 ( .A(n29817), .Z(n29818) );
  HS65_LH_BFX2 U5320 ( .A(n29814), .Z(n29819) );
  HS65_LH_IVX2 U5321 ( .A(n29826), .Z(n29820) );
  HS65_LH_IVX2 U5322 ( .A(n29820), .Z(n29821) );
  HS65_LH_IVX2 U5323 ( .A(n29828), .Z(n29822) );
  HS65_LH_IVX2 U5324 ( .A(n29822), .Z(n29823) );
  HS65_LH_BFX2 U5325 ( .A(n29819), .Z(n29824) );
  HS65_LH_IVX2 U5326 ( .A(n29831), .Z(n29825) );
  HS65_LH_IVX2 U5327 ( .A(n29825), .Z(n29826) );
  HS65_LH_IVX2 U5328 ( .A(n29833), .Z(n29827) );
  HS65_LH_IVX2 U5329 ( .A(n29827), .Z(n29828) );
  HS65_LH_BFX2 U5330 ( .A(n29824), .Z(n29829) );
  HS65_LH_IVX2 U5331 ( .A(n29836), .Z(n29830) );
  HS65_LH_IVX2 U5332 ( .A(n29830), .Z(n29831) );
  HS65_LH_IVX2 U5333 ( .A(n29838), .Z(n29832) );
  HS65_LH_IVX2 U5334 ( .A(n29832), .Z(n29833) );
  HS65_LH_BFX2 U5335 ( .A(n29829), .Z(n29834) );
  HS65_LH_IVX2 U5336 ( .A(n29841), .Z(n29835) );
  HS65_LH_IVX2 U5337 ( .A(n29835), .Z(n29836) );
  HS65_LH_IVX2 U5338 ( .A(n29843), .Z(n29837) );
  HS65_LH_IVX2 U5339 ( .A(n29837), .Z(n29838) );
  HS65_LH_BFX2 U5340 ( .A(n29834), .Z(n29839) );
  HS65_LH_IVX2 U5341 ( .A(n29846), .Z(n29840) );
  HS65_LH_IVX2 U5342 ( .A(n29840), .Z(n29841) );
  HS65_LH_IVX2 U5344 ( .A(n29848), .Z(n29842) );
  HS65_LH_IVX2 U5345 ( .A(n29842), .Z(n29843) );
  HS65_LH_BFX2 U5346 ( .A(n29839), .Z(n29844) );
  HS65_LH_IVX2 U5347 ( .A(n29853), .Z(n29845) );
  HS65_LH_IVX2 U5348 ( .A(n29845), .Z(n29846) );
  HS65_LH_IVX2 U5349 ( .A(n29851), .Z(n29847) );
  HS65_LH_IVX2 U5350 ( .A(n29847), .Z(n29848) );
  HS65_LH_BFX2 U5351 ( .A(n29844), .Z(n29849) );
  HS65_LH_IVX2 U5352 ( .A(n29858), .Z(n29850) );
  HS65_LH_IVX2 U5353 ( .A(n29850), .Z(n29851) );
  HS65_LH_IVX2 U5354 ( .A(n29856), .Z(n29852) );
  HS65_LH_IVX2 U5355 ( .A(n29852), .Z(n29853) );
  HS65_LH_BFX2 U5356 ( .A(n29849), .Z(n29854) );
  HS65_LH_IVX2 U5357 ( .A(n29861), .Z(n29855) );
  HS65_LH_IVX2 U5358 ( .A(n29855), .Z(n29856) );
  HS65_LH_BFX2 U5359 ( .A(n29854), .Z(n29857) );
  HS65_LH_BFX2 U5360 ( .A(n29864), .Z(n29858) );
  HS65_LH_BFX2 U5361 ( .A(n29857), .Z(n29859) );
  HS65_LH_IVX2 U5362 ( .A(n18023), .Z(n29860) );
  HS65_LH_IVX2 U5363 ( .A(n29860), .Z(n29861) );
  HS65_LH_IVX2 U5364 ( .A(n29859), .Z(n29862) );
  HS65_LH_IVX2 U5365 ( .A(n29862), .Z(n29863) );
  HS65_LH_BFX2 U5366 ( .A(n18024), .Z(n29864) );
  HS65_LH_BFX2 U5367 ( .A(n29867), .Z(n29865) );
  HS65_LH_IVX2 U5368 ( .A(n29874), .Z(n29866) );
  HS65_LH_IVX2 U5369 ( .A(n29866), .Z(n29867) );
  HS65_LH_BFX2 U5370 ( .A(n29870), .Z(n29868) );
  HS65_LH_BFX2 U5371 ( .A(n18044), .Z(n29869) );
  HS65_LH_BFX2 U5372 ( .A(n29873), .Z(n29870) );
  HS65_LH_BFX2 U5373 ( .A(n29869), .Z(n29871) );
  HS65_LH_IVX2 U5374 ( .A(n29877), .Z(n29872) );
  HS65_LH_IVX2 U5375 ( .A(n29872), .Z(n29873) );
  HS65_LH_BFX2 U5376 ( .A(n38748), .Z(n29874) );
  HS65_LH_BFX2 U5377 ( .A(n29871), .Z(n29875) );
  HS65_LH_IVX2 U5378 ( .A(n38808), .Z(n29876) );
  HS65_LH_IVX2 U5379 ( .A(n29876), .Z(n29877) );
  HS65_LH_BFX2 U5380 ( .A(n29881), .Z(n29878) );
  HS65_LH_BFX2 U5381 ( .A(n29883), .Z(n29879) );
  HS65_LH_IVX2 U5382 ( .A(n29888), .Z(n29880) );
  HS65_LH_IVX2 U5384 ( .A(n29880), .Z(n29881) );
  HS65_LH_IVX2 U5385 ( .A(n29886), .Z(n29882) );
  HS65_LH_IVX2 U5386 ( .A(n29882), .Z(n29883) );
  HS65_LH_BFX2 U5387 ( .A(n18048), .Z(n29884) );
  HS65_LH_IVX2 U5388 ( .A(n29891), .Z(n29885) );
  HS65_LH_IVX2 U5389 ( .A(n29885), .Z(n29886) );
  HS65_LH_BFX2 U5390 ( .A(n29884), .Z(n29887) );
  HS65_LH_BFX2 U5391 ( .A(n29892), .Z(n29888) );
  HS65_LH_BFX2 U5392 ( .A(n29887), .Z(n29889) );
  HS65_LH_IVX2 U5393 ( .A(n29895), .Z(n29890) );
  HS65_LH_IVX2 U5394 ( .A(n29890), .Z(n29891) );
  HS65_LH_BFX2 U5395 ( .A(n29896), .Z(n29892) );
  HS65_LH_BFX2 U5396 ( .A(n29889), .Z(n29893) );
  HS65_LH_IVX2 U5397 ( .A(n29899), .Z(n29894) );
  HS65_LH_IVX2 U5398 ( .A(n29894), .Z(n29895) );
  HS65_LH_BFX2 U5399 ( .A(n29900), .Z(n29896) );
  HS65_LH_BFX2 U5400 ( .A(n29893), .Z(n29897) );
  HS65_LH_IVX2 U5401 ( .A(n38775), .Z(n29898) );
  HS65_LH_IVX2 U5402 ( .A(n29898), .Z(n29899) );
  HS65_LH_BFX2 U5403 ( .A(n38756), .Z(n29900) );
  HS65_LH_BFX2 U5404 ( .A(n29904), .Z(n29901) );
  HS65_LH_BFX2 U5405 ( .A(n29905), .Z(n29902) );
  HS65_LH_BFX2 U5406 ( .A(n38740), .Z(n29903) );
  HS65_LH_BFX2 U5407 ( .A(n38743), .Z(n29904) );
  HS65_LH_BFX2 U5408 ( .A(n38754), .Z(n29905) );
  HS65_LH_BFX2 U5409 ( .A(n29908), .Z(n29906) );
  HS65_LH_IVX2 U5411 ( .A(n29913), .Z(n29907) );
  HS65_LH_IVX2 U5412 ( .A(n29907), .Z(n29908) );
  HS65_LH_BFX2 U5413 ( .A(n29911), .Z(n29909) );
  HS65_LH_BFX2 U5414 ( .A(n18052), .Z(n29910) );
  HS65_LH_BFX2 U5415 ( .A(n29914), .Z(n29911) );
  HS65_LH_BFX2 U5416 ( .A(n29910), .Z(n29912) );
  HS65_LH_BFX2 U5417 ( .A(n29916), .Z(n29913) );
  HS65_LH_BFX2 U5418 ( .A(n29917), .Z(n29914) );
  HS65_LH_BFX2 U5419 ( .A(n29912), .Z(n29915) );
  HS65_LH_BFX2 U5420 ( .A(n29919), .Z(n29916) );
  HS65_LH_BFX2 U5421 ( .A(n29920), .Z(n29917) );
  HS65_LH_BFX2 U5422 ( .A(n29915), .Z(n29918) );
  HS65_LH_BFX2 U5423 ( .A(n29922), .Z(n29919) );
  HS65_LH_BFX2 U5424 ( .A(n29923), .Z(n29920) );
  HS65_LH_BFX2 U5425 ( .A(n29918), .Z(n29921) );
  HS65_LH_BFX2 U5426 ( .A(n29925), .Z(n29922) );
  HS65_LH_BFX2 U5427 ( .A(n29926), .Z(n29923) );
  HS65_LH_BFX2 U5428 ( .A(n29921), .Z(n29924) );
  HS65_LH_BFX2 U5429 ( .A(n29930), .Z(n29925) );
  HS65_LH_BFX2 U5430 ( .A(n29929), .Z(n29926) );
  HS65_LH_BFX2 U5431 ( .A(n29924), .Z(n29927) );
  HS65_LH_IVX2 U5432 ( .A(n29933), .Z(n29928) );
  HS65_LH_IVX2 U5433 ( .A(n29928), .Z(n29929) );
  HS65_LH_BFX2 U5434 ( .A(n29934), .Z(n29930) );
  HS65_LH_BFX2 U5435 ( .A(n29927), .Z(n29931) );
  HS65_LH_IVX2 U5436 ( .A(n38799), .Z(n29932) );
  HS65_LH_IVX2 U5437 ( .A(n29932), .Z(n29933) );
  HS65_LH_BFX2 U5438 ( .A(n38772), .Z(n29934) );
  HS65_LH_BFX2 U5439 ( .A(n29937), .Z(n29935) );
  HS65_LH_IVX2 U5440 ( .A(n29942), .Z(n29936) );
  HS65_LH_IVX2 U5441 ( .A(n29936), .Z(n29937) );
  HS65_LH_BFX2 U5442 ( .A(n18046), .Z(n29938) );
  HS65_LH_BFX2 U5443 ( .A(n29941), .Z(n29939) );
  HS65_LH_BFX2 U5444 ( .A(n29938), .Z(n29940) );
  HS65_LH_BFX2 U5445 ( .A(n29944), .Z(n29941) );
  HS65_LH_BFX2 U5446 ( .A(n29945), .Z(n29942) );
  HS65_LH_BFX2 U5447 ( .A(n29940), .Z(n29943) );
  HS65_LH_BFX2 U5448 ( .A(n29949), .Z(n29944) );
  HS65_LH_BFX2 U5449 ( .A(n29948), .Z(n29945) );
  HS65_LH_BFX2 U5450 ( .A(n29943), .Z(n29946) );
  HS65_LH_IVX2 U5451 ( .A(n29952), .Z(n29947) );
  HS65_LH_IVX2 U5452 ( .A(n29947), .Z(n29948) );
  HS65_LH_BFX2 U5453 ( .A(n29953), .Z(n29949) );
  HS65_LH_BFX2 U5454 ( .A(n29946), .Z(n29950) );
  HS65_LH_IVX2 U5455 ( .A(n38800), .Z(n29951) );
  HS65_LH_IVX2 U5456 ( .A(n29951), .Z(n29952) );
  HS65_LH_BFX2 U5457 ( .A(n38770), .Z(n29953) );
  HS65_LH_BFX2 U5458 ( .A(n39018), .Z(n29954) );
  HS65_LH_IVX2 U5459 ( .A(n18058), .Z(n39065) );
  HS65_LH_BFX2 U5460 ( .A(n29960), .Z(n29955) );
  HS65_LH_BFX2 U5461 ( .A(n29958), .Z(n29956) );
  HS65_LH_IVX2 U5462 ( .A(n29963), .Z(n29957) );
  HS65_LH_IVX2 U5463 ( .A(n29957), .Z(n29958) );
  HS65_LH_IVX2 U5464 ( .A(n29965), .Z(n29959) );
  HS65_LH_IVX2 U5465 ( .A(n29959), .Z(n29960) );
  HS65_LH_BFX2 U5466 ( .A(n18057), .Z(n29961) );
  HS65_LH_IVX2 U5467 ( .A(n29968), .Z(n29962) );
  HS65_LH_IVX2 U5468 ( .A(n29962), .Z(n29963) );
  HS65_LH_IVX2 U5469 ( .A(n29970), .Z(n29964) );
  HS65_LH_IVX2 U5470 ( .A(n29964), .Z(n29965) );
  HS65_LH_BFX2 U5471 ( .A(n29961), .Z(n29966) );
  HS65_LH_IVX2 U5472 ( .A(n29973), .Z(n29967) );
  HS65_LH_IVX2 U5473 ( .A(n29967), .Z(n29968) );
  HS65_LH_IVX2 U5474 ( .A(n29975), .Z(n29969) );
  HS65_LH_IVX2 U5475 ( .A(n29969), .Z(n29970) );
  HS65_LH_BFX2 U5476 ( .A(n29966), .Z(n29971) );
  HS65_LH_IVX2 U5477 ( .A(n29978), .Z(n29972) );
  HS65_LH_IVX2 U5478 ( .A(n29972), .Z(n29973) );
  HS65_LH_IVX2 U5479 ( .A(n29980), .Z(n29974) );
  HS65_LH_IVX2 U5480 ( .A(n29974), .Z(n29975) );
  HS65_LH_BFX2 U5481 ( .A(n29971), .Z(n29976) );
  HS65_LH_IVX2 U5482 ( .A(n29984), .Z(n29977) );
  HS65_LH_IVX2 U5483 ( .A(n29977), .Z(n29978) );
  HS65_LH_IVX2 U5484 ( .A(n29986), .Z(n29979) );
  HS65_LH_IVX2 U5485 ( .A(n29979), .Z(n29980) );
  HS65_LH_BFX2 U5486 ( .A(n29976), .Z(n29981) );
  HS65_LH_BFX2 U5487 ( .A(n29981), .Z(n29982) );
  HS65_LH_IVX2 U5488 ( .A(n29989), .Z(n29983) );
  HS65_LH_IVX2 U5489 ( .A(n29983), .Z(n29984) );
  HS65_LH_IVX2 U5490 ( .A(n29991), .Z(n29985) );
  HS65_LH_IVX2 U5491 ( .A(n29985), .Z(n29986) );
  HS65_LH_BFX2 U5492 ( .A(n29982), .Z(n29987) );
  HS65_LH_IVX2 U5493 ( .A(n29994), .Z(n29988) );
  HS65_LH_IVX2 U5494 ( .A(n29988), .Z(n29989) );
  HS65_LH_IVX2 U5495 ( .A(n29996), .Z(n29990) );
  HS65_LH_IVX2 U5496 ( .A(n29990), .Z(n29991) );
  HS65_LH_BFX2 U5497 ( .A(n29987), .Z(n29992) );
  HS65_LH_IVX2 U5498 ( .A(n29999), .Z(n29993) );
  HS65_LH_IVX2 U5499 ( .A(n29993), .Z(n29994) );
  HS65_LH_IVX2 U5500 ( .A(n30001), .Z(n29995) );
  HS65_LH_IVX2 U5501 ( .A(n29995), .Z(n29996) );
  HS65_LH_BFX2 U5502 ( .A(n29992), .Z(n29997) );
  HS65_LH_IVX2 U5503 ( .A(n38735), .Z(n29998) );
  HS65_LH_IVX2 U5504 ( .A(n29998), .Z(n29999) );
  HS65_LH_IVX2 U5505 ( .A(n38738), .Z(n30000) );
  HS65_LH_IVX2 U5506 ( .A(n30000), .Z(n30001) );
  HS65_LH_BFX2 U5507 ( .A(n29997), .Z(n30002) );
  HS65_LH_BFX2 U5508 ( .A(n30006), .Z(n30003) );
  HS65_LH_BFX2 U5509 ( .A(n18050), .Z(n30004) );
  HS65_LH_BFX2 U5510 ( .A(n30008), .Z(n30005) );
  HS65_LH_BFX2 U5511 ( .A(n30009), .Z(n30006) );
  HS65_LH_BFX2 U5512 ( .A(n30004), .Z(n30007) );
  HS65_LH_BFX2 U5513 ( .A(n30011), .Z(n30008) );
  HS65_LH_BFX2 U5514 ( .A(n30012), .Z(n30009) );
  HS65_LH_BFX2 U5515 ( .A(n30007), .Z(n30010) );
  HS65_LH_BFX2 U5516 ( .A(n30014), .Z(n30011) );
  HS65_LH_BFX2 U5517 ( .A(n30015), .Z(n30012) );
  HS65_LH_BFX2 U5518 ( .A(n30010), .Z(n30013) );
  HS65_LH_BFX2 U5519 ( .A(n30017), .Z(n30014) );
  HS65_LH_BFX2 U5520 ( .A(n30018), .Z(n30015) );
  HS65_LH_BFX2 U5521 ( .A(n30013), .Z(n30016) );
  HS65_LH_BFX2 U5522 ( .A(n30020), .Z(n30017) );
  HS65_LH_BFX2 U5523 ( .A(n30021), .Z(n30018) );
  HS65_LH_BFX2 U5524 ( .A(n30016), .Z(n30019) );
  HS65_LH_BFX2 U5525 ( .A(n30025), .Z(n30020) );
  HS65_LH_BFX2 U5526 ( .A(n30026), .Z(n30021) );
  HS65_LH_BFX2 U5527 ( .A(n30019), .Z(n30022) );
  HS65_LH_IVX2 U5528 ( .A(n38955), .Z(n30023) );
  HS65_LH_IVX2 U5529 ( .A(n30023), .Z(n30024) );
  HS65_LH_BFX2 U5530 ( .A(n38749), .Z(n30025) );
  HS65_LH_BFX2 U5531 ( .A(n38767), .Z(n30026) );
  HS65_LH_BFX2 U5532 ( .A(n30062), .Z(n30027) );
  HS65_LH_IVX2 U5533 ( .A(n18063), .Z(n38982) );
  HS65_LH_BFX2 U5534 ( .A(n30033), .Z(n30028) );
  HS65_LH_BFX2 U5535 ( .A(n30031), .Z(n30029) );
  HS65_LH_IVX2 U5542 ( .A(n30036), .Z(n30030) );
  HS65_LH_IVX2 U5543 ( .A(n30030), .Z(n30031) );
  HS65_LH_IVX2 U5544 ( .A(n30038), .Z(n30032) );
  HS65_LH_IVX2 U5545 ( .A(n30032), .Z(n30033) );
  HS65_LH_BFX2 U5546 ( .A(n18061), .Z(n30034) );
  HS65_LH_IVX2 U5547 ( .A(n30041), .Z(n30035) );
  HS65_LH_IVX2 U5548 ( .A(n30035), .Z(n30036) );
  HS65_LH_IVX2 U5549 ( .A(n30043), .Z(n30037) );
  HS65_LH_IVX2 U5550 ( .A(n30037), .Z(n30038) );
  HS65_LH_BFX2 U5551 ( .A(n30034), .Z(n30039) );
  HS65_LH_IVX2 U5552 ( .A(n30046), .Z(n30040) );
  HS65_LH_IVX2 U5553 ( .A(n30040), .Z(n30041) );
  HS65_LH_IVX2 U5554 ( .A(n30048), .Z(n30042) );
  HS65_LH_IVX2 U5555 ( .A(n30042), .Z(n30043) );
  HS65_LH_BFX2 U5556 ( .A(n30039), .Z(n30044) );
  HS65_LH_IVX2 U5557 ( .A(n30051), .Z(n30045) );
  HS65_LH_IVX2 U5558 ( .A(n30045), .Z(n30046) );
  HS65_LH_IVX2 U5559 ( .A(n30053), .Z(n30047) );
  HS65_LH_IVX2 U5560 ( .A(n30047), .Z(n30048) );
  HS65_LH_BFX2 U5561 ( .A(n30044), .Z(n30049) );
  HS65_LH_IVX2 U5562 ( .A(n30057), .Z(n30050) );
  HS65_LH_IVX2 U5563 ( .A(n30050), .Z(n30051) );
  HS65_LH_IVX2 U5564 ( .A(n30059), .Z(n30052) );
  HS65_LH_IVX2 U5565 ( .A(n30052), .Z(n30053) );
  HS65_LH_BFX2 U5566 ( .A(n30049), .Z(n30054) );
  HS65_LH_BFX2 U5567 ( .A(n30054), .Z(n30055) );
  HS65_LH_IVX2 U5568 ( .A(n30064), .Z(n30056) );
  HS65_LH_IVX2 U5569 ( .A(n30056), .Z(n30057) );
  HS65_LH_IVX2 U5570 ( .A(n30066), .Z(n30058) );
  HS65_LH_IVX2 U5571 ( .A(n30058), .Z(n30059) );
  HS65_LH_BFX2 U5572 ( .A(n30055), .Z(n30060) );
  HS65_LH_IVX2 U5573 ( .A(n38998), .Z(n30061) );
  HS65_LH_IVX2 U5574 ( .A(n30061), .Z(n30062) );
  HS65_LH_IVX2 U5575 ( .A(n30069), .Z(n30063) );
  HS65_LH_IVX2 U5576 ( .A(n30063), .Z(n30064) );
  HS65_LH_IVX2 U5577 ( .A(n30071), .Z(n30065) );
  HS65_LH_IVX2 U5578 ( .A(n30065), .Z(n30066) );
  HS65_LH_BFX2 U5579 ( .A(n30060), .Z(n30067) );
  HS65_LH_IVX2 U5580 ( .A(n30074), .Z(n30068) );
  HS65_LH_IVX2 U5581 ( .A(n30068), .Z(n30069) );
  HS65_LH_IVX2 U5582 ( .A(n30076), .Z(n30070) );
  HS65_LH_IVX2 U5583 ( .A(n30070), .Z(n30071) );
  HS65_LH_BFX2 U5584 ( .A(n30067), .Z(n30072) );
  HS65_LH_IVX2 U5585 ( .A(n30079), .Z(n30073) );
  HS65_LH_IVX2 U5586 ( .A(n30073), .Z(n30074) );
  HS65_LH_IVX2 U5587 ( .A(n30081), .Z(n30075) );
  HS65_LH_IVX2 U5588 ( .A(n30075), .Z(n30076) );
  HS65_LH_BFX2 U5589 ( .A(n30072), .Z(n30077) );
  HS65_LH_IVX2 U5590 ( .A(n30084), .Z(n30078) );
  HS65_LH_IVX2 U5591 ( .A(n30078), .Z(n30079) );
  HS65_LH_IVX2 U5592 ( .A(n30086), .Z(n30080) );
  HS65_LH_IVX2 U5593 ( .A(n30080), .Z(n30081) );
  HS65_LH_BFX2 U5594 ( .A(n30077), .Z(n30082) );
  HS65_LH_IVX2 U5595 ( .A(n30089), .Z(n30083) );
  HS65_LH_IVX2 U5596 ( .A(n30083), .Z(n30084) );
  HS65_LH_IVX2 U5597 ( .A(n30091), .Z(n30085) );
  HS65_LH_IVX2 U5598 ( .A(n30085), .Z(n30086) );
  HS65_LH_BFX2 U5599 ( .A(n30082), .Z(n30087) );
  HS65_LH_IVX2 U5600 ( .A(n38758), .Z(n30088) );
  HS65_LH_IVX2 U5601 ( .A(n30088), .Z(n30089) );
  HS65_LH_IVX2 U5602 ( .A(n38760), .Z(n30090) );
  HS65_LH_IVX2 U5603 ( .A(n30090), .Z(n30091) );
  HS65_LH_BFX2 U5605 ( .A(n30095), .Z(n30092) );
  HS65_LH_BFX2 U5606 ( .A(n30096), .Z(n30093) );
  HS65_LH_BFX2 U5607 ( .A(n18054), .Z(n30094) );
  HS65_LH_BFX2 U5608 ( .A(n30098), .Z(n30095) );
  HS65_LH_BFX2 U5609 ( .A(n30099), .Z(n30096) );
  HS65_LH_BFX2 U5610 ( .A(n30094), .Z(n30097) );
  HS65_LH_BFX2 U5611 ( .A(n30101), .Z(n30098) );
  HS65_LH_BFX2 U5612 ( .A(n30102), .Z(n30099) );
  HS65_LH_BFX2 U5613 ( .A(n30097), .Z(n30100) );
  HS65_LH_BFX2 U5614 ( .A(n30104), .Z(n30101) );
  HS65_LH_BFX2 U5615 ( .A(n30105), .Z(n30102) );
  HS65_LH_BFX2 U5616 ( .A(n30100), .Z(n30103) );
  HS65_LH_BFX2 U5617 ( .A(n30107), .Z(n30104) );
  HS65_LH_BFX2 U5618 ( .A(n30108), .Z(n30105) );
  HS65_LH_BFX2 U5619 ( .A(n30103), .Z(n30106) );
  HS65_LH_BFX2 U5620 ( .A(n30110), .Z(n30107) );
  HS65_LH_BFX2 U5621 ( .A(n30111), .Z(n30108) );
  HS65_LH_BFX2 U5622 ( .A(n30106), .Z(n30109) );
  HS65_LH_BFX2 U5623 ( .A(n30113), .Z(n30110) );
  HS65_LH_BFX2 U5624 ( .A(n30114), .Z(n30111) );
  HS65_LH_BFX2 U5625 ( .A(n30109), .Z(n30112) );
  HS65_LH_BFX2 U5626 ( .A(n30116), .Z(n30113) );
  HS65_LH_BFX2 U5627 ( .A(n30117), .Z(n30114) );
  HS65_LH_BFX2 U5628 ( .A(n30112), .Z(n30115) );
  HS65_LH_BFX2 U5629 ( .A(n30121), .Z(n30116) );
  HS65_LH_BFX2 U5630 ( .A(n30120), .Z(n30117) );
  HS65_LH_BFX2 U5631 ( .A(n30115), .Z(n30118) );
  HS65_LH_IVX2 U5632 ( .A(n30124), .Z(n30119) );
  HS65_LH_IVX2 U5633 ( .A(n30119), .Z(n30120) );
  HS65_LH_BFX2 U5634 ( .A(n38747), .Z(n30121) );
  HS65_LH_BFX2 U5635 ( .A(n30118), .Z(n30122) );
  HS65_LH_IVX2 U5636 ( .A(n38806), .Z(n30123) );
  HS65_LH_IVX2 U5637 ( .A(n30123), .Z(n30124) );
  HS65_LH_BFX2 U5638 ( .A(n38899), .Z(n30125) );
  HS65_LH_IVX2 U5639 ( .A(n18068), .Z(n38882) );
  HS65_LH_BFX2 U5640 ( .A(n30131), .Z(n30126) );
  HS65_LH_BFX2 U5641 ( .A(n30129), .Z(n30127) );
  HS65_LH_IVX2 U5642 ( .A(n30134), .Z(n30128) );
  HS65_LH_IVX2 U5643 ( .A(n30128), .Z(n30129) );
  HS65_LH_IVX2 U5644 ( .A(n30136), .Z(n30130) );
  HS65_LH_IVX2 U5645 ( .A(n30130), .Z(n30131) );
  HS65_LH_BFX2 U5646 ( .A(n18066), .Z(n30132) );
  HS65_LH_IVX2 U5647 ( .A(n30139), .Z(n30133) );
  HS65_LH_IVX2 U5648 ( .A(n30133), .Z(n30134) );
  HS65_LH_IVX2 U5649 ( .A(n30141), .Z(n30135) );
  HS65_LH_IVX2 U5650 ( .A(n30135), .Z(n30136) );
  HS65_LH_BFX2 U5651 ( .A(n30132), .Z(n30137) );
  HS65_LH_IVX2 U5652 ( .A(n30144), .Z(n30138) );
  HS65_LH_IVX2 U5653 ( .A(n30138), .Z(n30139) );
  HS65_LH_IVX2 U5654 ( .A(n30146), .Z(n30140) );
  HS65_LH_IVX2 U5655 ( .A(n30140), .Z(n30141) );
  HS65_LH_BFX2 U5656 ( .A(n30137), .Z(n30142) );
  HS65_LH_IVX2 U5657 ( .A(n30149), .Z(n30143) );
  HS65_LH_IVX2 U5658 ( .A(n30143), .Z(n30144) );
  HS65_LH_IVX2 U5659 ( .A(n30151), .Z(n30145) );
  HS65_LH_IVX2 U5660 ( .A(n30145), .Z(n30146) );
  HS65_LH_BFX2 U5661 ( .A(n30142), .Z(n30147) );
  HS65_LH_IVX2 U5662 ( .A(n30154), .Z(n30148) );
  HS65_LH_IVX2 U5663 ( .A(n30148), .Z(n30149) );
  HS65_LH_IVX2 U5664 ( .A(n30156), .Z(n30150) );
  HS65_LH_IVX2 U5665 ( .A(n30150), .Z(n30151) );
  HS65_LH_BFX2 U5666 ( .A(n30147), .Z(n30152) );
  HS65_LH_IVX2 U5667 ( .A(n30160), .Z(n30153) );
  HS65_LH_IVX2 U5669 ( .A(n30153), .Z(n30154) );
  HS65_LH_IVX2 U5670 ( .A(n30162), .Z(n30155) );
  HS65_LH_IVX2 U5671 ( .A(n30155), .Z(n30156) );
  HS65_LH_BFX2 U5672 ( .A(n30152), .Z(n30157) );
  HS65_LH_BFX2 U5673 ( .A(n30157), .Z(n30158) );
  HS65_LH_IVX2 U5674 ( .A(n30165), .Z(n30159) );
  HS65_LH_IVX2 U5675 ( .A(n30159), .Z(n30160) );
  HS65_LH_IVX2 U5676 ( .A(n30167), .Z(n30161) );
  HS65_LH_IVX2 U5677 ( .A(n30161), .Z(n30162) );
  HS65_LH_BFX2 U5678 ( .A(n30158), .Z(n30163) );
  HS65_LH_IVX2 U5679 ( .A(n30170), .Z(n30164) );
  HS65_LH_IVX2 U5680 ( .A(n30164), .Z(n30165) );
  HS65_LH_IVX2 U5681 ( .A(n30172), .Z(n30166) );
  HS65_LH_IVX2 U5682 ( .A(n30166), .Z(n30167) );
  HS65_LH_BFX2 U5683 ( .A(n30163), .Z(n30168) );
  HS65_LH_IVX2 U5684 ( .A(n30175), .Z(n30169) );
  HS65_LH_IVX2 U5685 ( .A(n30169), .Z(n30170) );
  HS65_LH_IVX2 U5686 ( .A(n30177), .Z(n30171) );
  HS65_LH_IVX2 U5687 ( .A(n30171), .Z(n30172) );
  HS65_LH_BFX2 U5688 ( .A(n30168), .Z(n30173) );
  HS65_LH_IVX2 U5689 ( .A(n30180), .Z(n30174) );
  HS65_LH_IVX2 U5690 ( .A(n30174), .Z(n30175) );
  HS65_LH_IVX2 U5691 ( .A(n30182), .Z(n30176) );
  HS65_LH_IVX2 U5692 ( .A(n30176), .Z(n30177) );
  HS65_LH_BFX2 U5693 ( .A(n30173), .Z(n30178) );
  HS65_LH_IVX2 U5694 ( .A(n30185), .Z(n30179) );
  HS65_LH_IVX2 U5695 ( .A(n30179), .Z(n30180) );
  HS65_LH_IVX2 U5696 ( .A(n30187), .Z(n30181) );
  HS65_LH_IVX2 U5697 ( .A(n30181), .Z(n30182) );
  HS65_LH_BFX2 U5698 ( .A(n30178), .Z(n30183) );
  HS65_LH_IVX2 U5699 ( .A(n30190), .Z(n30184) );
  HS65_LH_IVX2 U5700 ( .A(n30184), .Z(n30185) );
  HS65_LH_IVX2 U5701 ( .A(n30192), .Z(n30186) );
  HS65_LH_IVX2 U5702 ( .A(n30186), .Z(n30187) );
  HS65_LH_BFX2 U5703 ( .A(n30183), .Z(n30188) );
  HS65_LH_IVX2 U5704 ( .A(n30195), .Z(n30189) );
  HS65_LH_IVX2 U5705 ( .A(n30189), .Z(n30190) );
  HS65_LH_IVX2 U5706 ( .A(n30197), .Z(n30191) );
  HS65_LH_IVX2 U5707 ( .A(n30191), .Z(n30192) );
  HS65_LH_BFX2 U5708 ( .A(n30188), .Z(n30193) );
  HS65_LH_IVX2 U5709 ( .A(n38742), .Z(n30194) );
  HS65_LH_IVX2 U5710 ( .A(n30194), .Z(n30195) );
  HS65_LH_IVX2 U5711 ( .A(n38745), .Z(n30196) );
  HS65_LH_IVX2 U5712 ( .A(n30196), .Z(n30197) );
  HS65_LH_BFX2 U5713 ( .A(n30193), .Z(n30198) );
  HS65_LH_BFX2 U5714 ( .A(n30202), .Z(n30199) );
  HS65_LH_BFX2 U5715 ( .A(n30203), .Z(n30200) );
  HS65_LH_BFX2 U5716 ( .A(n18059), .Z(n30201) );
  HS65_LH_BFX2 U5717 ( .A(n30205), .Z(n30202) );
  HS65_LH_BFX2 U5718 ( .A(n30206), .Z(n30203) );
  HS65_LH_BFX2 U5719 ( .A(n30201), .Z(n30204) );
  HS65_LH_BFX2 U5720 ( .A(n30208), .Z(n30205) );
  HS65_LH_BFX2 U5721 ( .A(n30209), .Z(n30206) );
  HS65_LH_BFX2 U5722 ( .A(n30204), .Z(n30207) );
  HS65_LH_BFX2 U5723 ( .A(n30211), .Z(n30208) );
  HS65_LH_BFX2 U5724 ( .A(n30212), .Z(n30209) );
  HS65_LH_BFX2 U5725 ( .A(n30207), .Z(n30210) );
  HS65_LH_BFX2 U5726 ( .A(n30214), .Z(n30211) );
  HS65_LH_BFX2 U5727 ( .A(n30215), .Z(n30212) );
  HS65_LH_BFX2 U5728 ( .A(n30210), .Z(n30213) );
  HS65_LH_BFX2 U5729 ( .A(n30217), .Z(n30214) );
  HS65_LH_BFX2 U5730 ( .A(n30218), .Z(n30215) );
  HS65_LH_BFX2 U5731 ( .A(n30213), .Z(n30216) );
  HS65_LH_BFX2 U5732 ( .A(n30220), .Z(n30217) );
  HS65_LH_BFX2 U5733 ( .A(n30221), .Z(n30218) );
  HS65_LH_BFX2 U5734 ( .A(n30216), .Z(n30219) );
  HS65_LH_BFX2 U5736 ( .A(n30223), .Z(n30220) );
  HS65_LH_BFX2 U5737 ( .A(n30224), .Z(n30221) );
  HS65_LH_BFX2 U5738 ( .A(n30219), .Z(n30222) );
  HS65_LH_BFX2 U5739 ( .A(n30226), .Z(n30223) );
  HS65_LH_BFX2 U5740 ( .A(n30227), .Z(n30224) );
  HS65_LH_BFX2 U5741 ( .A(n30222), .Z(n30225) );
  HS65_LH_BFX2 U5742 ( .A(n30229), .Z(n30226) );
  HS65_LH_BFX2 U5743 ( .A(n30230), .Z(n30227) );
  HS65_LH_BFX2 U5744 ( .A(n30225), .Z(n30228) );
  HS65_LH_BFX2 U5745 ( .A(n30232), .Z(n30229) );
  HS65_LH_BFX2 U5746 ( .A(n30233), .Z(n30230) );
  HS65_LH_BFX2 U5747 ( .A(n30228), .Z(n30231) );
  HS65_LH_BFX2 U5748 ( .A(n30237), .Z(n30232) );
  HS65_LH_BFX2 U5749 ( .A(n30236), .Z(n30233) );
  HS65_LH_BFX2 U5750 ( .A(n30231), .Z(n30234) );
  HS65_LH_IVX2 U5751 ( .A(n38773), .Z(n30235) );
  HS65_LH_IVX2 U5752 ( .A(n30235), .Z(n30236) );
  HS65_LH_BFX2 U5753 ( .A(n38753), .Z(n30237) );
  HS65_LH_BFX2 U5754 ( .A(n38782), .Z(n30238) );
  HS65_LH_IVX2 U5755 ( .A(n18073), .Z(n38764) );
  HS65_LH_BFX2 U5756 ( .A(n30244), .Z(n30239) );
  HS65_LH_BFX2 U5757 ( .A(n30242), .Z(n30240) );
  HS65_LH_IVX2 U5758 ( .A(n30247), .Z(n30241) );
  HS65_LH_IVX2 U5759 ( .A(n30241), .Z(n30242) );
  HS65_LH_IVX2 U5760 ( .A(n30249), .Z(n30243) );
  HS65_LH_IVX2 U5761 ( .A(n30243), .Z(n30244) );
  HS65_LH_BFX2 U5762 ( .A(n18071), .Z(n30245) );
  HS65_LH_IVX2 U5763 ( .A(n30252), .Z(n30246) );
  HS65_LH_IVX2 U5764 ( .A(n30246), .Z(n30247) );
  HS65_LH_IVX2 U5765 ( .A(n30254), .Z(n30248) );
  HS65_LH_IVX2 U5766 ( .A(n30248), .Z(n30249) );
  HS65_LH_BFX2 U5767 ( .A(n30245), .Z(n30250) );
  HS65_LH_IVX2 U5768 ( .A(n30257), .Z(n30251) );
  HS65_LH_IVX2 U5769 ( .A(n30251), .Z(n30252) );
  HS65_LH_IVX2 U5770 ( .A(n30259), .Z(n30253) );
  HS65_LH_IVX2 U5771 ( .A(n30253), .Z(n30254) );
  HS65_LH_BFX2 U5772 ( .A(n30250), .Z(n30255) );
  HS65_LH_IVX2 U5773 ( .A(n30262), .Z(n30256) );
  HS65_LH_IVX2 U5774 ( .A(n30256), .Z(n30257) );
  HS65_LH_IVX2 U5775 ( .A(n30264), .Z(n30258) );
  HS65_LH_IVX2 U5776 ( .A(n30258), .Z(n30259) );
  HS65_LH_BFX2 U5777 ( .A(n30255), .Z(n30260) );
  HS65_LH_IVX2 U5778 ( .A(n30267), .Z(n30261) );
  HS65_LH_IVX2 U5779 ( .A(n30261), .Z(n30262) );
  HS65_LH_IVX2 U5780 ( .A(n30269), .Z(n30263) );
  HS65_LH_IVX2 U5781 ( .A(n30263), .Z(n30264) );
  HS65_LH_BFX2 U5782 ( .A(n30260), .Z(n30265) );
  HS65_LH_IVX2 U5783 ( .A(n30273), .Z(n30266) );
  HS65_LH_IVX2 U5784 ( .A(n30266), .Z(n30267) );
  HS65_LH_IVX2 U5785 ( .A(n30275), .Z(n30268) );
  HS65_LH_IVX2 U5786 ( .A(n30268), .Z(n30269) );
  HS65_LH_BFX2 U5787 ( .A(n30265), .Z(n30270) );
  HS65_LH_BFX2 U5788 ( .A(n30270), .Z(n30271) );
  HS65_LH_IVX2 U5789 ( .A(n30278), .Z(n30272) );
  HS65_LH_IVX2 U5790 ( .A(n30272), .Z(n30273) );
  HS65_LH_IVX2 U5791 ( .A(n30280), .Z(n30274) );
  HS65_LH_IVX2 U5792 ( .A(n30274), .Z(n30275) );
  HS65_LH_BFX2 U5793 ( .A(n30271), .Z(n30276) );
  HS65_LH_IVX2 U5794 ( .A(n30283), .Z(n30277) );
  HS65_LH_IVX2 U5795 ( .A(n30277), .Z(n30278) );
  HS65_LH_IVX2 U5796 ( .A(n30285), .Z(n30279) );
  HS65_LH_IVX2 U5797 ( .A(n30279), .Z(n30280) );
  HS65_LH_BFX2 U5798 ( .A(n30276), .Z(n30281) );
  HS65_LH_IVX2 U5799 ( .A(n30288), .Z(n30282) );
  HS65_LH_IVX2 U5800 ( .A(n30282), .Z(n30283) );
  HS65_LH_IVX2 U5802 ( .A(n30290), .Z(n30284) );
  HS65_LH_IVX2 U5805 ( .A(n30284), .Z(n30285) );
  HS65_LH_BFX2 U5806 ( .A(n30281), .Z(n30286) );
  HS65_LH_IVX2 U5807 ( .A(n30293), .Z(n30287) );
  HS65_LH_IVX2 U5808 ( .A(n30287), .Z(n30288) );
  HS65_LH_IVX2 U5809 ( .A(n30295), .Z(n30289) );
  HS65_LH_IVX2 U5810 ( .A(n30289), .Z(n30290) );
  HS65_LH_BFX2 U5811 ( .A(n30286), .Z(n30291) );
  HS65_LH_IVX2 U5812 ( .A(n30298), .Z(n30292) );
  HS65_LH_IVX2 U5813 ( .A(n30292), .Z(n30293) );
  HS65_LH_IVX2 U5814 ( .A(n30300), .Z(n30294) );
  HS65_LH_IVX2 U5815 ( .A(n30294), .Z(n30295) );
  HS65_LH_BFX2 U5816 ( .A(n30291), .Z(n30296) );
  HS65_LH_IVX2 U5817 ( .A(n30303), .Z(n30297) );
  HS65_LH_IVX2 U5818 ( .A(n30297), .Z(n30298) );
  HS65_LH_IVX2 U5819 ( .A(n30305), .Z(n30299) );
  HS65_LH_IVX2 U5820 ( .A(n30299), .Z(n30300) );
  HS65_LH_BFX2 U5821 ( .A(n30296), .Z(n30301) );
  HS65_LH_IVX2 U5822 ( .A(n30308), .Z(n30302) );
  HS65_LH_IVX2 U5823 ( .A(n30302), .Z(n30303) );
  HS65_LH_IVX2 U5824 ( .A(n30310), .Z(n30304) );
  HS65_LH_IVX2 U5825 ( .A(n30304), .Z(n30305) );
  HS65_LH_BFX2 U5826 ( .A(n30301), .Z(n30306) );
  HS65_LH_IVX2 U5827 ( .A(n30313), .Z(n30307) );
  HS65_LH_IVX2 U5828 ( .A(n30307), .Z(n30308) );
  HS65_LH_IVX2 U5829 ( .A(n30315), .Z(n30309) );
  HS65_LH_IVX2 U5830 ( .A(n30309), .Z(n30310) );
  HS65_LH_BFX2 U5831 ( .A(n30306), .Z(n30311) );
  HS65_LH_IVX2 U5832 ( .A(n30318), .Z(n30312) );
  HS65_LH_IVX2 U5833 ( .A(n30312), .Z(n30313) );
  HS65_LH_IVX2 U5834 ( .A(n30320), .Z(n30314) );
  HS65_LH_IVX2 U5835 ( .A(n30314), .Z(n30315) );
  HS65_LH_BFX2 U5836 ( .A(n30311), .Z(n30316) );
  HS65_LH_IVX2 U5837 ( .A(n38755), .Z(n30317) );
  HS65_LH_IVX2 U5838 ( .A(n30317), .Z(n30318) );
  HS65_LH_IVX2 U5839 ( .A(n30323), .Z(n30319) );
  HS65_LH_IVX2 U5840 ( .A(n30319), .Z(n30320) );
  HS65_LH_BFX2 U5841 ( .A(n30316), .Z(n30321) );
  HS65_LH_IVX2 U5842 ( .A(n38765), .Z(n30322) );
  HS65_LH_IVX2 U5843 ( .A(n30322), .Z(n30323) );
  HS65_LH_BFX2 U5844 ( .A(n30327), .Z(n30324) );
  HS65_LH_BFX2 U5845 ( .A(n30328), .Z(n30325) );
  HS65_LH_BFX2 U5846 ( .A(n18064), .Z(n30326) );
  HS65_LH_BFX2 U5847 ( .A(n30330), .Z(n30327) );
  HS65_LH_BFX2 U5848 ( .A(n30331), .Z(n30328) );
  HS65_LH_BFX2 U5849 ( .A(n30326), .Z(n30329) );
  HS65_LH_BFX2 U5850 ( .A(n30333), .Z(n30330) );
  HS65_LH_BFX2 U5851 ( .A(n30334), .Z(n30331) );
  HS65_LH_BFX2 U5852 ( .A(n30329), .Z(n30332) );
  HS65_LH_BFX2 U5853 ( .A(n30336), .Z(n30333) );
  HS65_LH_BFX2 U5854 ( .A(n30337), .Z(n30334) );
  HS65_LH_BFX2 U5855 ( .A(n30332), .Z(n30335) );
  HS65_LH_BFX2 U5856 ( .A(n30339), .Z(n30336) );
  HS65_LH_BFX2 U5857 ( .A(n30340), .Z(n30337) );
  HS65_LH_BFX2 U5858 ( .A(n30335), .Z(n30338) );
  HS65_LH_BFX2 U5859 ( .A(n30342), .Z(n30339) );
  HS65_LH_BFX2 U5860 ( .A(n30343), .Z(n30340) );
  HS65_LH_BFX2 U5861 ( .A(n30338), .Z(n30341) );
  HS65_LH_BFX2 U5862 ( .A(n30345), .Z(n30342) );
  HS65_LH_BFX2 U5863 ( .A(n30346), .Z(n30343) );
  HS65_LH_BFX2 U5864 ( .A(n30341), .Z(n30344) );
  HS65_LH_BFX2 U5865 ( .A(n30348), .Z(n30345) );
  HS65_LH_BFX2 U5866 ( .A(n30349), .Z(n30346) );
  HS65_LH_BFX2 U5868 ( .A(n30344), .Z(n30347) );
  HS65_LH_BFX2 U5869 ( .A(n30351), .Z(n30348) );
  HS65_LH_BFX2 U5870 ( .A(n30352), .Z(n30349) );
  HS65_LH_BFX2 U5871 ( .A(n30347), .Z(n30350) );
  HS65_LH_BFX2 U5872 ( .A(n30354), .Z(n30351) );
  HS65_LH_BFX2 U5873 ( .A(n30355), .Z(n30352) );
  HS65_LH_BFX2 U5874 ( .A(n30350), .Z(n30353) );
  HS65_LH_BFX2 U5875 ( .A(n30357), .Z(n30354) );
  HS65_LH_BFX2 U5876 ( .A(n30358), .Z(n30355) );
  HS65_LH_BFX2 U5877 ( .A(n30353), .Z(n30356) );
  HS65_LH_BFX2 U5878 ( .A(n30360), .Z(n30357) );
  HS65_LH_BFX2 U5879 ( .A(n30361), .Z(n30358) );
  HS65_LH_BFX2 U5880 ( .A(n30356), .Z(n30359) );
  HS65_LH_BFX2 U5881 ( .A(n30363), .Z(n30360) );
  HS65_LH_BFX2 U5882 ( .A(n30364), .Z(n30361) );
  HS65_LH_BFX2 U5883 ( .A(n30359), .Z(n30362) );
  HS65_LH_BFX2 U5884 ( .A(n30366), .Z(n30363) );
  HS65_LH_BFX2 U5885 ( .A(n30367), .Z(n30364) );
  HS65_LH_BFX2 U5886 ( .A(n30362), .Z(n30365) );
  HS65_LH_BFX2 U5887 ( .A(n30371), .Z(n30366) );
  HS65_LH_BFX2 U5888 ( .A(n30370), .Z(n30367) );
  HS65_LH_BFX2 U5889 ( .A(n30365), .Z(n30368) );
  HS65_LH_IVX2 U5890 ( .A(n38798), .Z(n30369) );
  HS65_LH_IVX2 U5891 ( .A(n30369), .Z(n30370) );
  HS65_LH_BFX2 U5892 ( .A(n38771), .Z(n30371) );
  HS65_LH_BFX2 U5893 ( .A(n30464), .Z(n30372) );
  HS65_LH_IVX2 U5894 ( .A(n18078), .Z(n30461) );
  HS65_LH_BFX2 U5895 ( .A(n30378), .Z(n30373) );
  HS65_LH_BFX2 U5896 ( .A(n30376), .Z(n30374) );
  HS65_LH_IVX2 U5897 ( .A(n30381), .Z(n30375) );
  HS65_LH_IVX2 U5898 ( .A(n30375), .Z(n30376) );
  HS65_LH_IVX2 U5899 ( .A(n30383), .Z(n30377) );
  HS65_LH_IVX2 U5900 ( .A(n30377), .Z(n30378) );
  HS65_LH_BFX2 U5901 ( .A(n18076), .Z(n30379) );
  HS65_LH_IVX2 U5902 ( .A(n30386), .Z(n30380) );
  HS65_LH_IVX2 U5903 ( .A(n30380), .Z(n30381) );
  HS65_LH_IVX2 U5904 ( .A(n30388), .Z(n30382) );
  HS65_LH_IVX2 U5905 ( .A(n30382), .Z(n30383) );
  HS65_LH_BFX2 U5906 ( .A(n30379), .Z(n30384) );
  HS65_LH_IVX2 U5907 ( .A(n30391), .Z(n30385) );
  HS65_LH_IVX2 U5908 ( .A(n30385), .Z(n30386) );
  HS65_LH_IVX2 U5909 ( .A(n30393), .Z(n30387) );
  HS65_LH_IVX2 U5910 ( .A(n30387), .Z(n30388) );
  HS65_LH_BFX2 U5911 ( .A(n30384), .Z(n30389) );
  HS65_LH_IVX2 U5912 ( .A(n30396), .Z(n30390) );
  HS65_LH_IVX2 U5913 ( .A(n30390), .Z(n30391) );
  HS65_LH_IVX2 U5914 ( .A(n30398), .Z(n30392) );
  HS65_LH_IVX2 U5915 ( .A(n30392), .Z(n30393) );
  HS65_LH_BFX2 U5917 ( .A(n30389), .Z(n30394) );
  HS65_LH_IVX2 U5919 ( .A(n30401), .Z(n30395) );
  HS65_LH_IVX2 U5921 ( .A(n30395), .Z(n30396) );
  HS65_LH_IVX2 U5923 ( .A(n30403), .Z(n30397) );
  HS65_LH_IVX2 U5925 ( .A(n30397), .Z(n30398) );
  HS65_LH_BFX2 U5927 ( .A(n30394), .Z(n30399) );
  HS65_LH_IVX2 U5929 ( .A(n30407), .Z(n30400) );
  HS65_LH_IVX2 U5931 ( .A(n30400), .Z(n30401) );
  HS65_LH_IVX2 U5937 ( .A(n30409), .Z(n30402) );
  HS65_LH_IVX2 U5938 ( .A(n30402), .Z(n30403) );
  HS65_LH_BFX2 U5939 ( .A(n30399), .Z(n30404) );
  HS65_LH_BFX2 U5940 ( .A(n30404), .Z(n30405) );
  HS65_LH_IVX2 U5941 ( .A(n30412), .Z(n30406) );
  HS65_LH_IVX2 U5942 ( .A(n30406), .Z(n30407) );
  HS65_LH_IVX2 U5943 ( .A(n30414), .Z(n30408) );
  HS65_LH_IVX2 U5944 ( .A(n30408), .Z(n30409) );
  HS65_LH_BFX2 U5945 ( .A(n30405), .Z(n30410) );
  HS65_LH_IVX2 U5946 ( .A(n30417), .Z(n30411) );
  HS65_LH_IVX2 U5947 ( .A(n30411), .Z(n30412) );
  HS65_LH_IVX2 U5948 ( .A(n30419), .Z(n30413) );
  HS65_LH_IVX2 U5949 ( .A(n30413), .Z(n30414) );
  HS65_LH_BFX2 U5950 ( .A(n30410), .Z(n30415) );
  HS65_LH_IVX2 U5951 ( .A(n30422), .Z(n30416) );
  HS65_LH_IVX2 U5952 ( .A(n30416), .Z(n30417) );
  HS65_LH_IVX2 U5953 ( .A(n30424), .Z(n30418) );
  HS65_LH_IVX2 U5954 ( .A(n30418), .Z(n30419) );
  HS65_LH_BFX2 U5955 ( .A(n30415), .Z(n30420) );
  HS65_LH_IVX2 U5956 ( .A(n30427), .Z(n30421) );
  HS65_LH_IVX2 U5957 ( .A(n30421), .Z(n30422) );
  HS65_LH_IVX2 U5958 ( .A(n30429), .Z(n30423) );
  HS65_LH_IVX2 U5959 ( .A(n30423), .Z(n30424) );
  HS65_LH_BFX2 U5960 ( .A(n30420), .Z(n30425) );
  HS65_LH_IVX2 U5961 ( .A(n30432), .Z(n30426) );
  HS65_LH_IVX2 U5962 ( .A(n30426), .Z(n30427) );
  HS65_LH_IVX2 U5963 ( .A(n30434), .Z(n30428) );
  HS65_LH_IVX2 U5964 ( .A(n30428), .Z(n30429) );
  HS65_LH_BFX2 U5965 ( .A(n30425), .Z(n30430) );
  HS65_LH_IVX2 U5966 ( .A(n30437), .Z(n30431) );
  HS65_LH_IVX2 U5967 ( .A(n30431), .Z(n30432) );
  HS65_LH_IVX2 U5968 ( .A(n30439), .Z(n30433) );
  HS65_LH_IVX2 U5969 ( .A(n30433), .Z(n30434) );
  HS65_LH_BFX2 U5970 ( .A(n30430), .Z(n30435) );
  HS65_LH_IVX2 U5971 ( .A(n30442), .Z(n30436) );
  HS65_LH_IVX2 U5972 ( .A(n30436), .Z(n30437) );
  HS65_LH_IVX2 U5973 ( .A(n30444), .Z(n30438) );
  HS65_LH_IVX2 U5974 ( .A(n30438), .Z(n30439) );
  HS65_LH_BFX2 U5976 ( .A(n30435), .Z(n30440) );
  HS65_LH_IVX2 U5977 ( .A(n30447), .Z(n30441) );
  HS65_LH_IVX2 U5978 ( .A(n30441), .Z(n30442) );
  HS65_LH_IVX2 U5979 ( .A(n30449), .Z(n30443) );
  HS65_LH_IVX2 U5980 ( .A(n30443), .Z(n30444) );
  HS65_LH_BFX2 U5981 ( .A(n30440), .Z(n30445) );
  HS65_LH_IVX2 U5982 ( .A(n30452), .Z(n30446) );
  HS65_LH_IVX2 U5983 ( .A(n30446), .Z(n30447) );
  HS65_LH_IVX2 U5984 ( .A(n30454), .Z(n30448) );
  HS65_LH_IVX2 U5985 ( .A(n30448), .Z(n30449) );
  HS65_LH_BFX2 U5986 ( .A(n30445), .Z(n30450) );
  HS65_LH_IVX2 U5987 ( .A(n30459), .Z(n30451) );
  HS65_LH_IVX2 U5988 ( .A(n30451), .Z(n30452) );
  HS65_LH_IVX2 U5989 ( .A(n30457), .Z(n30453) );
  HS65_LH_IVX2 U5990 ( .A(n30453), .Z(n30454) );
  HS65_LH_BFX2 U5991 ( .A(n30450), .Z(n30455) );
  HS65_LH_IVX2 U5992 ( .A(n30462), .Z(n30456) );
  HS65_LH_IVX2 U5993 ( .A(n30456), .Z(n30457) );
  HS65_LH_BFX2 U5994 ( .A(n30455), .Z(n30458) );
  HS65_LH_BFX2 U5995 ( .A(n39294), .Z(n30459) );
  HS65_LH_BFX2 U5996 ( .A(n30458), .Z(n30460) );
  HS65_LH_IVX2 U5997 ( .A(n30461), .Z(n30462) );
  HS65_LH_IVX2 U5998 ( .A(n30460), .Z(n30463) );
  HS65_LH_IVX2 U5999 ( .A(n30463), .Z(n30464) );
  HS65_LH_BFX2 U6000 ( .A(n30468), .Z(n30465) );
  HS65_LH_BFX2 U6001 ( .A(n30469), .Z(n30466) );
  HS65_LH_BFX2 U6002 ( .A(n18069), .Z(n30467) );
  HS65_LH_BFX2 U6003 ( .A(n30471), .Z(n30468) );
  HS65_LH_BFX2 U6004 ( .A(n30472), .Z(n30469) );
  HS65_LH_BFX2 U6005 ( .A(n30467), .Z(n30470) );
  HS65_LH_BFX2 U6006 ( .A(n30474), .Z(n30471) );
  HS65_LH_BFX2 U6007 ( .A(n30475), .Z(n30472) );
  HS65_LH_BFX2 U6008 ( .A(n30470), .Z(n30473) );
  HS65_LH_BFX2 U6009 ( .A(n30477), .Z(n30474) );
  HS65_LH_BFX2 U6010 ( .A(n30478), .Z(n30475) );
  HS65_LH_BFX2 U6011 ( .A(n30473), .Z(n30476) );
  HS65_LH_BFX2 U6012 ( .A(n30480), .Z(n30477) );
  HS65_LH_BFX2 U6013 ( .A(n30481), .Z(n30478) );
  HS65_LH_BFX2 U6014 ( .A(n30476), .Z(n30479) );
  HS65_LH_BFX2 U6015 ( .A(n30483), .Z(n30480) );
  HS65_LH_BFX2 U6016 ( .A(n30484), .Z(n30481) );
  HS65_LH_BFX2 U6017 ( .A(n30479), .Z(n30482) );
  HS65_LH_BFX2 U6018 ( .A(n30486), .Z(n30483) );
  HS65_LH_BFX2 U6019 ( .A(n30487), .Z(n30484) );
  HS65_LH_BFX2 U6020 ( .A(n30482), .Z(n30485) );
  HS65_LH_BFX2 U6021 ( .A(n30489), .Z(n30486) );
  HS65_LH_BFX2 U6022 ( .A(n30490), .Z(n30487) );
  HS65_LH_BFX2 U6023 ( .A(n30485), .Z(n30488) );
  HS65_LH_BFX2 U6024 ( .A(n30492), .Z(n30489) );
  HS65_LH_BFX2 U6025 ( .A(n30493), .Z(n30490) );
  HS65_LH_BFX2 U6026 ( .A(n30488), .Z(n30491) );
  HS65_LH_BFX2 U6027 ( .A(n30495), .Z(n30492) );
  HS65_LH_BFX2 U6028 ( .A(n30496), .Z(n30493) );
  HS65_LH_BFX2 U6029 ( .A(n30491), .Z(n30494) );
  HS65_LH_BFX2 U6030 ( .A(n30498), .Z(n30495) );
  HS65_LH_BFX2 U6031 ( .A(n30499), .Z(n30496) );
  HS65_LH_BFX2 U6032 ( .A(n30494), .Z(n30497) );
  HS65_LH_BFX2 U6035 ( .A(n30501), .Z(n30498) );
  HS65_LH_BFX2 U6036 ( .A(n30502), .Z(n30499) );
  HS65_LH_BFX2 U6037 ( .A(n30497), .Z(n30500) );
  HS65_LH_BFX2 U6038 ( .A(n30504), .Z(n30501) );
  HS65_LH_BFX2 U6039 ( .A(n30505), .Z(n30502) );
  HS65_LH_BFX2 U6040 ( .A(n30500), .Z(n30503) );
  HS65_LH_BFX2 U6041 ( .A(n30507), .Z(n30504) );
  HS65_LH_BFX2 U6042 ( .A(n30508), .Z(n30505) );
  HS65_LH_BFX2 U6043 ( .A(n30503), .Z(n30506) );
  HS65_LH_BFX2 U6044 ( .A(n30510), .Z(n30507) );
  HS65_LH_BFX2 U6045 ( .A(n30511), .Z(n30508) );
  HS65_LH_BFX2 U6046 ( .A(n30506), .Z(n30509) );
  HS65_LH_BFX2 U6047 ( .A(n30513), .Z(n30510) );
  HS65_LH_BFX2 U6048 ( .A(n30514), .Z(n30511) );
  HS65_LH_BFX2 U6049 ( .A(n30509), .Z(n30512) );
  HS65_LH_BFX2 U6050 ( .A(n30516), .Z(n30513) );
  HS65_LH_BFX2 U6051 ( .A(n30517), .Z(n30514) );
  HS65_LH_BFX2 U6052 ( .A(n30512), .Z(n30515) );
  HS65_LH_BFX2 U6053 ( .A(n38750), .Z(n30516) );
  HS65_LH_BFX2 U6054 ( .A(n30520), .Z(n30517) );
  HS65_LH_BFX2 U6055 ( .A(n30515), .Z(n30518) );
  HS65_LH_IVX2 U6056 ( .A(n38812), .Z(n30519) );
  HS65_LH_IVX2 U6057 ( .A(n30519), .Z(n30520) );
  HS65_LH_BFX2 U6058 ( .A(n30524), .Z(n30521) );
  HS65_LH_BFX2 U6059 ( .A(n30525), .Z(n30522) );
  HS65_LH_BFX2 U6060 ( .A(n18079), .Z(n30523) );
  HS65_LH_BFX2 U6061 ( .A(n30527), .Z(n30524) );
  HS65_LH_BFX2 U6062 ( .A(n30528), .Z(n30525) );
  HS65_LH_BFX2 U6063 ( .A(n30523), .Z(n30526) );
  HS65_LH_BFX2 U6064 ( .A(n30530), .Z(n30527) );
  HS65_LH_BFX2 U6065 ( .A(n30531), .Z(n30528) );
  HS65_LH_BFX2 U6066 ( .A(n30526), .Z(n30529) );
  HS65_LH_BFX2 U6067 ( .A(n30533), .Z(n30530) );
  HS65_LH_BFX2 U6068 ( .A(n30534), .Z(n30531) );
  HS65_LH_BFX2 U6069 ( .A(n30529), .Z(n30532) );
  HS65_LH_BFX2 U6070 ( .A(n30536), .Z(n30533) );
  HS65_LH_BFX2 U6071 ( .A(n30537), .Z(n30534) );
  HS65_LH_BFX2 U6072 ( .A(n30532), .Z(n30535) );
  HS65_LH_BFX2 U6073 ( .A(n30539), .Z(n30536) );
  HS65_LH_BFX2 U6074 ( .A(n30540), .Z(n30537) );
  HS65_LH_BFX2 U6075 ( .A(n30535), .Z(n30538) );
  HS65_LH_BFX2 U6076 ( .A(n30542), .Z(n30539) );
  HS65_LH_BFX2 U6077 ( .A(n30543), .Z(n30540) );
  HS65_LH_BFX2 U6078 ( .A(n30538), .Z(n30541) );
  HS65_LH_BFX2 U6079 ( .A(n30545), .Z(n30542) );
  HS65_LH_BFX2 U6080 ( .A(n30546), .Z(n30543) );
  HS65_LH_BFX2 U6081 ( .A(n30541), .Z(n30544) );
  HS65_LH_BFX2 U6082 ( .A(n30548), .Z(n30545) );
  HS65_LH_BFX2 U6083 ( .A(n30549), .Z(n30546) );
  HS65_LH_BFX2 U6084 ( .A(n30544), .Z(n30547) );
  HS65_LH_BFX2 U6085 ( .A(n30551), .Z(n30548) );
  HS65_LH_BFX2 U6086 ( .A(n30552), .Z(n30549) );
  HS65_LH_BFX2 U6087 ( .A(n30547), .Z(n30550) );
  HS65_LH_BFX2 U6088 ( .A(n30554), .Z(n30551) );
  HS65_LH_BFX2 U6089 ( .A(n30555), .Z(n30552) );
  HS65_LH_BFX2 U6090 ( .A(n30550), .Z(n30553) );
  HS65_LH_BFX2 U6091 ( .A(n30557), .Z(n30554) );
  HS65_LH_BFX2 U6092 ( .A(n30558), .Z(n30555) );
  HS65_LH_BFX2 U6093 ( .A(n30553), .Z(n30556) );
  HS65_LH_BFX2 U6094 ( .A(n30560), .Z(n30557) );
  HS65_LH_BFX2 U6095 ( .A(n30561), .Z(n30558) );
  HS65_LH_BFX2 U6096 ( .A(n30556), .Z(n30559) );
  HS65_LH_BFX2 U6097 ( .A(n30563), .Z(n30560) );
  HS65_LH_BFX2 U6098 ( .A(n30564), .Z(n30561) );
  HS65_LH_BFX2 U6099 ( .A(n30559), .Z(n30562) );
  HS65_LH_BFX2 U6100 ( .A(n30566), .Z(n30563) );
  HS65_LH_BFX2 U6101 ( .A(n30567), .Z(n30564) );
  HS65_LH_BFX2 U6102 ( .A(n30562), .Z(n30565) );
  HS65_LH_BFX2 U6103 ( .A(n30569), .Z(n30566) );
  HS65_LH_BFX2 U6104 ( .A(n30570), .Z(n30567) );
  HS65_LH_BFX2 U6105 ( .A(n30565), .Z(n30568) );
  HS65_LH_BFX2 U6106 ( .A(n30572), .Z(n30569) );
  HS65_LH_BFX2 U6107 ( .A(n30573), .Z(n30570) );
  HS65_LH_BFX2 U6109 ( .A(n30568), .Z(n30571) );
  HS65_LH_BFX2 U6110 ( .A(n30575), .Z(n30572) );
  HS65_LH_BFX2 U6111 ( .A(n30576), .Z(n30573) );
  HS65_LH_BFX2 U6112 ( .A(n30571), .Z(n30574) );
  HS65_LH_BFX2 U6113 ( .A(n30582), .Z(n30575) );
  HS65_LH_BFX2 U6114 ( .A(n30579), .Z(n30576) );
  HS65_LH_BFX2 U6115 ( .A(n30574), .Z(n30577) );
  HS65_LH_IVX2 U6116 ( .A(n18080), .Z(n30578) );
  HS65_LH_IVX2 U6117 ( .A(n30578), .Z(n30579) );
  HS65_LH_IVX2 U6118 ( .A(n30577), .Z(n30580) );
  HS65_LH_IVX2 U6119 ( .A(n30580), .Z(n30581) );
  HS65_LH_BFX2 U6120 ( .A(n17678), .Z(n30582) );
  HS65_LH_BFX2 U6121 ( .A(n30586), .Z(n30583) );
  HS65_LH_BFX2 U6122 ( .A(n30587), .Z(n30584) );
  HS65_LH_BFX2 U6123 ( .A(n18074), .Z(n30585) );
  HS65_LH_BFX2 U6124 ( .A(n30589), .Z(n30586) );
  HS65_LH_BFX2 U6125 ( .A(n30590), .Z(n30587) );
  HS65_LH_BFX2 U6126 ( .A(n30585), .Z(n30588) );
  HS65_LH_BFX2 U6127 ( .A(n30592), .Z(n30589) );
  HS65_LH_BFX2 U6128 ( .A(n30593), .Z(n30590) );
  HS65_LH_BFX2 U6129 ( .A(n30588), .Z(n30591) );
  HS65_LH_BFX2 U6130 ( .A(n30595), .Z(n30592) );
  HS65_LH_BFX2 U6131 ( .A(n30596), .Z(n30593) );
  HS65_LH_BFX2 U6132 ( .A(n30591), .Z(n30594) );
  HS65_LH_BFX2 U6133 ( .A(n30598), .Z(n30595) );
  HS65_LH_BFX2 U6134 ( .A(n30599), .Z(n30596) );
  HS65_LH_BFX2 U6135 ( .A(n30594), .Z(n30597) );
  HS65_LH_BFX2 U6136 ( .A(n30601), .Z(n30598) );
  HS65_LH_BFX2 U6137 ( .A(n30602), .Z(n30599) );
  HS65_LH_BFX2 U6138 ( .A(n30597), .Z(n30600) );
  HS65_LH_BFX2 U6139 ( .A(n30604), .Z(n30601) );
  HS65_LH_BFX2 U6140 ( .A(n30605), .Z(n30602) );
  HS65_LH_BFX2 U6141 ( .A(n30600), .Z(n30603) );
  HS65_LH_BFX2 U6142 ( .A(n30607), .Z(n30604) );
  HS65_LH_BFX2 U6143 ( .A(n30608), .Z(n30605) );
  HS65_LH_BFX2 U6144 ( .A(n30603), .Z(n30606) );
  HS65_LH_BFX2 U6145 ( .A(n30610), .Z(n30607) );
  HS65_LH_BFX2 U6146 ( .A(n30611), .Z(n30608) );
  HS65_LH_BFX2 U6147 ( .A(n30606), .Z(n30609) );
  HS65_LH_BFX2 U6148 ( .A(n30613), .Z(n30610) );
  HS65_LH_BFX2 U6149 ( .A(n30614), .Z(n30611) );
  HS65_LH_BFX2 U6150 ( .A(n30609), .Z(n30612) );
  HS65_LH_BFX2 U6151 ( .A(n30616), .Z(n30613) );
  HS65_LH_BFX2 U6152 ( .A(n30617), .Z(n30614) );
  HS65_LH_BFX2 U6153 ( .A(n30612), .Z(n30615) );
  HS65_LH_BFX2 U6154 ( .A(n30619), .Z(n30616) );
  HS65_LH_BFX2 U6155 ( .A(n30620), .Z(n30617) );
  HS65_LH_BFX2 U6160 ( .A(n30615), .Z(n30618) );
  HS65_LH_BFX2 U6161 ( .A(n30622), .Z(n30619) );
  HS65_LH_BFX2 U6162 ( .A(n30623), .Z(n30620) );
  HS65_LH_BFX2 U6164 ( .A(n30618), .Z(n30621) );
  HS65_LH_BFX2 U6165 ( .A(n30625), .Z(n30622) );
  HS65_LH_BFX2 U6166 ( .A(n30626), .Z(n30623) );
  HS65_LH_BFX2 U6168 ( .A(n30621), .Z(n30624) );
  HS65_LH_BFX2 U6170 ( .A(n30628), .Z(n30625) );
  HS65_LH_BFX2 U6172 ( .A(n30629), .Z(n30626) );
  HS65_LH_BFX2 U6178 ( .A(n30624), .Z(n30627) );
  HS65_LH_BFX2 U6179 ( .A(n30631), .Z(n30628) );
  HS65_LH_BFX2 U6180 ( .A(n30632), .Z(n30629) );
  HS65_LH_BFX2 U6181 ( .A(n30627), .Z(n30630) );
  HS65_LH_BFX2 U6182 ( .A(n30634), .Z(n30631) );
  HS65_LH_BFX2 U6183 ( .A(n30635), .Z(n30632) );
  HS65_LH_BFX2 U6184 ( .A(n30630), .Z(n30633) );
  HS65_LH_BFX2 U6185 ( .A(n30637), .Z(n30634) );
  HS65_LH_BFX2 U6186 ( .A(n30638), .Z(n30635) );
  HS65_LH_BFX2 U6187 ( .A(n30633), .Z(n30636) );
  HS65_LH_BFX2 U6188 ( .A(n30644), .Z(n30637) );
  HS65_LH_BFX2 U6189 ( .A(n30641), .Z(n30638) );
  HS65_LH_BFX2 U6190 ( .A(n30636), .Z(n30639) );
  HS65_LH_IVX2 U6191 ( .A(n18075), .Z(n30640) );
  HS65_LH_IVX2 U6192 ( .A(n30640), .Z(n30641) );
  HS65_LH_IVX2 U6193 ( .A(n30639), .Z(n30642) );
  HS65_LH_IVX2 U6194 ( .A(n30642), .Z(n30643) );
  HS65_LH_BFX2 U6195 ( .A(n17674), .Z(n30644) );
  HS65_LH_BFX2 U6196 ( .A(n30737), .Z(n30645) );
  HS65_LH_IVX2 U6197 ( .A(n18084), .Z(n30734) );
  HS65_LH_BFX2 U6198 ( .A(n30651), .Z(n30646) );
  HS65_LH_BFX2 U6199 ( .A(n30649), .Z(n30647) );
  HS65_LH_IVX2 U6200 ( .A(n30654), .Z(n30648) );
  HS65_LH_IVX2 U6201 ( .A(n30648), .Z(n30649) );
  HS65_LH_IVX2 U6202 ( .A(n30656), .Z(n30650) );
  HS65_LH_IVX2 U6203 ( .A(n30650), .Z(n30651) );
  HS65_LH_BFX2 U6204 ( .A(n18083), .Z(n30652) );
  HS65_LH_IVX2 U6205 ( .A(n30659), .Z(n30653) );
  HS65_LH_IVX2 U6206 ( .A(n30653), .Z(n30654) );
  HS65_LH_IVX2 U6207 ( .A(n30661), .Z(n30655) );
  HS65_LH_IVX2 U6208 ( .A(n30655), .Z(n30656) );
  HS65_LH_BFX2 U6209 ( .A(n30652), .Z(n30657) );
  HS65_LH_IVX2 U6210 ( .A(n30664), .Z(n30658) );
  HS65_LH_IVX2 U6211 ( .A(n30658), .Z(n30659) );
  HS65_LH_IVX2 U6212 ( .A(n30666), .Z(n30660) );
  HS65_LH_IVX2 U6213 ( .A(n30660), .Z(n30661) );
  HS65_LH_BFX2 U6214 ( .A(n30657), .Z(n30662) );
  HS65_LH_IVX2 U6215 ( .A(n30669), .Z(n30663) );
  HS65_LH_IVX2 U6216 ( .A(n30663), .Z(n30664) );
  HS65_LH_IVX2 U6217 ( .A(n30671), .Z(n30665) );
  HS65_LH_IVX2 U6218 ( .A(n30665), .Z(n30666) );
  HS65_LH_BFX2 U6219 ( .A(n30662), .Z(n30667) );
  HS65_LH_IVX2 U6220 ( .A(n30674), .Z(n30668) );
  HS65_LH_IVX2 U6221 ( .A(n30668), .Z(n30669) );
  HS65_LH_IVX2 U6222 ( .A(n30676), .Z(n30670) );
  HS65_LH_IVX2 U6223 ( .A(n30670), .Z(n30671) );
  HS65_LH_BFX2 U6224 ( .A(n30667), .Z(n30672) );
  HS65_LH_IVX2 U6225 ( .A(n30680), .Z(n30673) );
  HS65_LH_IVX2 U6226 ( .A(n30673), .Z(n30674) );
  HS65_LH_IVX2 U6227 ( .A(n30682), .Z(n30675) );
  HS65_LH_IVX2 U6228 ( .A(n30675), .Z(n30676) );
  HS65_LH_BFX2 U6229 ( .A(n30672), .Z(n30677) );
  HS65_LH_BFX2 U6230 ( .A(n30677), .Z(n30678) );
  HS65_LH_IVX2 U6231 ( .A(n30685), .Z(n30679) );
  HS65_LH_IVX2 U6232 ( .A(n30679), .Z(n30680) );
  HS65_LH_IVX2 U6233 ( .A(n30687), .Z(n30681) );
  HS65_LH_IVX2 U6234 ( .A(n30681), .Z(n30682) );
  HS65_LH_BFX2 U6235 ( .A(n30678), .Z(n30683) );
  HS65_LH_IVX2 U6236 ( .A(n30690), .Z(n30684) );
  HS65_LH_IVX2 U6237 ( .A(n30684), .Z(n30685) );
  HS65_LH_IVX2 U6238 ( .A(n30692), .Z(n30686) );
  HS65_LH_IVX2 U6239 ( .A(n30686), .Z(n30687) );
  HS65_LH_BFX2 U6240 ( .A(n30683), .Z(n30688) );
  HS65_LH_IVX2 U6241 ( .A(n30695), .Z(n30689) );
  HS65_LH_IVX2 U6242 ( .A(n30689), .Z(n30690) );
  HS65_LH_IVX2 U6243 ( .A(n30697), .Z(n30691) );
  HS65_LH_IVX2 U6244 ( .A(n30691), .Z(n30692) );
  HS65_LH_BFX2 U6245 ( .A(n30688), .Z(n30693) );
  HS65_LH_IVX2 U6246 ( .A(n30700), .Z(n30694) );
  HS65_LH_IVX2 U6247 ( .A(n30694), .Z(n30695) );
  HS65_LH_IVX2 U6248 ( .A(n30702), .Z(n30696) );
  HS65_LH_IVX2 U6249 ( .A(n30696), .Z(n30697) );
  HS65_LH_BFX2 U6250 ( .A(n30693), .Z(n30698) );
  HS65_LH_IVX2 U6251 ( .A(n30705), .Z(n30699) );
  HS65_LH_IVX2 U6252 ( .A(n30699), .Z(n30700) );
  HS65_LH_IVX2 U6253 ( .A(n30707), .Z(n30701) );
  HS65_LH_IVX2 U6254 ( .A(n30701), .Z(n30702) );
  HS65_LH_BFX2 U6255 ( .A(n30698), .Z(n30703) );
  HS65_LH_IVX2 U6256 ( .A(n30710), .Z(n30704) );
  HS65_LH_IVX2 U6257 ( .A(n30704), .Z(n30705) );
  HS65_LH_IVX2 U6258 ( .A(n30712), .Z(n30706) );
  HS65_LH_IVX2 U6259 ( .A(n30706), .Z(n30707) );
  HS65_LH_BFX2 U6260 ( .A(n30703), .Z(n30708) );
  HS65_LH_IVX2 U6261 ( .A(n30715), .Z(n30709) );
  HS65_LH_IVX2 U6262 ( .A(n30709), .Z(n30710) );
  HS65_LH_IVX2 U6263 ( .A(n30717), .Z(n30711) );
  HS65_LH_IVX2 U6264 ( .A(n30711), .Z(n30712) );
  HS65_LH_BFX2 U6265 ( .A(n30708), .Z(n30713) );
  HS65_LH_IVX2 U6266 ( .A(n30720), .Z(n30714) );
  HS65_LH_IVX2 U6267 ( .A(n30714), .Z(n30715) );
  HS65_LH_IVX2 U6268 ( .A(n30722), .Z(n30716) );
  HS65_LH_IVX2 U6269 ( .A(n30716), .Z(n30717) );
  HS65_LH_BFX2 U6270 ( .A(n30713), .Z(n30718) );
  HS65_LH_IVX2 U6271 ( .A(n30725), .Z(n30719) );
  HS65_LH_IVX2 U6272 ( .A(n30719), .Z(n30720) );
  HS65_LH_IVX2 U6273 ( .A(n30727), .Z(n30721) );
  HS65_LH_IVX2 U6274 ( .A(n30721), .Z(n30722) );
  HS65_LH_BFX2 U6275 ( .A(n30718), .Z(n30723) );
  HS65_LH_IVX2 U6276 ( .A(n30732), .Z(n30724) );
  HS65_LH_IVX2 U6277 ( .A(n30724), .Z(n30725) );
  HS65_LH_IVX2 U6278 ( .A(n30730), .Z(n30726) );
  HS65_LH_IVX2 U6279 ( .A(n30726), .Z(n30727) );
  HS65_LH_BFX2 U6280 ( .A(n30723), .Z(n30728) );
  HS65_LH_IVX2 U6281 ( .A(n30735), .Z(n30729) );
  HS65_LH_IVX2 U6282 ( .A(n30729), .Z(n30730) );
  HS65_LH_BFX2 U6283 ( .A(n30728), .Z(n30731) );
  HS65_LH_BFX2 U6284 ( .A(n39296), .Z(n30732) );
  HS65_LH_BFX2 U6285 ( .A(n30731), .Z(n30733) );
  HS65_LH_IVX2 U6286 ( .A(n30734), .Z(n30735) );
  HS65_LH_IVX2 U6287 ( .A(n30733), .Z(n30736) );
  HS65_LH_IVX2 U6288 ( .A(n30736), .Z(n30737) );
  HS65_LH_BFX2 U6289 ( .A(n30743), .Z(n30738) );
  HS65_LH_BFX2 U6290 ( .A(n30741), .Z(n30739) );
  HS65_LH_IVX2 U6291 ( .A(n30746), .Z(n30740) );
  HS65_LH_IVX2 U6292 ( .A(n30740), .Z(n30741) );
  HS65_LH_IVX2 U6293 ( .A(n30748), .Z(n30742) );
  HS65_LH_IVX2 U6294 ( .A(n30742), .Z(n30743) );
  HS65_LH_BFX2 U6295 ( .A(n18087), .Z(n30744) );
  HS65_LH_IVX2 U6296 ( .A(n30751), .Z(n30745) );
  HS65_LH_IVX2 U6297 ( .A(n30745), .Z(n30746) );
  HS65_LH_IVX2 U6298 ( .A(n30753), .Z(n30747) );
  HS65_LH_IVX2 U6299 ( .A(n30747), .Z(n30748) );
  HS65_LH_BFX2 U6300 ( .A(n30744), .Z(n30749) );
  HS65_LH_IVX2 U6301 ( .A(n30756), .Z(n30750) );
  HS65_LH_IVX2 U6302 ( .A(n30750), .Z(n30751) );
  HS65_LH_IVX2 U6303 ( .A(n30758), .Z(n30752) );
  HS65_LH_IVX2 U6304 ( .A(n30752), .Z(n30753) );
  HS65_LH_BFX2 U6305 ( .A(n30749), .Z(n30754) );
  HS65_LH_IVX2 U6306 ( .A(n30761), .Z(n30755) );
  HS65_LH_IVX2 U6308 ( .A(n30755), .Z(n30756) );
  HS65_LH_IVX2 U6309 ( .A(n30763), .Z(n30757) );
  HS65_LH_IVX2 U6310 ( .A(n30757), .Z(n30758) );
  HS65_LH_BFX2 U6311 ( .A(n30754), .Z(n30759) );
  HS65_LH_IVX2 U6312 ( .A(n30766), .Z(n30760) );
  HS65_LH_IVX2 U6313 ( .A(n30760), .Z(n30761) );
  HS65_LH_IVX2 U6314 ( .A(n30768), .Z(n30762) );
  HS65_LH_IVX2 U6315 ( .A(n30762), .Z(n30763) );
  HS65_LH_BFX2 U6316 ( .A(n30759), .Z(n30764) );
  HS65_LH_IVX2 U6317 ( .A(n30772), .Z(n30765) );
  HS65_LH_IVX2 U6318 ( .A(n30765), .Z(n30766) );
  HS65_LH_IVX2 U6319 ( .A(n30774), .Z(n30767) );
  HS65_LH_IVX2 U6320 ( .A(n30767), .Z(n30768) );
  HS65_LH_BFX2 U6321 ( .A(n30764), .Z(n30769) );
  HS65_LH_BFX2 U6322 ( .A(n30769), .Z(n30770) );
  HS65_LH_IVX2 U6323 ( .A(n30777), .Z(n30771) );
  HS65_LH_IVX2 U6324 ( .A(n30771), .Z(n30772) );
  HS65_LH_IVX2 U6325 ( .A(n30779), .Z(n30773) );
  HS65_LH_IVX2 U6326 ( .A(n30773), .Z(n30774) );
  HS65_LH_BFX2 U6327 ( .A(n30770), .Z(n30775) );
  HS65_LH_IVX2 U6328 ( .A(n30782), .Z(n30776) );
  HS65_LH_IVX2 U6329 ( .A(n30776), .Z(n30777) );
  HS65_LH_IVX2 U6330 ( .A(n30784), .Z(n30778) );
  HS65_LH_IVX2 U6331 ( .A(n30778), .Z(n30779) );
  HS65_LH_BFX2 U6332 ( .A(n30775), .Z(n30780) );
  HS65_LH_IVX2 U6333 ( .A(n30787), .Z(n30781) );
  HS65_LH_IVX2 U6334 ( .A(n30781), .Z(n30782) );
  HS65_LH_IVX2 U6335 ( .A(n30789), .Z(n30783) );
  HS65_LH_IVX2 U6336 ( .A(n30783), .Z(n30784) );
  HS65_LH_BFX2 U6337 ( .A(n30780), .Z(n30785) );
  HS65_LH_IVX2 U6338 ( .A(n30792), .Z(n30786) );
  HS65_LH_IVX2 U6339 ( .A(n30786), .Z(n30787) );
  HS65_LH_IVX2 U6340 ( .A(n30794), .Z(n30788) );
  HS65_LH_IVX2 U6341 ( .A(n30788), .Z(n30789) );
  HS65_LH_BFX2 U6342 ( .A(n30785), .Z(n30790) );
  HS65_LH_IVX2 U6343 ( .A(n30797), .Z(n30791) );
  HS65_LH_IVX2 U6344 ( .A(n30791), .Z(n30792) );
  HS65_LH_IVX2 U6345 ( .A(n30799), .Z(n30793) );
  HS65_LH_IVX2 U6346 ( .A(n30793), .Z(n30794) );
  HS65_LH_BFX2 U6347 ( .A(n30790), .Z(n30795) );
  HS65_LH_IVX2 U6348 ( .A(n30802), .Z(n30796) );
  HS65_LH_IVX2 U6349 ( .A(n30796), .Z(n30797) );
  HS65_LH_IVX2 U6350 ( .A(n30804), .Z(n30798) );
  HS65_LH_IVX2 U6351 ( .A(n30798), .Z(n30799) );
  HS65_LH_BFX2 U6352 ( .A(n30795), .Z(n30800) );
  HS65_LH_IVX2 U6353 ( .A(n30807), .Z(n30801) );
  HS65_LH_IVX2 U6354 ( .A(n30801), .Z(n30802) );
  HS65_LH_IVX2 U6355 ( .A(n30809), .Z(n30803) );
  HS65_LH_IVX2 U6356 ( .A(n30803), .Z(n30804) );
  HS65_LH_BFX2 U6357 ( .A(n30800), .Z(n30805) );
  HS65_LH_IVX2 U6358 ( .A(n30812), .Z(n30806) );
  HS65_LH_IVX2 U6359 ( .A(n30806), .Z(n30807) );
  HS65_LH_IVX2 U6360 ( .A(n30814), .Z(n30808) );
  HS65_LH_IVX2 U6361 ( .A(n30808), .Z(n30809) );
  HS65_LH_BFX2 U6362 ( .A(n30805), .Z(n30810) );
  HS65_LH_IVX2 U6363 ( .A(n30819), .Z(n30811) );
  HS65_LH_IVX2 U6364 ( .A(n30811), .Z(n30812) );
  HS65_LH_IVX2 U6365 ( .A(n30817), .Z(n30813) );
  HS65_LH_IVX2 U6366 ( .A(n30813), .Z(n30814) );
  HS65_LH_BFX2 U6367 ( .A(n30810), .Z(n30815) );
  HS65_LH_IVX2 U6368 ( .A(n30824), .Z(n30816) );
  HS65_LH_IVX2 U6369 ( .A(n30816), .Z(n30817) );
  HS65_LH_IVX2 U6370 ( .A(n30822), .Z(n30818) );
  HS65_LH_IVX2 U6372 ( .A(n30818), .Z(n30819) );
  HS65_LH_BFX2 U6373 ( .A(n30815), .Z(n30820) );
  HS65_LH_IVX2 U6374 ( .A(n30827), .Z(n30821) );
  HS65_LH_IVX2 U6375 ( .A(n30821), .Z(n30822) );
  HS65_LH_BFX2 U6376 ( .A(n30820), .Z(n30823) );
  HS65_LH_BFX2 U6377 ( .A(n39295), .Z(n30824) );
  HS65_LH_BFX2 U6378 ( .A(n30823), .Z(n30825) );
  HS65_LH_IVX2 U6379 ( .A(n18088), .Z(n30826) );
  HS65_LH_IVX2 U6380 ( .A(n30826), .Z(n30827) );
  HS65_LH_IVX2 U6381 ( .A(n30825), .Z(n30828) );
  HS65_LH_IVX2 U6382 ( .A(n30828), .Z(n30829) );
  HS65_LH_BFX2 U6383 ( .A(n30833), .Z(n30830) );
  HS65_LH_BFX2 U6384 ( .A(n30834), .Z(n30831) );
  HS65_LH_BFX2 U6385 ( .A(n18017), .Z(n30832) );
  HS65_LH_BFX2 U6386 ( .A(n30836), .Z(n30833) );
  HS65_LH_BFX2 U6387 ( .A(n30837), .Z(n30834) );
  HS65_LH_BFX2 U6388 ( .A(n30832), .Z(n30835) );
  HS65_LH_BFX2 U6389 ( .A(n30839), .Z(n30836) );
  HS65_LH_BFX2 U6390 ( .A(n30840), .Z(n30837) );
  HS65_LH_BFX2 U6391 ( .A(n30835), .Z(n30838) );
  HS65_LH_BFX2 U6392 ( .A(n30842), .Z(n30839) );
  HS65_LH_BFX2 U6393 ( .A(n30843), .Z(n30840) );
  HS65_LH_BFX2 U6394 ( .A(n30838), .Z(n30841) );
  HS65_LH_BFX2 U6395 ( .A(n30845), .Z(n30842) );
  HS65_LH_BFX2 U6396 ( .A(n30846), .Z(n30843) );
  HS65_LH_BFX2 U6397 ( .A(n30841), .Z(n30844) );
  HS65_LH_BFX2 U6398 ( .A(n30848), .Z(n30845) );
  HS65_LH_BFX2 U6399 ( .A(n30849), .Z(n30846) );
  HS65_LH_BFX2 U6400 ( .A(n30844), .Z(n30847) );
  HS65_LH_BFX2 U6401 ( .A(n30851), .Z(n30848) );
  HS65_LH_BFX2 U6402 ( .A(n30852), .Z(n30849) );
  HS65_LH_BFX2 U6403 ( .A(n30847), .Z(n30850) );
  HS65_LH_BFX2 U6404 ( .A(n30854), .Z(n30851) );
  HS65_LH_BFX2 U6405 ( .A(n30855), .Z(n30852) );
  HS65_LH_BFX2 U6406 ( .A(n30850), .Z(n30853) );
  HS65_LH_BFX2 U6407 ( .A(n30857), .Z(n30854) );
  HS65_LH_BFX2 U6408 ( .A(n30858), .Z(n30855) );
  HS65_LH_BFX2 U6409 ( .A(n30853), .Z(n30856) );
  HS65_LH_BFX2 U6410 ( .A(n30860), .Z(n30857) );
  HS65_LH_BFX2 U6411 ( .A(n30861), .Z(n30858) );
  HS65_LH_BFX2 U6412 ( .A(n30856), .Z(n30859) );
  HS65_LH_BFX2 U6413 ( .A(n30863), .Z(n30860) );
  HS65_LH_BFX2 U6414 ( .A(n30864), .Z(n30861) );
  HS65_LH_BFX2 U6415 ( .A(n30859), .Z(n30862) );
  HS65_LH_BFX2 U6416 ( .A(n30866), .Z(n30863) );
  HS65_LH_BFX2 U6417 ( .A(n30867), .Z(n30864) );
  HS65_LH_BFX2 U6418 ( .A(n30862), .Z(n30865) );
  HS65_LH_BFX2 U6419 ( .A(n30869), .Z(n30866) );
  HS65_LH_BFX2 U6420 ( .A(n30870), .Z(n30867) );
  HS65_LH_BFX2 U6421 ( .A(n30865), .Z(n30868) );
  HS65_LH_BFX2 U6422 ( .A(n30872), .Z(n30869) );
  HS65_LH_BFX2 U6423 ( .A(n30873), .Z(n30870) );
  HS65_LH_BFX2 U6424 ( .A(n30868), .Z(n30871) );
  HS65_LH_BFX2 U6425 ( .A(n30875), .Z(n30872) );
  HS65_LH_BFX2 U6426 ( .A(n30876), .Z(n30873) );
  HS65_LH_BFX2 U6427 ( .A(n30871), .Z(n30874) );
  HS65_LH_BFX2 U6428 ( .A(n30878), .Z(n30875) );
  HS65_LH_BFX2 U6429 ( .A(n30879), .Z(n30876) );
  HS65_LH_BFX2 U6430 ( .A(n30874), .Z(n30877) );
  HS65_LH_BFX2 U6431 ( .A(n30881), .Z(n30878) );
  HS65_LH_BFX2 U6432 ( .A(n30882), .Z(n30879) );
  HS65_LH_BFX2 U6433 ( .A(n30877), .Z(n30880) );
  HS65_LH_BFX2 U6434 ( .A(n30884), .Z(n30881) );
  HS65_LH_BFX2 U6435 ( .A(n30885), .Z(n30882) );
  HS65_LH_BFX2 U6436 ( .A(n30880), .Z(n30883) );
  HS65_LH_BFX2 U6437 ( .A(n30891), .Z(n30884) );
  HS65_LH_BFX2 U6438 ( .A(n30888), .Z(n30885) );
  HS65_LH_BFX2 U6439 ( .A(n30883), .Z(n30886) );
  HS65_LH_IVX2 U6440 ( .A(n18018), .Z(n30887) );
  HS65_LH_IVX2 U6441 ( .A(n30887), .Z(n30888) );
  HS65_LH_IVX2 U6442 ( .A(n30886), .Z(n30889) );
  HS65_LH_IVX2 U6443 ( .A(n30889), .Z(n30890) );
  HS65_LH_BFX2 U6444 ( .A(n17682), .Z(n30891) );
  HS65_LH_IVX2 U6445 ( .A(n36977), .Z(n30892) );
  HS65_LH_IVX2 U6446 ( .A(n30892), .Z(n30893) );
  HS65_LH_BFX2 U6447 ( .A(n30896), .Z(n30894) );
  HS65_LH_BFX2 U6448 ( .A(n18040), .Z(n30895) );
  HS65_LH_BFX2 U6449 ( .A(n36978), .Z(n30896) );
  HS65_LH_BFX2 U6450 ( .A(n30895), .Z(n30897) );
  HS65_LH_BFX2 U6451 ( .A(n30901), .Z(n30898) );
  HS65_LH_BFX2 U6452 ( .A(n30903), .Z(n30899) );
  HS65_LH_IVX2 U6453 ( .A(n30906), .Z(n30900) );
  HS65_LH_IVX2 U6454 ( .A(n30900), .Z(n30901) );
  HS65_LH_IVX2 U6455 ( .A(n30908), .Z(n30902) );
  HS65_LH_IVX2 U6456 ( .A(n30902), .Z(n30903) );
  HS65_LH_BFX2 U6457 ( .A(n18019), .Z(n30904) );
  HS65_LH_IVX2 U6458 ( .A(n30911), .Z(n30905) );
  HS65_LH_IVX2 U6459 ( .A(n30905), .Z(n30906) );
  HS65_LH_IVX2 U6460 ( .A(n30914), .Z(n30907) );
  HS65_LH_IVX2 U6461 ( .A(n30907), .Z(n30908) );
  HS65_LH_BFX2 U6462 ( .A(n30904), .Z(n30909) );
  HS65_LH_IVX2 U6463 ( .A(n30917), .Z(n30910) );
  HS65_LH_IVX2 U6464 ( .A(n30910), .Z(n30911) );
  HS65_LH_BFX2 U6465 ( .A(n30909), .Z(n30912) );
  HS65_LH_IVX2 U6466 ( .A(n30919), .Z(n30913) );
  HS65_LH_IVX2 U6467 ( .A(n30913), .Z(n30914) );
  HS65_LH_BFX2 U6468 ( .A(n30912), .Z(n30915) );
  HS65_LH_IVX2 U6469 ( .A(n30922), .Z(n30916) );
  HS65_LH_IVX2 U6470 ( .A(n30916), .Z(n30917) );
  HS65_LH_IVX2 U6471 ( .A(n30924), .Z(n30918) );
  HS65_LH_IVX2 U6472 ( .A(n30918), .Z(n30919) );
  HS65_LH_BFX2 U6473 ( .A(n30915), .Z(n30920) );
  HS65_LH_IVX2 U6474 ( .A(n30927), .Z(n30921) );
  HS65_LH_IVX2 U6475 ( .A(n30921), .Z(n30922) );
  HS65_LH_IVX2 U6476 ( .A(n30929), .Z(n30923) );
  HS65_LH_IVX2 U6477 ( .A(n30923), .Z(n30924) );
  HS65_LH_BFX2 U6478 ( .A(n30920), .Z(n30925) );
  HS65_LH_IVX2 U6479 ( .A(n30932), .Z(n30926) );
  HS65_LH_IVX2 U6480 ( .A(n30926), .Z(n30927) );
  HS65_LH_IVX2 U6481 ( .A(n30934), .Z(n30928) );
  HS65_LH_IVX2 U6482 ( .A(n30928), .Z(n30929) );
  HS65_LH_BFX2 U6483 ( .A(n30925), .Z(n30930) );
  HS65_LH_IVX2 U6484 ( .A(n30937), .Z(n30931) );
  HS65_LH_IVX2 U6485 ( .A(n30931), .Z(n30932) );
  HS65_LH_IVX2 U6486 ( .A(n30939), .Z(n30933) );
  HS65_LH_IVX2 U6487 ( .A(n30933), .Z(n30934) );
  HS65_LH_BFX2 U6488 ( .A(n30930), .Z(n30935) );
  HS65_LH_IVX2 U6489 ( .A(n30942), .Z(n30936) );
  HS65_LH_IVX2 U6490 ( .A(n30936), .Z(n30937) );
  HS65_LH_IVX2 U6491 ( .A(n30944), .Z(n30938) );
  HS65_LH_IVX2 U6492 ( .A(n30938), .Z(n30939) );
  HS65_LH_BFX2 U6493 ( .A(n30935), .Z(n30940) );
  HS65_LH_IVX2 U6494 ( .A(n30947), .Z(n30941) );
  HS65_LH_IVX2 U6495 ( .A(n30941), .Z(n30942) );
  HS65_LH_IVX2 U6496 ( .A(n30949), .Z(n30943) );
  HS65_LH_IVX2 U6497 ( .A(n30943), .Z(n30944) );
  HS65_LH_BFX2 U6498 ( .A(n30940), .Z(n30945) );
  HS65_LH_IVX2 U6499 ( .A(n30952), .Z(n30946) );
  HS65_LH_IVX2 U6500 ( .A(n30946), .Z(n30947) );
  HS65_LH_IVX2 U6501 ( .A(n30954), .Z(n30948) );
  HS65_LH_IVX2 U6502 ( .A(n30948), .Z(n30949) );
  HS65_LH_BFX2 U6504 ( .A(n30945), .Z(n30950) );
  HS65_LH_IVX2 U6505 ( .A(n30957), .Z(n30951) );
  HS65_LH_IVX2 U6506 ( .A(n30951), .Z(n30952) );
  HS65_LH_IVX2 U6507 ( .A(n30959), .Z(n30953) );
  HS65_LH_IVX2 U6508 ( .A(n30953), .Z(n30954) );
  HS65_LH_BFX2 U6509 ( .A(n30950), .Z(n30955) );
  HS65_LH_IVX2 U6510 ( .A(n30962), .Z(n30956) );
  HS65_LH_IVX2 U6511 ( .A(n30956), .Z(n30957) );
  HS65_LH_IVX2 U6512 ( .A(n30964), .Z(n30958) );
  HS65_LH_IVX2 U6513 ( .A(n30958), .Z(n30959) );
  HS65_LH_BFX2 U6514 ( .A(n30955), .Z(n30960) );
  HS65_LH_IVX2 U6515 ( .A(n30967), .Z(n30961) );
  HS65_LH_IVX2 U6516 ( .A(n30961), .Z(n30962) );
  HS65_LH_IVX2 U6517 ( .A(n30969), .Z(n30963) );
  HS65_LH_IVX2 U6518 ( .A(n30963), .Z(n30964) );
  HS65_LH_BFX2 U6519 ( .A(n30960), .Z(n30965) );
  HS65_LH_IVX2 U6520 ( .A(n30974), .Z(n30966) );
  HS65_LH_IVX2 U6521 ( .A(n30966), .Z(n30967) );
  HS65_LH_IVX2 U6522 ( .A(n30973), .Z(n30968) );
  HS65_LH_IVX2 U6523 ( .A(n30968), .Z(n30969) );
  HS65_LH_BFX2 U6524 ( .A(n30965), .Z(n30970) );
  HS65_LH_BFX2 U6525 ( .A(n30970), .Z(n30971) );
  HS65_LH_IVX2 U6526 ( .A(n30977), .Z(n30972) );
  HS65_LH_IVX2 U6527 ( .A(n30972), .Z(n30973) );
  HS65_LH_BFX2 U6528 ( .A(n30978), .Z(n30974) );
  HS65_LH_BFX2 U6529 ( .A(n30971), .Z(n30975) );
  HS65_LH_IVX2 U6530 ( .A(n14109), .Z(n30976) );
  HS65_LH_IVX2 U6531 ( .A(n30976), .Z(n30977) );
  HS65_LH_BFX2 U6532 ( .A(n30980), .Z(n30978) );
  HS65_LH_BFX2 U6533 ( .A(n30975), .Z(n30979) );
  HS65_LH_BFX2 U6534 ( .A(n30983), .Z(n30980) );
  HS65_LH_BFX2 U6535 ( .A(n30979), .Z(n30981) );
  HS65_LH_IVX2 U6536 ( .A(n18020), .Z(n30982) );
  HS65_LH_IVX2 U6537 ( .A(n30982), .Z(n30983) );
  HS65_LH_IVX2 U6538 ( .A(n30981), .Z(n30984) );
  HS65_LH_IVX2 U6539 ( .A(n30984), .Z(n30985) );
  HS65_LH_BFX2 U6540 ( .A(n30989), .Z(n30986) );
  HS65_LH_BFX2 U6541 ( .A(n30990), .Z(n30987) );
  HS65_LH_BFX2 U6542 ( .A(n18025), .Z(n30988) );
  HS65_LH_BFX2 U6543 ( .A(n30992), .Z(n30989) );
  HS65_LH_BFX2 U6544 ( .A(n30993), .Z(n30990) );
  HS65_LH_BFX2 U6545 ( .A(n30988), .Z(n30991) );
  HS65_LH_BFX2 U6546 ( .A(n30995), .Z(n30992) );
  HS65_LH_BFX2 U6547 ( .A(n30996), .Z(n30993) );
  HS65_LH_BFX2 U6548 ( .A(n30991), .Z(n30994) );
  HS65_LH_BFX2 U6549 ( .A(n30998), .Z(n30995) );
  HS65_LH_BFX2 U6550 ( .A(n30999), .Z(n30996) );
  HS65_LH_BFX2 U6551 ( .A(n30994), .Z(n30997) );
  HS65_LH_BFX2 U6552 ( .A(n31001), .Z(n30998) );
  HS65_LH_BFX2 U6553 ( .A(n31002), .Z(n30999) );
  HS65_LH_BFX2 U6554 ( .A(n30997), .Z(n31000) );
  HS65_LH_BFX2 U6555 ( .A(n31004), .Z(n31001) );
  HS65_LH_BFX2 U6556 ( .A(n31005), .Z(n31002) );
  HS65_LH_BFX2 U6557 ( .A(n31000), .Z(n31003) );
  HS65_LH_BFX2 U6558 ( .A(n31007), .Z(n31004) );
  HS65_LH_BFX2 U6559 ( .A(n31008), .Z(n31005) );
  HS65_LH_BFX2 U6560 ( .A(n31003), .Z(n31006) );
  HS65_LH_BFX2 U6561 ( .A(n31010), .Z(n31007) );
  HS65_LH_BFX2 U6562 ( .A(n31011), .Z(n31008) );
  HS65_LH_BFX2 U6563 ( .A(n31006), .Z(n31009) );
  HS65_LH_BFX2 U6564 ( .A(n31013), .Z(n31010) );
  HS65_LH_BFX2 U6565 ( .A(n31014), .Z(n31011) );
  HS65_LH_BFX2 U6566 ( .A(n31009), .Z(n31012) );
  HS65_LH_BFX2 U6567 ( .A(n31016), .Z(n31013) );
  HS65_LH_BFX2 U6568 ( .A(n31017), .Z(n31014) );
  HS65_LH_BFX2 U6570 ( .A(n31012), .Z(n31015) );
  HS65_LH_BFX2 U6571 ( .A(n31019), .Z(n31016) );
  HS65_LH_BFX2 U6572 ( .A(n31020), .Z(n31017) );
  HS65_LH_BFX2 U6573 ( .A(n31015), .Z(n31018) );
  HS65_LH_BFX2 U6574 ( .A(n31022), .Z(n31019) );
  HS65_LH_BFX2 U6575 ( .A(n31023), .Z(n31020) );
  HS65_LH_BFX2 U6576 ( .A(n31018), .Z(n31021) );
  HS65_LH_BFX2 U6577 ( .A(n31025), .Z(n31022) );
  HS65_LH_BFX2 U6578 ( .A(n31026), .Z(n31023) );
  HS65_LH_BFX2 U6579 ( .A(n31021), .Z(n31024) );
  HS65_LH_BFX2 U6580 ( .A(n31028), .Z(n31025) );
  HS65_LH_BFX2 U6581 ( .A(n31029), .Z(n31026) );
  HS65_LH_BFX2 U6582 ( .A(n31024), .Z(n31027) );
  HS65_LH_BFX2 U6583 ( .A(n31031), .Z(n31028) );
  HS65_LH_BFX2 U6584 ( .A(n31032), .Z(n31029) );
  HS65_LH_BFX2 U6585 ( .A(n31027), .Z(n31030) );
  HS65_LH_BFX2 U6586 ( .A(n31034), .Z(n31031) );
  HS65_LH_BFX2 U6587 ( .A(n31035), .Z(n31032) );
  HS65_LH_BFX2 U6588 ( .A(n31030), .Z(n31033) );
  HS65_LH_BFX2 U6589 ( .A(n31037), .Z(n31034) );
  HS65_LH_BFX2 U6590 ( .A(n31038), .Z(n31035) );
  HS65_LH_BFX2 U6591 ( .A(n31033), .Z(n31036) );
  HS65_LH_BFX2 U6592 ( .A(n31040), .Z(n31037) );
  HS65_LH_BFX2 U6593 ( .A(n31041), .Z(n31038) );
  HS65_LH_BFX2 U6594 ( .A(n31036), .Z(n31039) );
  HS65_LH_BFX2 U6595 ( .A(n31043), .Z(n31040) );
  HS65_LH_BFX2 U6596 ( .A(n31044), .Z(n31041) );
  HS65_LH_BFX2 U6597 ( .A(n31039), .Z(n31042) );
  HS65_LH_BFX2 U6598 ( .A(n14105), .Z(n31043) );
  HS65_LH_BFX2 U6599 ( .A(n31047), .Z(n31044) );
  HS65_LH_BFX2 U6600 ( .A(n31042), .Z(n31045) );
  HS65_LH_IVX2 U6601 ( .A(n18026), .Z(n31046) );
  HS65_LH_IVX2 U6602 ( .A(n31046), .Z(n31047) );
  HS65_LH_IVX2 U6603 ( .A(n31045), .Z(n31048) );
  HS65_LH_IVX2 U6604 ( .A(n31048), .Z(n31049) );
  HS65_LH_BFX2 U6605 ( .A(n31053), .Z(n31050) );
  HS65_LH_BFX2 U6606 ( .A(n31054), .Z(n31051) );
  HS65_LH_BFX2 U6607 ( .A(n18030), .Z(n31052) );
  HS65_LH_BFX2 U6608 ( .A(n31056), .Z(n31053) );
  HS65_LH_BFX2 U6609 ( .A(n31057), .Z(n31054) );
  HS65_LH_BFX2 U6610 ( .A(n31052), .Z(n31055) );
  HS65_LH_BFX2 U6611 ( .A(n31059), .Z(n31056) );
  HS65_LH_BFX2 U6612 ( .A(n31060), .Z(n31057) );
  HS65_LH_BFX2 U6613 ( .A(n31055), .Z(n31058) );
  HS65_LH_BFX2 U6614 ( .A(n31062), .Z(n31059) );
  HS65_LH_BFX2 U6615 ( .A(n31063), .Z(n31060) );
  HS65_LH_BFX2 U6616 ( .A(n31058), .Z(n31061) );
  HS65_LH_BFX2 U6617 ( .A(n31065), .Z(n31062) );
  HS65_LH_BFX2 U6618 ( .A(n31066), .Z(n31063) );
  HS65_LH_BFX2 U6619 ( .A(n31061), .Z(n31064) );
  HS65_LH_BFX2 U6620 ( .A(n31068), .Z(n31065) );
  HS65_LH_BFX2 U6621 ( .A(n31069), .Z(n31066) );
  HS65_LH_BFX2 U6622 ( .A(n31064), .Z(n31067) );
  HS65_LH_BFX2 U6623 ( .A(n31071), .Z(n31068) );
  HS65_LH_BFX2 U6624 ( .A(n31072), .Z(n31069) );
  HS65_LH_BFX2 U6625 ( .A(n31067), .Z(n31070) );
  HS65_LH_BFX2 U6626 ( .A(n31074), .Z(n31071) );
  HS65_LH_BFX2 U6627 ( .A(n31075), .Z(n31072) );
  HS65_LH_BFX2 U6628 ( .A(n31070), .Z(n31073) );
  HS65_LH_BFX2 U6629 ( .A(n31077), .Z(n31074) );
  HS65_LH_BFX2 U6630 ( .A(n31078), .Z(n31075) );
  HS65_LH_BFX2 U6631 ( .A(n31073), .Z(n31076) );
  HS65_LH_BFX2 U6632 ( .A(n31080), .Z(n31077) );
  HS65_LH_BFX2 U6633 ( .A(n31081), .Z(n31078) );
  HS65_LH_BFX2 U6634 ( .A(n31076), .Z(n31079) );
  HS65_LH_BFX2 U6636 ( .A(n31083), .Z(n31080) );
  HS65_LH_BFX2 U6637 ( .A(n31084), .Z(n31081) );
  HS65_LH_BFX2 U6638 ( .A(n31079), .Z(n31082) );
  HS65_LH_BFX2 U6639 ( .A(n31086), .Z(n31083) );
  HS65_LH_BFX2 U6640 ( .A(n31087), .Z(n31084) );
  HS65_LH_BFX2 U6641 ( .A(n31082), .Z(n31085) );
  HS65_LH_BFX2 U6642 ( .A(n31089), .Z(n31086) );
  HS65_LH_BFX2 U6643 ( .A(n31090), .Z(n31087) );
  HS65_LH_BFX2 U6644 ( .A(n31085), .Z(n31088) );
  HS65_LH_BFX2 U6645 ( .A(n31092), .Z(n31089) );
  HS65_LH_BFX2 U6646 ( .A(n31093), .Z(n31090) );
  HS65_LH_BFX2 U6647 ( .A(n31088), .Z(n31091) );
  HS65_LH_BFX2 U6648 ( .A(n31095), .Z(n31092) );
  HS65_LH_BFX2 U6649 ( .A(n31096), .Z(n31093) );
  HS65_LH_BFX2 U6650 ( .A(n31091), .Z(n31094) );
  HS65_LH_BFX2 U6651 ( .A(n31098), .Z(n31095) );
  HS65_LH_BFX2 U6652 ( .A(n31099), .Z(n31096) );
  HS65_LH_BFX2 U6653 ( .A(n31094), .Z(n31097) );
  HS65_LH_BFX2 U6654 ( .A(n31101), .Z(n31098) );
  HS65_LH_BFX2 U6655 ( .A(n31102), .Z(n31099) );
  HS65_LH_BFX2 U6656 ( .A(n31097), .Z(n31100) );
  HS65_LH_BFX2 U6657 ( .A(n31104), .Z(n31101) );
  HS65_LH_BFX2 U6658 ( .A(n31105), .Z(n31102) );
  HS65_LH_BFX2 U6659 ( .A(n31100), .Z(n31103) );
  HS65_LH_BFX2 U6660 ( .A(n31107), .Z(n31104) );
  HS65_LH_BFX2 U6661 ( .A(n31108), .Z(n31105) );
  HS65_LH_BFX2 U6662 ( .A(n31103), .Z(n31106) );
  HS65_LH_BFX2 U6663 ( .A(n14103), .Z(n31107) );
  HS65_LH_BFX2 U6664 ( .A(n31111), .Z(n31108) );
  HS65_LH_BFX2 U6665 ( .A(n31106), .Z(n31109) );
  HS65_LH_IVX2 U6666 ( .A(n18031), .Z(n31110) );
  HS65_LH_IVX2 U6667 ( .A(n31110), .Z(n31111) );
  HS65_LH_IVX2 U6668 ( .A(n31109), .Z(n31112) );
  HS65_LH_IVX2 U6669 ( .A(n31112), .Z(n31113) );
  HS65_LH_BFX2 U6670 ( .A(n39526), .Z(n31114) );
  HS65_LH_BFX2 U6671 ( .A(n31118), .Z(n31115) );
  HS65_LH_BFX2 U6672 ( .A(n31119), .Z(n31116) );
  HS65_LH_BFX2 U6673 ( .A(n18035), .Z(n31117) );
  HS65_LH_BFX2 U6674 ( .A(n31121), .Z(n31118) );
  HS65_LH_BFX2 U6675 ( .A(n31122), .Z(n31119) );
  HS65_LH_BFX2 U6676 ( .A(n31117), .Z(n31120) );
  HS65_LH_BFX2 U6677 ( .A(n31124), .Z(n31121) );
  HS65_LH_BFX2 U6678 ( .A(n31125), .Z(n31122) );
  HS65_LH_BFX2 U6679 ( .A(n31120), .Z(n31123) );
  HS65_LH_BFX2 U6680 ( .A(n31127), .Z(n31124) );
  HS65_LH_BFX2 U6681 ( .A(n31128), .Z(n31125) );
  HS65_LH_BFX2 U6682 ( .A(n31123), .Z(n31126) );
  HS65_LH_BFX2 U6683 ( .A(n31130), .Z(n31127) );
  HS65_LH_BFX2 U6684 ( .A(n31131), .Z(n31128) );
  HS65_LH_BFX2 U6685 ( .A(n31126), .Z(n31129) );
  HS65_LH_BFX2 U6686 ( .A(n31133), .Z(n31130) );
  HS65_LH_BFX2 U6687 ( .A(n31134), .Z(n31131) );
  HS65_LH_BFX2 U6688 ( .A(n31129), .Z(n31132) );
  HS65_LH_BFX2 U6689 ( .A(n31136), .Z(n31133) );
  HS65_LH_BFX2 U6690 ( .A(n31137), .Z(n31134) );
  HS65_LH_BFX2 U6691 ( .A(n31132), .Z(n31135) );
  HS65_LH_BFX2 U6692 ( .A(n31139), .Z(n31136) );
  HS65_LH_BFX2 U6693 ( .A(n31140), .Z(n31137) );
  HS65_LH_BFX2 U6694 ( .A(n31135), .Z(n31138) );
  HS65_LH_BFX2 U6695 ( .A(n31142), .Z(n31139) );
  HS65_LH_BFX2 U6696 ( .A(n31143), .Z(n31140) );
  HS65_LH_BFX2 U6697 ( .A(n31138), .Z(n31141) );
  HS65_LH_BFX2 U6698 ( .A(n31145), .Z(n31142) );
  HS65_LH_BFX2 U6699 ( .A(n31146), .Z(n31143) );
  HS65_LH_BFX2 U6700 ( .A(n31141), .Z(n31144) );
  HS65_LH_BFX2 U6702 ( .A(n31148), .Z(n31145) );
  HS65_LH_BFX2 U6703 ( .A(n31149), .Z(n31146) );
  HS65_LH_BFX2 U6704 ( .A(n31144), .Z(n31147) );
  HS65_LH_BFX2 U6725 ( .A(n31151), .Z(n31148) );
  HS65_LH_BFX2 U6726 ( .A(n31152), .Z(n31149) );
  HS65_LH_BFX2 U6727 ( .A(n31147), .Z(n31150) );
  HS65_LH_BFX2 U6728 ( .A(n31154), .Z(n31151) );
  HS65_LH_BFX2 U6729 ( .A(n31155), .Z(n31152) );
  HS65_LH_BFX2 U6730 ( .A(n31150), .Z(n31153) );
  HS65_LH_BFX2 U6731 ( .A(n31157), .Z(n31154) );
  HS65_LH_BFX2 U6732 ( .A(n31158), .Z(n31155) );
  HS65_LH_BFX2 U6733 ( .A(n31153), .Z(n31156) );
  HS65_LH_BFX2 U6734 ( .A(n31160), .Z(n31157) );
  HS65_LH_BFX2 U6735 ( .A(n31161), .Z(n31158) );
  HS65_LH_BFX2 U6736 ( .A(n31156), .Z(n31159) );
  HS65_LH_BFX2 U6737 ( .A(n31163), .Z(n31160) );
  HS65_LH_BFX2 U6738 ( .A(n31164), .Z(n31161) );
  HS65_LH_BFX2 U6739 ( .A(n31159), .Z(n31162) );
  HS65_LH_BFX2 U6740 ( .A(n31166), .Z(n31163) );
  HS65_LH_BFX2 U6741 ( .A(n31167), .Z(n31164) );
  HS65_LH_BFX2 U6742 ( .A(n31162), .Z(n31165) );
  HS65_LH_BFX2 U6743 ( .A(n31169), .Z(n31166) );
  HS65_LH_BFX2 U6744 ( .A(n31170), .Z(n31167) );
  HS65_LH_BFX2 U6745 ( .A(n31165), .Z(n31168) );
  HS65_LH_BFX2 U6746 ( .A(n31172), .Z(n31169) );
  HS65_LH_BFX2 U6747 ( .A(n31173), .Z(n31170) );
  HS65_LH_BFX2 U6748 ( .A(n31168), .Z(n31171) );
  HS65_LH_BFX2 U6749 ( .A(n14101), .Z(n31172) );
  HS65_LH_BFX2 U6751 ( .A(n31176), .Z(n31173) );
  HS65_LH_BFX2 U6752 ( .A(n31171), .Z(n31174) );
  HS65_LH_IVX2 U6754 ( .A(n18036), .Z(n31175) );
  HS65_LH_IVX2 U6755 ( .A(n31175), .Z(n31176) );
  HS65_LH_IVX2 U6757 ( .A(n31174), .Z(n31177) );
  HS65_LH_IVX2 U6760 ( .A(n31177), .Z(n31178) );
  HS65_LH_IVX2 U6761 ( .A(n31201), .Z(n31179) );
  HS65_LH_IVX2 U6763 ( .A(n31179), .Z(n31180) );
  HS65_LH_IVX2 U6764 ( .A(n31203), .Z(n31181) );
  HS65_LH_IVX2 U6766 ( .A(n31181), .Z(n31182) );
  HS65_LH_IVX2 U6767 ( .A(n31205), .Z(n31183) );
  HS65_LH_IVX2 U6769 ( .A(n31183), .Z(n31184) );
  HS65_LH_AOI12X2 U6770 ( .A(n17305), .B(n17567), .C(n17434), .Z(n270) );
  HS65_LH_BFX2 U6772 ( .A(n35420), .Z(n31185) );
  HS65_LH_IVX2 U6773 ( .A(n31208), .Z(n31186) );
  HS65_LH_IVX2 U6775 ( .A(n31186), .Z(n31187) );
  HS65_LH_BFX2 U6776 ( .A(n31192), .Z(n31188) );
  HS65_LH_BFX2 U6778 ( .A(n31194), .Z(n31189) );
  HS65_LH_BFX2 U6779 ( .A(n31196), .Z(n31190) );
  HS65_LH_IVX2 U6781 ( .A(n35229), .Z(n31191) );
  HS65_LH_IVX2 U6782 ( .A(n31191), .Z(n31192) );
  HS65_LH_IVX2 U6784 ( .A(n35654), .Z(n31193) );
  HS65_LH_IVX2 U6785 ( .A(n31193), .Z(n31194) );
  HS65_LH_IVX2 U6787 ( .A(n35263), .Z(n31195) );
  HS65_LH_IVX2 U6788 ( .A(n31195), .Z(n31196) );
  HS65_LH_BFX2 U6790 ( .A(n17373), .Z(n31197) );
  HS65_LH_IVX2 U6791 ( .A(n35224), .Z(n31198) );
  HS65_LH_IVX2 U6793 ( .A(n31198), .Z(n31199) );
  HS65_LH_IVX2 U6794 ( .A(n35237), .Z(n31200) );
  HS65_LH_IVX2 U6796 ( .A(n31200), .Z(n31201) );
  HS65_LH_IVX2 U6797 ( .A(n35239), .Z(n31202) );
  HS65_LH_IVX2 U6799 ( .A(n31202), .Z(n31203) );
  HS65_LH_IVX2 U6800 ( .A(n35241), .Z(n31204) );
  HS65_LH_IVX2 U6802 ( .A(n31204), .Z(n31205) );
  HS65_LH_BFX2 U6803 ( .A(n31185), .Z(n31206) );
  HS65_LH_IVX2 U6805 ( .A(n31209), .Z(n31207) );
  HS65_LH_IVX2 U6806 ( .A(n31207), .Z(n31208) );
  HS65_LH_BFX2 U6808 ( .A(n31210), .Z(n31209) );
  HS65_LH_BFX2 U6810 ( .A(n31211), .Z(n31210) );
  HS65_LH_BFX2 U6815 ( .A(n31212), .Z(n31211) );
  HS65_LH_BFX2 U6816 ( .A(n31213), .Z(n31212) );
  HS65_LH_BFX2 U6817 ( .A(n31214), .Z(n31213) );
  HS65_LH_BFX2 U6818 ( .A(n31215), .Z(n31214) );
  HS65_LH_BFX2 U6819 ( .A(n35574), .Z(n31215) );
  HS65_LH_BFX2 U6820 ( .A(n31218), .Z(n31216) );
  HS65_LH_IVX2 U6821 ( .A(n31221), .Z(n31217) );
  HS65_LH_IVX2 U6822 ( .A(n31217), .Z(n31218) );
  HS65_LH_BFX2 U6823 ( .A(n31220), .Z(n31219) );
  HS65_LH_BFX2 U6824 ( .A(n31222), .Z(n31220) );
  HS65_LH_BFX2 U6825 ( .A(n31223), .Z(n31221) );
  HS65_LH_BFX2 U6826 ( .A(n31224), .Z(n31222) );
  HS65_LH_BFX2 U6827 ( .A(n31225), .Z(n31223) );
  HS65_LH_BFX2 U6828 ( .A(n31226), .Z(n31224) );
  HS65_LH_BFX2 U6829 ( .A(n31227), .Z(n31225) );
  HS65_LH_BFX2 U6830 ( .A(n31228), .Z(n31226) );
  HS65_LH_BFX2 U6831 ( .A(n31229), .Z(n31227) );
  HS65_LH_BFX2 U6832 ( .A(n31230), .Z(n31228) );
  HS65_LH_BFX2 U6833 ( .A(n31231), .Z(n31229) );
  HS65_LH_BFX2 U6834 ( .A(n31232), .Z(n31230) );
  HS65_LH_BFX2 U6835 ( .A(n31233), .Z(n31231) );
  HS65_LH_BFX2 U6836 ( .A(n31234), .Z(n31232) );
  HS65_LH_BFX2 U6837 ( .A(n31235), .Z(n31233) );
  HS65_LH_BFX2 U6838 ( .A(n31236), .Z(n31234) );
  HS65_LH_BFX2 U6839 ( .A(n31237), .Z(n31235) );
  HS65_LH_BFX2 U6840 ( .A(n31238), .Z(n31236) );
  HS65_LH_BFX2 U6842 ( .A(n31239), .Z(n31237) );
  HS65_LH_BFX2 U6843 ( .A(n31240), .Z(n31238) );
  HS65_LH_BFX2 U6844 ( .A(n31241), .Z(n31239) );
  HS65_LH_BFX2 U6845 ( .A(n31242), .Z(n31240) );
  HS65_LH_BFX2 U6846 ( .A(n31243), .Z(n31241) );
  HS65_LH_BFX2 U6847 ( .A(n31244), .Z(n31242) );
  HS65_LH_BFX2 U6848 ( .A(n31245), .Z(n31243) );
  HS65_LH_BFX2 U6849 ( .A(n31246), .Z(n31244) );
  HS65_LH_BFX2 U6850 ( .A(n31247), .Z(n31245) );
  HS65_LH_BFX2 U6851 ( .A(n31248), .Z(n31246) );
  HS65_LH_BFX2 U6852 ( .A(n31249), .Z(n31247) );
  HS65_LH_BFX2 U6853 ( .A(n31250), .Z(n31248) );
  HS65_LH_BFX2 U6854 ( .A(n31251), .Z(n31249) );
  HS65_LH_BFX2 U6855 ( .A(n31252), .Z(n31250) );
  HS65_LH_BFX2 U6856 ( .A(n31253), .Z(n31251) );
  HS65_LH_BFX2 U6857 ( .A(n31254), .Z(n31252) );
  HS65_LH_BFX2 U6858 ( .A(n31255), .Z(n31253) );
  HS65_LH_BFX2 U6859 ( .A(n31256), .Z(n31254) );
  HS65_LH_BFX2 U6860 ( .A(n31257), .Z(n31255) );
  HS65_LH_BFX2 U6861 ( .A(n14485), .Z(n31256) );
  HS65_LH_BFX2 U6862 ( .A(n31258), .Z(n31257) );
  HS65_LH_BFX2 U6863 ( .A(n17956), .Z(n31258) );
  HS65_LH_BFX2 U6864 ( .A(n31260), .Z(n31259) );
  HS65_LH_BFX2 U6865 ( .A(n31261), .Z(n31260) );
  HS65_LH_BFX2 U6866 ( .A(n31262), .Z(n31261) );
  HS65_LH_BFX2 U6867 ( .A(n31263), .Z(n31262) );
  HS65_LH_BFX2 U6868 ( .A(n31264), .Z(n31263) );
  HS65_LH_BFX2 U6869 ( .A(n31265), .Z(n31264) );
  HS65_LH_BFX2 U6870 ( .A(n31266), .Z(n31265) );
  HS65_LH_BFX2 U6871 ( .A(n31267), .Z(n31266) );
  HS65_LH_BFX2 U6872 ( .A(n31268), .Z(n31267) );
  HS65_LH_BFX2 U6873 ( .A(n31269), .Z(n31268) );
  HS65_LH_BFX2 U6874 ( .A(n31270), .Z(n31269) );
  HS65_LH_BFX2 U6875 ( .A(n31271), .Z(n31270) );
  HS65_LH_BFX2 U6876 ( .A(n31272), .Z(n31271) );
  HS65_LH_BFX2 U6877 ( .A(n31273), .Z(n31272) );
  HS65_LH_BFX2 U6878 ( .A(n31274), .Z(n31273) );
  HS65_LH_BFX2 U6879 ( .A(n31275), .Z(n31274) );
  HS65_LH_BFX2 U6880 ( .A(n15566), .Z(n31275) );
  HS65_LH_AOI12X2 U6881 ( .A(n17591), .B(n14524), .C(n14523), .Z(n14541) );
  HS65_LH_BFX2 U6882 ( .A(n14541), .Z(n31276) );
  HS65_LH_BFX2 U6883 ( .A(n31278), .Z(n31277) );
  HS65_LH_BFX2 U6884 ( .A(n31279), .Z(n31278) );
  HS65_LH_BFX2 U6885 ( .A(n31280), .Z(n31279) );
  HS65_LH_BFX2 U6886 ( .A(n31281), .Z(n31280) );
  HS65_LH_BFX2 U6887 ( .A(n31282), .Z(n31281) );
  HS65_LH_BFX2 U6888 ( .A(n31283), .Z(n31282) );
  HS65_LH_BFX2 U6889 ( .A(n31284), .Z(n31283) );
  HS65_LH_BFX2 U6890 ( .A(n31285), .Z(n31284) );
  HS65_LH_BFX2 U6891 ( .A(n31286), .Z(n31285) );
  HS65_LH_BFX2 U6892 ( .A(n31287), .Z(n31286) );
  HS65_LH_BFX2 U6893 ( .A(n31288), .Z(n31287) );
  HS65_LH_BFX2 U6894 ( .A(n31289), .Z(n31288) );
  HS65_LH_BFX2 U6895 ( .A(n31290), .Z(n31289) );
  HS65_LH_BFX2 U6896 ( .A(n31291), .Z(n31290) );
  HS65_LH_BFX2 U6897 ( .A(n31292), .Z(n31291) );
  HS65_LH_BFX2 U6898 ( .A(n31293), .Z(n31292) );
  HS65_LH_BFX2 U6904 ( .A(n31276), .Z(n31293) );
  HS65_LH_OAI12X2 U6905 ( .A(n15395), .B(n32759), .C(n17638), .Z(n14523) );
  HS65_LH_BFX2 U6906 ( .A(n31297), .Z(n31294) );
  HS65_LH_BFX2 U6907 ( .A(n31298), .Z(n31295) );
  HS65_LH_BFX2 U6908 ( .A(n31299), .Z(n31296) );
  HS65_LH_BFX2 U6909 ( .A(n31300), .Z(n31297) );
  HS65_LH_BFX2 U6910 ( .A(n31301), .Z(n31298) );
  HS65_LH_BFX2 U6911 ( .A(n31302), .Z(n31299) );
  HS65_LH_BFX2 U6912 ( .A(n31303), .Z(n31300) );
  HS65_LH_BFX2 U6913 ( .A(n31304), .Z(n31301) );
  HS65_LH_BFX2 U6914 ( .A(n31305), .Z(n31302) );
  HS65_LH_BFX2 U6915 ( .A(n31306), .Z(n31303) );
  HS65_LH_BFX2 U6916 ( .A(n31307), .Z(n31304) );
  HS65_LH_BFX2 U6917 ( .A(n31308), .Z(n31305) );
  HS65_LH_BFX2 U6918 ( .A(n31309), .Z(n31306) );
  HS65_LH_BFX2 U6919 ( .A(n31310), .Z(n31307) );
  HS65_LH_BFX2 U6920 ( .A(n31311), .Z(n31308) );
  HS65_LH_BFX2 U6921 ( .A(n31312), .Z(n31309) );
  HS65_LH_BFX2 U6922 ( .A(n31313), .Z(n31310) );
  HS65_LH_BFX2 U6923 ( .A(n31314), .Z(n31311) );
  HS65_LH_BFX2 U6924 ( .A(n31315), .Z(n31312) );
  HS65_LH_BFX2 U6925 ( .A(n31316), .Z(n31313) );
  HS65_LH_BFX2 U6926 ( .A(n31317), .Z(n31314) );
  HS65_LH_BFX2 U6927 ( .A(n31318), .Z(n31315) );
  HS65_LH_BFX2 U6928 ( .A(n31319), .Z(n31316) );
  HS65_LH_BFX2 U6929 ( .A(n31320), .Z(n31317) );
  HS65_LH_BFX2 U6930 ( .A(n31321), .Z(n31318) );
  HS65_LH_BFX2 U6932 ( .A(n31322), .Z(n31319) );
  HS65_LH_BFX2 U6934 ( .A(n31323), .Z(n31320) );
  HS65_LH_BFX2 U6936 ( .A(n31324), .Z(n31321) );
  HS65_LH_BFX2 U6938 ( .A(n31325), .Z(n31322) );
  HS65_LH_BFX2 U6940 ( .A(n31326), .Z(n31323) );
  HS65_LH_BFX2 U6941 ( .A(n31327), .Z(n31324) );
  HS65_LH_BFX2 U6942 ( .A(n31328), .Z(n31325) );
  HS65_LH_BFX2 U6943 ( .A(n31329), .Z(n31326) );
  HS65_LH_BFX2 U6944 ( .A(n31330), .Z(n31327) );
  HS65_LH_BFX2 U6987 ( .A(n31331), .Z(n31328) );
  HS65_LH_BFX2 U6988 ( .A(n31332), .Z(n31329) );
  HS65_LH_BFX2 U6990 ( .A(n31333), .Z(n31330) );
  HS65_LH_BFX2 U6991 ( .A(n31334), .Z(n31331) );
  HS65_LH_BFX2 U6992 ( .A(n31335), .Z(n31332) );
  HS65_LH_BFX2 U6993 ( .A(n31336), .Z(n31333) );
  HS65_LH_BFX2 U6994 ( .A(n31337), .Z(n31334) );
  HS65_LH_BFX2 U6995 ( .A(n31338), .Z(n31335) );
  HS65_LH_BFX2 U6996 ( .A(n15563), .Z(n31336) );
  HS65_LH_BFX2 U6997 ( .A(n31339), .Z(n31337) );
  HS65_LH_BFX2 U6998 ( .A(n31340), .Z(n31338) );
  HS65_LH_BFX2 U6999 ( .A(n31341), .Z(n31339) );
  HS65_LH_BFX2 U7000 ( .A(n31342), .Z(n31340) );
  HS65_LH_BFX2 U7001 ( .A(n31343), .Z(n31341) );
  HS65_LH_BFX2 U7002 ( .A(n31344), .Z(n31342) );
  HS65_LH_BFX2 U7003 ( .A(n31345), .Z(n31343) );
  HS65_LH_BFX2 U7004 ( .A(n31346), .Z(n31344) );
  HS65_LH_BFX2 U7005 ( .A(n14907), .Z(n31345) );
  HS65_LH_BFX2 U7006 ( .A(n31347), .Z(n31346) );
  HS65_LH_BFX2 U7007 ( .A(n31348), .Z(n31347) );
  HS65_LH_BFX2 U7008 ( .A(n17905), .Z(n31348) );
  HS65_LH_IVX2 U7009 ( .A(n31351), .Z(n31349) );
  HS65_LH_IVX2 U7010 ( .A(n31349), .Z(n31350) );
  HS65_LH_BFX2 U7011 ( .A(n31352), .Z(n31351) );
  HS65_LH_BFX2 U7012 ( .A(n31353), .Z(n31352) );
  HS65_LH_BFX2 U7013 ( .A(n31354), .Z(n31353) );
  HS65_LH_BFX2 U7014 ( .A(n31355), .Z(n31354) );
  HS65_LH_BFX2 U7015 ( .A(n31356), .Z(n31355) );
  HS65_LH_BFX2 U7016 ( .A(n31357), .Z(n31356) );
  HS65_LH_BFX2 U7018 ( .A(n31358), .Z(n31357) );
  HS65_LH_BFX2 U7026 ( .A(n31359), .Z(n31358) );
  HS65_LH_BFX2 U7075 ( .A(n31360), .Z(n31359) );
  HS65_LH_BFX2 U7076 ( .A(n31361), .Z(n31360) );
  HS65_LH_BFX2 U7077 ( .A(n31362), .Z(n31361) );
  HS65_LH_BFX2 U7078 ( .A(n31363), .Z(n31362) );
  HS65_LH_BFX2 U7079 ( .A(n31364), .Z(n31363) );
  HS65_LH_BFX2 U7080 ( .A(n31365), .Z(n31364) );
  HS65_LH_BFX2 U7081 ( .A(n15718), .Z(n31365) );
  HS65_LH_BFX2 U7083 ( .A(n31367), .Z(n31366) );
  HS65_LH_BFX2 U7084 ( .A(n31368), .Z(n31367) );
  HS65_LH_BFX2 U7085 ( .A(n31369), .Z(n31368) );
  HS65_LH_BFX2 U7086 ( .A(n31370), .Z(n31369) );
  HS65_LH_BFX2 U7087 ( .A(n31371), .Z(n31370) );
  HS65_LH_BFX2 U7088 ( .A(n31372), .Z(n31371) );
  HS65_LH_BFX2 U7089 ( .A(n31373), .Z(n31372) );
  HS65_LH_BFX2 U7090 ( .A(n31374), .Z(n31373) );
  HS65_LH_BFX2 U7092 ( .A(n31375), .Z(n31374) );
  HS65_LH_BFX2 U7093 ( .A(n31376), .Z(n31375) );
  HS65_LH_BFX2 U7094 ( .A(n31377), .Z(n31376) );
  HS65_LH_BFX2 U7095 ( .A(n31378), .Z(n31377) );
  HS65_LH_BFX2 U7096 ( .A(n31379), .Z(n31378) );
  HS65_LH_BFX2 U7097 ( .A(n31380), .Z(n31379) );
  HS65_LH_BFX2 U7098 ( .A(n31381), .Z(n31380) );
  HS65_LH_BFX2 U7099 ( .A(n31382), .Z(n31381) );
  HS65_LH_BFX2 U7100 ( .A(n31383), .Z(n31382) );
  HS65_LH_BFX2 U7101 ( .A(n15568), .Z(n31383) );
  HS65_LH_BFX2 U7102 ( .A(n31385), .Z(n31384) );
  HS65_LH_BFX2 U7103 ( .A(n31386), .Z(n31385) );
  HS65_LH_BFX2 U7104 ( .A(n31387), .Z(n31386) );
  HS65_LH_BFX2 U7106 ( .A(n31388), .Z(n31387) );
  HS65_LH_BFX2 U7108 ( .A(n31389), .Z(n31388) );
  HS65_LH_BFX2 U7110 ( .A(n31390), .Z(n31389) );
  HS65_LH_BFX2 U7159 ( .A(n31391), .Z(n31390) );
  HS65_LH_BFX2 U7160 ( .A(n31392), .Z(n31391) );
  HS65_LH_BFX2 U7161 ( .A(n31393), .Z(n31392) );
  HS65_LH_BFX2 U7162 ( .A(n31394), .Z(n31393) );
  HS65_LH_BFX2 U7163 ( .A(n31395), .Z(n31394) );
  HS65_LH_BFX2 U7164 ( .A(n31396), .Z(n31395) );
  HS65_LH_BFX2 U7165 ( .A(n31397), .Z(n31396) );
  HS65_LH_BFX2 U7166 ( .A(n31398), .Z(n31397) );
  HS65_LH_BFX2 U7167 ( .A(n31399), .Z(n31398) );
  HS65_LH_BFX2 U7168 ( .A(n31400), .Z(n31399) );
  HS65_LH_BFX2 U7170 ( .A(n31401), .Z(n31400) );
  HS65_LH_BFX2 U7172 ( .A(n14539), .Z(n31401) );
  HS65_LH_BFX2 U7174 ( .A(n31403), .Z(n31402) );
  HS65_LH_BFX2 U7176 ( .A(n31404), .Z(n31403) );
  HS65_LH_BFX2 U7178 ( .A(n31405), .Z(n31404) );
  HS65_LH_BFX2 U7180 ( .A(n31406), .Z(n31405) );
  HS65_LH_BFX2 U7181 ( .A(n31407), .Z(n31406) );
  HS65_LH_BFX2 U7183 ( .A(n31408), .Z(n31407) );
  HS65_LH_BFX2 U7185 ( .A(n31409), .Z(n31408) );
  HS65_LH_BFX2 U7187 ( .A(n31410), .Z(n31409) );
  HS65_LH_BFX2 U7189 ( .A(n31411), .Z(n31410) );
  HS65_LH_BFX2 U7191 ( .A(n31412), .Z(n31411) );
  HS65_LH_BFX2 U7192 ( .A(n31413), .Z(n31412) );
  HS65_LH_BFX2 U7194 ( .A(n31414), .Z(n31413) );
  HS65_LH_BFX2 U7219 ( .A(n31415), .Z(n31414) );
  HS65_LH_BFX2 U7220 ( .A(n31416), .Z(n31415) );
  HS65_LH_BFX2 U7221 ( .A(n31417), .Z(n31416) );
  HS65_LH_BFX2 U7222 ( .A(n31418), .Z(n31417) );
  HS65_LH_BFX2 U7223 ( .A(n15576), .Z(n31418) );
  HS65_LH_BFX2 U7224 ( .A(n31420), .Z(n31419) );
  HS65_LH_BFX2 U7225 ( .A(n31421), .Z(n31420) );
  HS65_LH_BFX2 U7226 ( .A(n31422), .Z(n31421) );
  HS65_LH_BFX2 U7227 ( .A(n31423), .Z(n31422) );
  HS65_LH_BFX2 U7228 ( .A(n31424), .Z(n31423) );
  HS65_LH_BFX2 U7229 ( .A(n31425), .Z(n31424) );
  HS65_LH_BFX2 U7244 ( .A(n31426), .Z(n31425) );
  HS65_LH_BFX2 U7245 ( .A(n31427), .Z(n31426) );
  HS65_LH_BFX2 U7247 ( .A(n31428), .Z(n31427) );
  HS65_LH_BFX2 U7248 ( .A(n31429), .Z(n31428) );
  HS65_LH_BFX2 U7250 ( .A(n31430), .Z(n31429) );
  HS65_LH_BFX2 U7251 ( .A(n31431), .Z(n31430) );
  HS65_LH_BFX2 U7253 ( .A(n31432), .Z(n31431) );
  HS65_LH_BFX2 U7254 ( .A(n31433), .Z(n31432) );
  HS65_LH_BFX2 U7256 ( .A(n31434), .Z(n31433) );
  HS65_LH_BFX2 U7257 ( .A(n31435), .Z(n31434) );
  HS65_LH_BFX2 U7259 ( .A(n31436), .Z(n31435) );
  HS65_LH_BFX2 U7260 ( .A(n31437), .Z(n31436) );
  HS65_LH_BFX2 U7262 ( .A(n14266), .Z(n31437) );
  HS65_LH_BFX2 U7263 ( .A(n31439), .Z(n31438) );
  HS65_LH_BFX2 U7265 ( .A(n31440), .Z(n31439) );
  HS65_LH_BFX2 U7266 ( .A(n31441), .Z(n31440) );
  HS65_LH_BFX2 U7268 ( .A(n31442), .Z(n31441) );
  HS65_LH_BFX2 U7269 ( .A(n31443), .Z(n31442) );
  HS65_LH_BFX2 U7271 ( .A(n31444), .Z(n31443) );
  HS65_LH_BFX2 U7272 ( .A(n31445), .Z(n31444) );
  HS65_LH_BFX2 U7274 ( .A(n31446), .Z(n31445) );
  HS65_LH_BFX2 U7275 ( .A(n31447), .Z(n31446) );
  HS65_LH_BFX2 U7277 ( .A(n31448), .Z(n31447) );
  HS65_LH_BFX2 U7278 ( .A(n31449), .Z(n31448) );
  HS65_LH_BFX2 U7280 ( .A(n31450), .Z(n31449) );
  HS65_LH_BFX2 U7281 ( .A(n31451), .Z(n31450) );
  HS65_LH_BFX2 U7283 ( .A(n31452), .Z(n31451) );
  HS65_LH_BFX2 U7284 ( .A(n31453), .Z(n31452) );
  HS65_LH_BFX2 U7286 ( .A(n31454), .Z(n31453) );
  HS65_LH_BFX2 U7287 ( .A(n31455), .Z(n31454) );
  HS65_LH_BFX2 U7289 ( .A(n31456), .Z(n31455) );
  HS65_LH_BFX2 U7290 ( .A(n14268), .Z(n31456) );
  HS65_LH_BFX2 U7292 ( .A(n31458), .Z(n31457) );
  HS65_LH_BFX2 U7293 ( .A(n31459), .Z(n31458) );
  HS65_LH_BFX2 U7294 ( .A(n31460), .Z(n31459) );
  HS65_LH_BFX2 U7295 ( .A(n31461), .Z(n31460) );
  HS65_LH_BFX2 U7297 ( .A(n31462), .Z(n31461) );
  HS65_LH_BFX2 U7299 ( .A(n31463), .Z(n31462) );
  HS65_LH_BFX2 U7301 ( .A(n31464), .Z(n31463) );
  HS65_LH_BFX2 U7303 ( .A(n31465), .Z(n31464) );
  HS65_LH_BFX2 U7308 ( .A(n31466), .Z(n31465) );
  HS65_LH_BFX2 U7309 ( .A(n31467), .Z(n31466) );
  HS65_LH_BFX2 U7310 ( .A(n31468), .Z(n31467) );
  HS65_LH_BFX2 U7311 ( .A(n31469), .Z(n31468) );
  HS65_LH_BFX2 U7312 ( .A(n31470), .Z(n31469) );
  HS65_LH_BFX2 U7313 ( .A(n31471), .Z(n31470) );
  HS65_LH_BFX2 U7314 ( .A(n31472), .Z(n31471) );
  HS65_LH_BFX2 U7315 ( .A(n31473), .Z(n31472) );
  HS65_LH_BFX2 U7316 ( .A(n31474), .Z(n31473) );
  HS65_LH_BFX2 U7317 ( .A(n31475), .Z(n31474) );
  HS65_LH_BFX2 U7318 ( .A(n31476), .Z(n31475) );
  HS65_LH_BFX2 U7319 ( .A(n17247), .Z(n31476) );
  HS65_LH_BFX2 U7320 ( .A(n31478), .Z(n31477) );
  HS65_LH_BFX2 U7321 ( .A(n31479), .Z(n31478) );
  HS65_LH_BFX2 U7322 ( .A(n31480), .Z(n31479) );
  HS65_LH_BFX2 U7323 ( .A(n31481), .Z(n31480) );
  HS65_LH_BFX2 U7324 ( .A(n31482), .Z(n31481) );
  HS65_LH_BFX2 U7325 ( .A(n31483), .Z(n31482) );
  HS65_LH_BFX2 U7326 ( .A(n31484), .Z(n31483) );
  HS65_LH_BFX2 U7327 ( .A(n31485), .Z(n31484) );
  HS65_LH_BFX2 U7328 ( .A(n31486), .Z(n31485) );
  HS65_LH_BFX2 U7329 ( .A(n31487), .Z(n31486) );
  HS65_LH_BFX2 U7330 ( .A(n31488), .Z(n31487) );
  HS65_LH_BFX2 U7331 ( .A(n31489), .Z(n31488) );
  HS65_LH_BFX2 U7332 ( .A(n31490), .Z(n31489) );
  HS65_LH_BFX2 U7333 ( .A(n31491), .Z(n31490) );
  HS65_LH_BFX2 U7334 ( .A(n31492), .Z(n31491) );
  HS65_LH_BFX2 U7335 ( .A(n31493), .Z(n31492) );
  HS65_LH_BFX2 U7336 ( .A(n31494), .Z(n31493) );
  HS65_LH_BFX2 U7337 ( .A(n31495), .Z(n31494) );
  HS65_LH_BFX2 U7338 ( .A(n14263), .Z(n31495) );
  HS65_LH_BFX2 U7339 ( .A(n31497), .Z(n31496) );
  HS65_LH_BFX2 U7340 ( .A(n31498), .Z(n31497) );
  HS65_LH_BFX2 U7341 ( .A(n31499), .Z(n31498) );
  HS65_LH_BFX2 U7342 ( .A(n31500), .Z(n31499) );
  HS65_LH_BFX2 U7344 ( .A(n31501), .Z(n31500) );
  HS65_LH_BFX2 U7346 ( .A(n31502), .Z(n31501) );
  HS65_LH_BFX2 U7348 ( .A(n31503), .Z(n31502) );
  HS65_LH_BFX2 U7350 ( .A(n31504), .Z(n31503) );
  HS65_LH_BFX2 U7352 ( .A(n31505), .Z(n31504) );
  HS65_LH_BFX2 U7354 ( .A(n31506), .Z(n31505) );
  HS65_LH_BFX2 U7356 ( .A(n31507), .Z(n31506) );
  HS65_LH_BFX2 U7358 ( .A(n31508), .Z(n31507) );
  HS65_LH_BFX2 U7360 ( .A(n31509), .Z(n31508) );
  HS65_LH_BFX2 U7362 ( .A(n31510), .Z(n31509) );
  HS65_LH_BFX2 U7364 ( .A(n31511), .Z(n31510) );
  HS65_LH_BFX2 U7366 ( .A(n31512), .Z(n31511) );
  HS65_LH_BFX2 U7417 ( .A(n31513), .Z(n31512) );
  HS65_LH_BFX2 U7419 ( .A(n31514), .Z(n31513) );
  HS65_LH_BFX2 U7421 ( .A(n14264), .Z(n31514) );
  HS65_LH_BFX2 U7423 ( .A(n31516), .Z(n31515) );
  HS65_LH_BFX2 U7425 ( .A(n31517), .Z(n31516) );
  HS65_LH_BFX2 U7427 ( .A(n31518), .Z(n31517) );
  HS65_LH_BFX2 U7429 ( .A(n31519), .Z(n31518) );
  HS65_LH_BFX2 U7431 ( .A(n31520), .Z(n31519) );
  HS65_LH_BFX2 U7433 ( .A(n31521), .Z(n31520) );
  HS65_LH_BFX2 U7435 ( .A(n31522), .Z(n31521) );
  HS65_LH_BFX2 U7436 ( .A(n31523), .Z(n31522) );
  HS65_LH_BFX2 U7438 ( .A(n31524), .Z(n31523) );
  HS65_LH_BFX2 U7440 ( .A(n31525), .Z(n31524) );
  HS65_LH_BFX2 U7442 ( .A(n31526), .Z(n31525) );
  HS65_LH_BFX2 U7444 ( .A(n31527), .Z(n31526) );
  HS65_LH_BFX2 U7446 ( .A(n31528), .Z(n31527) );
  HS65_LH_BFX2 U7448 ( .A(n31529), .Z(n31528) );
  HS65_LH_BFX2 U7504 ( .A(n31530), .Z(n31529) );
  HS65_LH_BFX2 U7505 ( .A(n31531), .Z(n31530) );
  HS65_LH_BFX2 U7506 ( .A(n31532), .Z(n31531) );
  HS65_LH_BFX2 U7507 ( .A(n31533), .Z(n31532) );
  HS65_LH_BFX2 U7509 ( .A(n14267), .Z(n31533) );
  HS65_LH_BFX2 U7511 ( .A(n31535), .Z(n31534) );
  HS65_LH_BFX2 U7513 ( .A(n31536), .Z(n31535) );
  HS65_LH_BFX2 U7515 ( .A(n31537), .Z(n31536) );
  HS65_LH_BFX2 U7517 ( .A(n31538), .Z(n31537) );
  HS65_LH_BFX2 U7519 ( .A(n31539), .Z(n31538) );
  HS65_LH_BFX2 U7521 ( .A(n31540), .Z(n31539) );
  HS65_LH_BFX2 U7523 ( .A(n31541), .Z(n31540) );
  HS65_LH_BFX2 U7525 ( .A(n31542), .Z(n31541) );
  HS65_LH_BFX2 U7527 ( .A(n31543), .Z(n31542) );
  HS65_LH_BFX2 U7529 ( .A(n31544), .Z(n31543) );
  HS65_LH_BFX2 U7531 ( .A(n31545), .Z(n31544) );
  HS65_LH_BFX2 U7533 ( .A(n31546), .Z(n31545) );
  HS65_LH_BFX2 U7535 ( .A(n31547), .Z(n31546) );
  HS65_LH_BFX2 U7537 ( .A(n31548), .Z(n31547) );
  HS65_LH_BFX2 U7562 ( .A(n31549), .Z(n31548) );
  HS65_LH_BFX2 U7563 ( .A(n31550), .Z(n31549) );
  HS65_LH_BFX2 U7564 ( .A(n31551), .Z(n31550) );
  HS65_LH_BFX2 U7565 ( .A(n31552), .Z(n31551) );
  HS65_LH_BFX2 U7566 ( .A(n14301), .Z(n31552) );
  HS65_LH_BFX2 U7567 ( .A(n31554), .Z(n31553) );
  HS65_LH_BFX2 U7568 ( .A(n31555), .Z(n31554) );
  HS65_LH_BFX2 U7569 ( .A(n31556), .Z(n31555) );
  HS65_LH_BFX2 U7570 ( .A(n31557), .Z(n31556) );
  HS65_LH_BFX2 U7571 ( .A(n31558), .Z(n31557) );
  HS65_LH_BFX2 U7572 ( .A(n31559), .Z(n31558) );
  HS65_LH_BFX2 U7573 ( .A(n31560), .Z(n31559) );
  HS65_LH_BFX2 U7574 ( .A(n31561), .Z(n31560) );
  HS65_LH_BFX2 U7575 ( .A(n31562), .Z(n31561) );
  HS65_LH_BFX2 U7576 ( .A(n31563), .Z(n31562) );
  HS65_LH_BFX2 U7577 ( .A(n31564), .Z(n31563) );
  HS65_LH_BFX2 U7578 ( .A(n31565), .Z(n31564) );
  HS65_LH_BFX2 U7579 ( .A(n31566), .Z(n31565) );
  HS65_LH_BFX2 U7580 ( .A(n31567), .Z(n31566) );
  HS65_LH_BFX2 U7581 ( .A(n31568), .Z(n31567) );
  HS65_LH_BFX2 U7582 ( .A(n31569), .Z(n31568) );
  HS65_LH_BFX2 U7583 ( .A(n31570), .Z(n31569) );
  HS65_LH_BFX2 U7584 ( .A(n31571), .Z(n31570) );
  HS65_LH_BFX2 U7585 ( .A(n14265), .Z(n31571) );
  HS65_LH_BFX2 U7586 ( .A(n31574), .Z(n31572) );
  HS65_LH_IVX2 U7590 ( .A(n31576), .Z(n31573) );
  HS65_LH_IVX2 U7592 ( .A(n31573), .Z(n31574) );
  HS65_LH_BFX2 U7593 ( .A(n31580), .Z(n31575) );
  HS65_LH_BFX2 U7595 ( .A(n31577), .Z(n31576) );
  HS65_LH_BFX2 U7596 ( .A(n31578), .Z(n31577) );
  HS65_LH_BFX2 U7598 ( .A(n31579), .Z(n31578) );
  HS65_LH_BFX2 U7599 ( .A(n31575), .Z(n31579) );
  HS65_LH_BFX2 U7601 ( .A(n31581), .Z(n31580) );
  HS65_LH_BFX2 U7602 ( .A(n31582), .Z(n31581) );
  HS65_LH_BFX2 U7604 ( .A(n31583), .Z(n31582) );
  HS65_LH_BFX2 U7605 ( .A(n31584), .Z(n31583) );
  HS65_LH_BFX2 U7607 ( .A(n31585), .Z(n31584) );
  HS65_LH_BFX2 U7608 ( .A(n31586), .Z(n31585) );
  HS65_LH_BFX2 U7610 ( .A(n31587), .Z(n31586) );
  HS65_LH_BFX2 U7611 ( .A(n31588), .Z(n31587) );
  HS65_LH_BFX2 U7613 ( .A(n31589), .Z(n31588) );
  HS65_LH_BFX2 U7614 ( .A(n31590), .Z(n31589) );
  HS65_LH_BFX2 U7616 ( .A(n31591), .Z(n31590) );
  HS65_LH_BFX2 U7617 ( .A(n31592), .Z(n31591) );
  HS65_LH_BFX2 U7619 ( .A(n14255), .Z(n31592) );
  HS65_LH_BFX2 U7620 ( .A(n31595), .Z(n31593) );
  HS65_LH_BFX2 U7622 ( .A(n31602), .Z(n31594) );
  HS65_LH_BFX2 U7623 ( .A(n31596), .Z(n31595) );
  HS65_LH_BFX2 U7625 ( .A(n31597), .Z(n31596) );
  HS65_LH_BFX2 U7626 ( .A(n31598), .Z(n31597) );
  HS65_LH_BFX2 U7628 ( .A(n31599), .Z(n31598) );
  HS65_LH_BFX2 U7629 ( .A(n31600), .Z(n31599) );
  HS65_LH_BFX2 U7631 ( .A(n31601), .Z(n31600) );
  HS65_LH_BFX2 U7632 ( .A(n31594), .Z(n31601) );
  HS65_LH_BFX2 U7634 ( .A(n31603), .Z(n31602) );
  HS65_LH_BFX2 U7635 ( .A(n31604), .Z(n31603) );
  HS65_LH_BFX2 U7637 ( .A(n31605), .Z(n31604) );
  HS65_LH_BFX2 U7638 ( .A(n31606), .Z(n31605) );
  HS65_LH_BFX2 U7640 ( .A(n31607), .Z(n31606) );
  HS65_LH_BFX2 U7641 ( .A(n31608), .Z(n31607) );
  HS65_LH_BFX2 U7643 ( .A(n31609), .Z(n31608) );
  HS65_LH_BFX2 U7644 ( .A(n31610), .Z(n31609) );
  HS65_LH_BFX2 U7646 ( .A(n31611), .Z(n31610) );
  HS65_LH_BFX2 U7648 ( .A(n31612), .Z(n31611) );
  HS65_LH_BFX2 U7673 ( .A(n14258), .Z(n31612) );
  HS65_LH_BFX2 U7674 ( .A(n31615), .Z(n31613) );
  HS65_LH_IVX2 U7675 ( .A(n31617), .Z(n31614) );
  HS65_LH_IVX2 U7676 ( .A(n31614), .Z(n31615) );
  HS65_LH_BFX2 U7677 ( .A(n31627), .Z(n31616) );
  HS65_LH_BFX2 U7678 ( .A(n31618), .Z(n31617) );
  HS65_LH_BFX2 U7679 ( .A(n31619), .Z(n31618) );
  HS65_LH_BFX2 U7680 ( .A(n31620), .Z(n31619) );
  HS65_LH_BFX2 U7681 ( .A(n31621), .Z(n31620) );
  HS65_LH_BFX2 U7682 ( .A(n31622), .Z(n31621) );
  HS65_LH_BFX2 U7683 ( .A(n31623), .Z(n31622) );
  HS65_LH_BFX2 U7684 ( .A(n31624), .Z(n31623) );
  HS65_LH_BFX2 U7685 ( .A(n31625), .Z(n31624) );
  HS65_LH_BFX2 U7686 ( .A(n31626), .Z(n31625) );
  HS65_LH_BFX2 U7687 ( .A(n31616), .Z(n31626) );
  HS65_LH_BFX2 U7688 ( .A(n31628), .Z(n31627) );
  HS65_LH_BFX2 U7689 ( .A(n31629), .Z(n31628) );
  HS65_LH_BFX2 U7690 ( .A(n31630), .Z(n31629) );
  HS65_LH_BFX2 U7692 ( .A(n31631), .Z(n31630) );
  HS65_LH_BFX2 U7693 ( .A(n31632), .Z(n31631) );
  HS65_LH_BFX2 U7694 ( .A(n31633), .Z(n31632) );
  HS65_LH_BFX2 U7695 ( .A(n14259), .Z(n31633) );
  HS65_LH_BFX2 U7696 ( .A(n31636), .Z(n31634) );
  HS65_LH_BFX2 U7697 ( .A(n31648), .Z(n31635) );
  HS65_LH_BFX2 U7699 ( .A(n31637), .Z(n31636) );
  HS65_LH_BFX2 U7700 ( .A(n31638), .Z(n31637) );
  HS65_LH_BFX2 U7702 ( .A(n31639), .Z(n31638) );
  HS65_LH_BFX2 U7703 ( .A(n31640), .Z(n31639) );
  HS65_LH_BFX2 U7705 ( .A(n31641), .Z(n31640) );
  HS65_LH_BFX2 U7706 ( .A(n31642), .Z(n31641) );
  HS65_LH_BFX2 U7708 ( .A(n31643), .Z(n31642) );
  HS65_LH_BFX2 U7709 ( .A(n31644), .Z(n31643) );
  HS65_LH_BFX2 U7711 ( .A(n31645), .Z(n31644) );
  HS65_LH_BFX2 U7712 ( .A(n31646), .Z(n31645) );
  HS65_LH_BFX2 U7714 ( .A(n31647), .Z(n31646) );
  HS65_LH_BFX2 U7715 ( .A(n31635), .Z(n31647) );
  HS65_LH_BFX2 U7717 ( .A(n31649), .Z(n31648) );
  HS65_LH_BFX2 U7718 ( .A(n31650), .Z(n31649) );
  HS65_LH_BFX2 U7720 ( .A(n31651), .Z(n31650) );
  HS65_LH_BFX2 U7721 ( .A(n31652), .Z(n31651) );
  HS65_LH_BFX2 U7723 ( .A(n31653), .Z(n31652) );
  HS65_LH_BFX2 U7724 ( .A(n14260), .Z(n31653) );
  HS65_LH_BFX2 U7726 ( .A(n31656), .Z(n31654) );
  HS65_LH_IVX2 U7727 ( .A(n31658), .Z(n31655) );
  HS65_LH_IVX2 U7729 ( .A(n31655), .Z(n31656) );
  HS65_LH_BFX2 U7730 ( .A(n31671), .Z(n31657) );
  HS65_LH_BFX2 U7732 ( .A(n31659), .Z(n31658) );
  HS65_LH_BFX2 U7733 ( .A(n31660), .Z(n31659) );
  HS65_LH_BFX2 U7735 ( .A(n31661), .Z(n31660) );
  HS65_LH_BFX2 U7736 ( .A(n31662), .Z(n31661) );
  HS65_LH_BFX2 U7738 ( .A(n31663), .Z(n31662) );
  HS65_LH_BFX2 U7739 ( .A(n31664), .Z(n31663) );
  HS65_LH_BFX2 U7741 ( .A(n31665), .Z(n31664) );
  HS65_LH_BFX2 U7742 ( .A(n31666), .Z(n31665) );
  HS65_LH_BFX2 U7744 ( .A(n31667), .Z(n31666) );
  HS65_LH_BFX2 U7745 ( .A(n31668), .Z(n31667) );
  HS65_LH_BFX2 U7747 ( .A(n31669), .Z(n31668) );
  HS65_LH_BFX2 U7748 ( .A(n31670), .Z(n31669) );
  HS65_LH_BFX2 U7750 ( .A(n31657), .Z(n31670) );
  HS65_LH_BFX2 U7751 ( .A(n31672), .Z(n31671) );
  HS65_LH_BFX2 U7753 ( .A(n31673), .Z(n31672) );
  HS65_LH_BFX2 U7755 ( .A(n31674), .Z(n31673) );
  HS65_LH_BFX2 U7757 ( .A(n14276), .Z(n31674) );
  HS65_LH_BFX2 U7782 ( .A(n31676), .Z(n31675) );
  HS65_LH_BFX2 U7783 ( .A(n31677), .Z(n31676) );
  HS65_LH_BFX2 U7784 ( .A(n31678), .Z(n31677) );
  HS65_LH_BFX2 U7785 ( .A(n31679), .Z(n31678) );
  HS65_LH_BFX2 U7786 ( .A(n31680), .Z(n31679) );
  HS65_LH_BFX2 U7787 ( .A(n31681), .Z(n31680) );
  HS65_LH_BFX2 U7788 ( .A(n31682), .Z(n31681) );
  HS65_LH_BFX2 U7789 ( .A(n31683), .Z(n31682) );
  HS65_LH_BFX2 U7790 ( .A(n31684), .Z(n31683) );
  HS65_LH_BFX2 U7791 ( .A(n31685), .Z(n31684) );
  HS65_LH_BFX2 U7792 ( .A(n31686), .Z(n31685) );
  HS65_LH_BFX2 U7793 ( .A(n31687), .Z(n31686) );
  HS65_LH_BFX2 U7794 ( .A(n31688), .Z(n31687) );
  HS65_LH_BFX2 U7795 ( .A(n31689), .Z(n31688) );
  HS65_LH_BFX2 U7796 ( .A(n31691), .Z(n31689) );
  HS65_LH_BFX2 U7797 ( .A(n14261), .Z(n31690) );
  HS65_LH_BFX2 U7798 ( .A(n31693), .Z(n31691) );
  HS65_LH_BFX2 U7799 ( .A(n31690), .Z(n31692) );
  HS65_LH_BFX2 U7800 ( .A(n31694), .Z(n31693) );
  HS65_LH_BFX2 U7801 ( .A(n31692), .Z(n31694) );
  HS65_LH_BFX2 U7802 ( .A(n31697), .Z(n31695) );
  HS65_LH_IVX2 U7803 ( .A(n31699), .Z(n31696) );
  HS65_LH_IVX2 U7804 ( .A(n31696), .Z(n31697) );
  HS65_LH_BFX2 U7805 ( .A(n31715), .Z(n31698) );
  HS65_LH_BFX2 U7806 ( .A(n31700), .Z(n31699) );
  HS65_LH_BFX2 U7807 ( .A(n31701), .Z(n31700) );
  HS65_LH_BFX2 U7809 ( .A(n31702), .Z(n31701) );
  HS65_LH_BFX2 U7810 ( .A(n31703), .Z(n31702) );
  HS65_LH_BFX2 U7812 ( .A(n31704), .Z(n31703) );
  HS65_LH_BFX2 U7813 ( .A(n31705), .Z(n31704) );
  HS65_LH_BFX2 U7815 ( .A(n31706), .Z(n31705) );
  HS65_LH_BFX2 U7816 ( .A(n31707), .Z(n31706) );
  HS65_LH_BFX2 U7818 ( .A(n31708), .Z(n31707) );
  HS65_LH_BFX2 U7819 ( .A(n31710), .Z(n31708) );
  HS65_LH_BFX2 U7821 ( .A(n14262), .Z(n31709) );
  HS65_LH_BFX2 U7822 ( .A(n31712), .Z(n31710) );
  HS65_LH_BFX2 U7824 ( .A(n31709), .Z(n31711) );
  HS65_LH_BFX2 U7825 ( .A(n31714), .Z(n31712) );
  HS65_LH_BFX2 U7827 ( .A(n31711), .Z(n31713) );
  HS65_LH_BFX2 U7828 ( .A(n31698), .Z(n31714) );
  HS65_LH_BFX2 U7830 ( .A(n31713), .Z(n31715) );
  HS65_LH_BFX2 U7831 ( .A(n31741), .Z(n31716) );
  HS65_LH_BFX2 U7833 ( .A(n31720), .Z(n31717) );
  HS65_LH_BFX2 U7834 ( .A(n2358), .Z(n31718) );
  HS65_LH_IVX2 U7836 ( .A(n31769), .Z(n31719) );
  HS65_LH_IVX2 U7837 ( .A(n31719), .Z(n31720) );
  HS65_LH_IVX2 U7839 ( .A(n31725), .Z(n31721) );
  HS65_LH_IVX2 U7840 ( .A(n31721), .Z(n31722) );
  HS65_LH_BFX2 U7842 ( .A(n2357), .Z(n31723) );
  HS65_LH_BFX2 U7843 ( .A(n31723), .Z(n31724) );
  HS65_LH_BFX2 U7845 ( .A(n31727), .Z(n31725) );
  HS65_LH_BFX2 U7846 ( .A(n31724), .Z(n31726) );
  HS65_LH_BFX2 U7848 ( .A(n31729), .Z(n31727) );
  HS65_LH_BFX2 U7849 ( .A(n31726), .Z(n31728) );
  HS65_LH_BFX2 U7851 ( .A(n31731), .Z(n31729) );
  HS65_LH_BFX2 U7852 ( .A(n31728), .Z(n31730) );
  HS65_LH_BFX2 U7854 ( .A(n31733), .Z(n31731) );
  HS65_LH_BFX2 U7855 ( .A(n31730), .Z(n31732) );
  HS65_LH_BFX2 U7857 ( .A(n31735), .Z(n31733) );
  HS65_LH_BFX2 U7858 ( .A(n31732), .Z(n31734) );
  HS65_LH_BFX2 U7860 ( .A(n31738), .Z(n31735) );
  HS65_LH_BFX2 U7862 ( .A(n31734), .Z(n31736) );
  HS65_LH_IVX2 U7864 ( .A(n31743), .Z(n31737) );
  HS65_LH_IVX2 U7866 ( .A(n31737), .Z(n31738) );
  HS65_LH_BFX2 U7916 ( .A(n31736), .Z(n31739) );
  HS65_LH_IVX2 U7917 ( .A(n31739), .Z(n31740) );
  HS65_LH_IVX2 U7918 ( .A(n31740), .Z(n31741) );
  HS65_LH_IVX2 U7919 ( .A(n31718), .Z(n31742) );
  HS65_LH_IVX2 U7920 ( .A(n31742), .Z(n31743) );
  HS65_LH_BFX2 U7921 ( .A(n31745), .Z(n31744) );
  HS65_LH_BFX2 U7922 ( .A(n31746), .Z(n31745) );
  HS65_LH_BFX2 U7923 ( .A(n31747), .Z(n31746) );
  HS65_LH_BFX2 U7924 ( .A(n31748), .Z(n31747) );
  HS65_LH_BFX2 U7925 ( .A(n31749), .Z(n31748) );
  HS65_LH_BFX2 U7926 ( .A(n31750), .Z(n31749) );
  HS65_LH_BFX2 U7927 ( .A(n31751), .Z(n31750) );
  HS65_LH_BFX2 U7928 ( .A(n31752), .Z(n31751) );
  HS65_LH_BFX2 U7929 ( .A(n31753), .Z(n31752) );
  HS65_LH_BFX2 U7930 ( .A(n31754), .Z(n31753) );
  HS65_LH_BFX2 U7931 ( .A(n31755), .Z(n31754) );
  HS65_LH_BFX2 U7933 ( .A(n31756), .Z(n31755) );
  HS65_LH_BFX2 U7935 ( .A(n31757), .Z(n31756) );
  HS65_LH_BFX2 U7937 ( .A(n31758), .Z(n31757) );
  HS65_LH_BFX2 U7939 ( .A(n31759), .Z(n31758) );
  HS65_LH_BFX2 U7941 ( .A(n31760), .Z(n31759) );
  HS65_LH_BFX2 U7943 ( .A(n31761), .Z(n31760) );
  HS65_LH_BFX2 U7945 ( .A(n31762), .Z(n31761) );
  HS65_LH_BFX2 U7947 ( .A(n31763), .Z(n31762) );
  HS65_LH_BFX2 U7949 ( .A(n14269), .Z(n31763) );
  HS65_LH_BFX2 U8000 ( .A(n31800), .Z(n31764) );
  HS65_LH_NAND2X7 U8002 ( .A(n16774), .B(n16773), .Z(n16782) );
  HS65_LH_BFX2 U8004 ( .A(n31767), .Z(n31765) );
  HS65_LH_IVX2 U8006 ( .A(n17985), .Z(n31766) );
  HS65_LH_IVX2 U8008 ( .A(n31766), .Z(n31767) );
  HS65_LH_IVX2 U8010 ( .A(n31780), .Z(n31768) );
  HS65_LH_IVX2 U8012 ( .A(n31768), .Z(n31769) );
  HS65_LH_BFX2 U8014 ( .A(n31773), .Z(n31770) );
  HS65_LH_BFX2 U8016 ( .A(n31775), .Z(n31771) );
  HS65_LH_IVX2 U8018 ( .A(n31781), .Z(n31772) );
  HS65_LH_IVX2 U8020 ( .A(n31772), .Z(n31773) );
  HS65_LH_IVX2 U8022 ( .A(n31778), .Z(n31774) );
  HS65_LH_IVX2 U8024 ( .A(n31774), .Z(n31775) );
  HS65_LH_BFX2 U8026 ( .A(n1541), .Z(n31776) );
  HS65_LH_IVX2 U8028 ( .A(n33552), .Z(n31777) );
  HS65_LH_IVX2 U8030 ( .A(n31777), .Z(n31778) );
  HS65_LH_BFX2 U8032 ( .A(n31776), .Z(n31779) );
  HS65_LH_BFX2 U8082 ( .A(n31783), .Z(n31780) );
  HS65_LH_BFX2 U8083 ( .A(n31784), .Z(n31781) );
  HS65_LH_BFX2 U8084 ( .A(n31779), .Z(n31782) );
  HS65_LH_BFX2 U8085 ( .A(n31786), .Z(n31783) );
  HS65_LH_BFX2 U8086 ( .A(n31787), .Z(n31784) );
  HS65_LH_BFX2 U8087 ( .A(n31782), .Z(n31785) );
  HS65_LH_BFX2 U8088 ( .A(n31789), .Z(n31786) );
  HS65_LH_BFX2 U8089 ( .A(n31790), .Z(n31787) );
  HS65_LH_BFX2 U8090 ( .A(n31785), .Z(n31788) );
  HS65_LH_BFX2 U8091 ( .A(n31792), .Z(n31789) );
  HS65_LH_BFX2 U8092 ( .A(n31793), .Z(n31790) );
  HS65_LH_BFX2 U8093 ( .A(n31788), .Z(n31791) );
  HS65_LH_BFX2 U8094 ( .A(n31795), .Z(n31792) );
  HS65_LH_BFX2 U8095 ( .A(n31801), .Z(n31793) );
  HS65_LH_BFX2 U8096 ( .A(n31791), .Z(n31794) );
  HS65_LH_BFX2 U8097 ( .A(n31798), .Z(n31795) );
  HS65_LH_BFX2 U8098 ( .A(n16781), .Z(n31796) );
  HS65_LH_IVX2 U8099 ( .A(n31805), .Z(n31797) );
  HS65_LH_IVX2 U8100 ( .A(n31797), .Z(n31798) );
  HS65_LH_IVX2 U8101 ( .A(n31794), .Z(n31799) );
  HS65_LH_IVX2 U8103 ( .A(n31799), .Z(n31800) );
  HS65_LH_BFX2 U8105 ( .A(n31803), .Z(n31801) );
  HS65_LH_BFX2 U8107 ( .A(n31804), .Z(n31802) );
  HS65_LH_BFX2 U8109 ( .A(n31806), .Z(n31803) );
  HS65_LH_BFX2 U8111 ( .A(n16780), .Z(n31804) );
  HS65_LH_BFX2 U8113 ( .A(n31807), .Z(n31805) );
  HS65_LH_BFX2 U8115 ( .A(n1542), .Z(n31806) );
  HS65_LH_BFX2 U8140 ( .A(n31808), .Z(n31807) );
  HS65_LH_BFX2 U8141 ( .A(n31809), .Z(n31808) );
  HS65_LH_BFX2 U8142 ( .A(n17988), .Z(n31809) );
  HS65_LH_BFX2 U8143 ( .A(n31817), .Z(n31810) );
  HS65_LH_BFX2 U8144 ( .A(n31814), .Z(n31811) );
  HS65_LH_BFX2 U8145 ( .A(n17891), .Z(n31812) );
  HS65_LH_IVX2 U8146 ( .A(n31819), .Z(n31813) );
  HS65_LH_IVX2 U8147 ( .A(n31813), .Z(n31814) );
  HS65_LH_IVX2 U8148 ( .A(n31820), .Z(n31815) );
  HS65_LH_IVX2 U8149 ( .A(n31815), .Z(n31816) );
  HS65_LH_BFX2 U8150 ( .A(n31818), .Z(n31817) );
  HS65_LH_BFX2 U8151 ( .A(n31821), .Z(n31818) );
  HS65_LH_BFX2 U8152 ( .A(n31822), .Z(n31819) );
  HS65_LH_BFX2 U8153 ( .A(n31823), .Z(n31820) );
  HS65_LH_BFX2 U8154 ( .A(n31824), .Z(n31821) );
  HS65_LH_BFX2 U8155 ( .A(n31825), .Z(n31822) );
  HS65_LH_BFX2 U8156 ( .A(n31826), .Z(n31823) );
  HS65_LH_BFX2 U8157 ( .A(n31827), .Z(n31824) );
  HS65_LH_BFX2 U8158 ( .A(n31828), .Z(n31825) );
  HS65_LH_BFX2 U8159 ( .A(n31829), .Z(n31826) );
  HS65_LH_BFX2 U8160 ( .A(n31830), .Z(n31827) );
  HS65_LH_BFX2 U8161 ( .A(n31831), .Z(n31828) );
  HS65_LH_BFX2 U8162 ( .A(n31832), .Z(n31829) );
  HS65_LH_BFX2 U8163 ( .A(n31833), .Z(n31830) );
  HS65_LH_BFX2 U8164 ( .A(n31834), .Z(n31831) );
  HS65_LH_BFX2 U8166 ( .A(n31835), .Z(n31832) );
  HS65_LH_BFX2 U8167 ( .A(n31836), .Z(n31833) );
  HS65_LH_BFX2 U8169 ( .A(n31837), .Z(n31834) );
  HS65_LH_BFX2 U8170 ( .A(n31838), .Z(n31835) );
  HS65_LH_BFX2 U8172 ( .A(n31839), .Z(n31836) );
  HS65_LH_BFX2 U8173 ( .A(n31840), .Z(n31837) );
  HS65_LH_BFX2 U8175 ( .A(n31841), .Z(n31838) );
  HS65_LH_BFX2 U8176 ( .A(n31842), .Z(n31839) );
  HS65_LH_BFX2 U8178 ( .A(n31843), .Z(n31840) );
  HS65_LH_BFX2 U8179 ( .A(n31844), .Z(n31841) );
  HS65_LH_BFX2 U8181 ( .A(n31845), .Z(n31842) );
  HS65_LH_BFX2 U8182 ( .A(n31846), .Z(n31843) );
  HS65_LH_BFX2 U8184 ( .A(n31847), .Z(n31844) );
  HS65_LH_BFX2 U8185 ( .A(n31848), .Z(n31845) );
  HS65_LH_BFX2 U8187 ( .A(n31849), .Z(n31846) );
  HS65_LH_BFX2 U8188 ( .A(n31850), .Z(n31847) );
  HS65_LH_BFX2 U8190 ( .A(n31851), .Z(n31848) );
  HS65_LH_BFX2 U8191 ( .A(n31852), .Z(n31849) );
  HS65_LH_BFX2 U8193 ( .A(n31853), .Z(n31850) );
  HS65_LH_BFX2 U8194 ( .A(n31854), .Z(n31851) );
  HS65_LH_BFX2 U8196 ( .A(n31855), .Z(n31852) );
  HS65_LH_BFX2 U8197 ( .A(n31856), .Z(n31853) );
  HS65_LH_BFX2 U8199 ( .A(n31857), .Z(n31854) );
  HS65_LH_BFX2 U8200 ( .A(n15564), .Z(n31855) );
  HS65_LH_BFX2 U8202 ( .A(n31858), .Z(n31856) );
  HS65_LH_BFX2 U8203 ( .A(n31859), .Z(n31857) );
  HS65_LH_BFX2 U8205 ( .A(n31860), .Z(n31858) );
  HS65_LH_BFX2 U8206 ( .A(n31861), .Z(n31859) );
  HS65_LH_BFX2 U8208 ( .A(n31862), .Z(n31860) );
  HS65_LH_BFX2 U8209 ( .A(n31863), .Z(n31861) );
  HS65_LH_BFX2 U8211 ( .A(n31864), .Z(n31862) );
  HS65_LH_BFX2 U8212 ( .A(n14989), .Z(n31863) );
  HS65_LH_BFX2 U8214 ( .A(n31865), .Z(n31864) );
  HS65_LH_BFX2 U8215 ( .A(n31866), .Z(n31865) );
  HS65_LH_BFX2 U8217 ( .A(n31812), .Z(n31866) );
  HS65_LH_IVX2 U8223 ( .A(n31875), .Z(n31867) );
  HS65_LH_IVX2 U8228 ( .A(n31867), .Z(n31868) );
  HS65_LH_BFX2 U8229 ( .A(n31872), .Z(n31869) );
  HS65_LH_BFX2 U8230 ( .A(n17932), .Z(n31870) );
  HS65_LH_IVX2 U8231 ( .A(n31876), .Z(n31871) );
  HS65_LH_IVX2 U8232 ( .A(n31871), .Z(n31872) );
  HS65_LH_IVX2 U8233 ( .A(n31877), .Z(n31873) );
  HS65_LH_IVX2 U8234 ( .A(n31873), .Z(n31874) );
  HS65_LH_BFX2 U8235 ( .A(n31878), .Z(n31875) );
  HS65_LH_BFX2 U8236 ( .A(n31879), .Z(n31876) );
  HS65_LH_BFX2 U8237 ( .A(n31880), .Z(n31877) );
  HS65_LH_BFX2 U8238 ( .A(n31881), .Z(n31878) );
  HS65_LH_BFX2 U8239 ( .A(n31882), .Z(n31879) );
  HS65_LH_BFX2 U8240 ( .A(n31883), .Z(n31880) );
  HS65_LH_BFX2 U8241 ( .A(n31884), .Z(n31881) );
  HS65_LH_BFX2 U8242 ( .A(n31885), .Z(n31882) );
  HS65_LH_BFX2 U8243 ( .A(n31886), .Z(n31883) );
  HS65_LH_BFX2 U8244 ( .A(n31887), .Z(n31884) );
  HS65_LH_BFX2 U8245 ( .A(n31888), .Z(n31885) );
  HS65_LH_BFX2 U8246 ( .A(n31889), .Z(n31886) );
  HS65_LH_BFX2 U8247 ( .A(n31890), .Z(n31887) );
  HS65_LH_BFX2 U8248 ( .A(n31891), .Z(n31888) );
  HS65_LH_BFX2 U8249 ( .A(n31892), .Z(n31889) );
  HS65_LH_BFX2 U8250 ( .A(n31893), .Z(n31890) );
  HS65_LH_BFX2 U8251 ( .A(n31894), .Z(n31891) );
  HS65_LH_BFX2 U8272 ( .A(n31895), .Z(n31892) );
  HS65_LH_BFX2 U8273 ( .A(n31896), .Z(n31893) );
  HS65_LH_BFX2 U8274 ( .A(n31897), .Z(n31894) );
  HS65_LH_BFX2 U8275 ( .A(n31898), .Z(n31895) );
  HS65_LH_BFX2 U8276 ( .A(n31899), .Z(n31896) );
  HS65_LH_BFX2 U8277 ( .A(n31900), .Z(n31897) );
  HS65_LH_BFX2 U8278 ( .A(n31901), .Z(n31898) );
  HS65_LH_BFX2 U8279 ( .A(n31902), .Z(n31899) );
  HS65_LH_BFX2 U8280 ( .A(n31903), .Z(n31900) );
  HS65_LH_BFX2 U8281 ( .A(n31904), .Z(n31901) );
  HS65_LH_BFX2 U8282 ( .A(n31905), .Z(n31902) );
  HS65_LH_BFX2 U8283 ( .A(n31906), .Z(n31903) );
  HS65_LH_BFX2 U8284 ( .A(n31907), .Z(n31904) );
  HS65_LH_BFX2 U8285 ( .A(n31908), .Z(n31905) );
  HS65_LH_BFX2 U8286 ( .A(n31909), .Z(n31906) );
  HS65_LH_BFX2 U8297 ( .A(n31910), .Z(n31907) );
  HS65_LH_BFX2 U8298 ( .A(n31913), .Z(n31908) );
  HS65_LH_BFX2 U8300 ( .A(n31912), .Z(n31909) );
  HS65_LH_BFX2 U8301 ( .A(n31914), .Z(n31910) );
  HS65_LH_IVX2 U8303 ( .A(n31916), .Z(n31911) );
  HS65_LH_IVX2 U8304 ( .A(n31911), .Z(n31912) );
  HS65_LH_BFX2 U8306 ( .A(n31917), .Z(n31913) );
  HS65_LH_BFX2 U8307 ( .A(n31918), .Z(n31914) );
  HS65_LH_IVX2 U8309 ( .A(n15562), .Z(n31915) );
  HS65_LH_IVX2 U8310 ( .A(n31915), .Z(n31916) );
  HS65_LH_BFX2 U8312 ( .A(n31919), .Z(n31917) );
  HS65_LH_BFX2 U8313 ( .A(n31920), .Z(n31918) );
  HS65_LH_BFX2 U8315 ( .A(n31921), .Z(n31919) );
  HS65_LH_BFX2 U8316 ( .A(n31922), .Z(n31920) );
  HS65_LH_BFX2 U8318 ( .A(n31923), .Z(n31921) );
  HS65_LH_BFX2 U8320 ( .A(n31924), .Z(n31922) );
  HS65_LH_BFX2 U8321 ( .A(n31925), .Z(n31923) );
  HS65_LH_BFX2 U8323 ( .A(n31926), .Z(n31924) );
  HS65_LH_BFX2 U8324 ( .A(n14697), .Z(n31925) );
  HS65_LH_BFX2 U8326 ( .A(n31927), .Z(n31926) );
  HS65_LH_BFX2 U8327 ( .A(n31870), .Z(n31927) );
  HS65_LH_BFX2 U8329 ( .A(n33965), .Z(n31928) );
  HS65_LH_BFX2 U8330 ( .A(n33964), .Z(n31929) );
  HS65_LH_BFX2 U8332 ( .A(n31931), .Z(n31930) );
  HS65_LH_BFX2 U8333 ( .A(n31932), .Z(n31931) );
  HS65_LH_BFX2 U8335 ( .A(n31933), .Z(n31932) );
  HS65_LH_BFX2 U8336 ( .A(n31934), .Z(n31933) );
  HS65_LH_BFX2 U8338 ( .A(n31935), .Z(n31934) );
  HS65_LH_BFX2 U8339 ( .A(n31936), .Z(n31935) );
  HS65_LH_BFX2 U8341 ( .A(n31937), .Z(n31936) );
  HS65_LH_BFX2 U8342 ( .A(n31938), .Z(n31937) );
  HS65_LH_BFX2 U8344 ( .A(n31939), .Z(n31938) );
  HS65_LH_BFX2 U8345 ( .A(n31940), .Z(n31939) );
  HS65_LH_BFX2 U8347 ( .A(n31941), .Z(n31940) );
  HS65_LH_BFX2 U8348 ( .A(n31942), .Z(n31941) );
  HS65_LH_BFX2 U8350 ( .A(n31943), .Z(n31942) );
  HS65_LH_BFX2 U8352 ( .A(n31944), .Z(n31943) );
  HS65_LH_BFX2 U8354 ( .A(n31945), .Z(n31944) );
  HS65_LH_BFX2 U8405 ( .A(n31946), .Z(n31945) );
  HS65_LH_BFX2 U8407 ( .A(n31947), .Z(n31946) );
  HS65_LH_BFX2 U8409 ( .A(n31948), .Z(n31947) );
  HS65_LH_BFX2 U8411 ( .A(n31949), .Z(n31948) );
  HS65_LH_BFX2 U8413 ( .A(n31950), .Z(n31949) );
  HS65_LH_BFX2 U8415 ( .A(n14275), .Z(n31950) );
  HS65_LH_BFX2 U8417 ( .A(n31952), .Z(n31951) );
  HS65_LH_BFX2 U8419 ( .A(n31953), .Z(n31952) );
  HS65_LH_BFX2 U8421 ( .A(n31954), .Z(n31953) );
  HS65_LH_BFX2 U8423 ( .A(n31955), .Z(n31954) );
  HS65_LH_BFX2 U8425 ( .A(n31956), .Z(n31955) );
  HS65_LH_BFX2 U8429 ( .A(n31957), .Z(n31956) );
  HS65_LH_BFX2 U8431 ( .A(n31958), .Z(n31957) );
  HS65_LH_BFX2 U8433 ( .A(n31959), .Z(n31958) );
  HS65_LH_BFX2 U8435 ( .A(n31960), .Z(n31959) );
  HS65_LH_BFX2 U8437 ( .A(n31961), .Z(n31960) );
  HS65_LH_BFX2 U8462 ( .A(n31962), .Z(n31961) );
  HS65_LH_BFX2 U8463 ( .A(n31963), .Z(n31962) );
  HS65_LH_BFX2 U8464 ( .A(n31964), .Z(n31963) );
  HS65_LH_BFX2 U8465 ( .A(n31965), .Z(n31964) );
  HS65_LH_BFX2 U8466 ( .A(n31966), .Z(n31965) );
  HS65_LH_BFX2 U8467 ( .A(n31967), .Z(n31966) );
  HS65_LH_BFX2 U8468 ( .A(n31968), .Z(n31967) );
  HS65_LH_BFX2 U8469 ( .A(n31969), .Z(n31968) );
  HS65_LH_BFX2 U8470 ( .A(n31970), .Z(n31969) );
  HS65_LH_BFX2 U8471 ( .A(n31971), .Z(n31970) );
  HS65_LH_BFX2 U8472 ( .A(n14270), .Z(n31971) );
  HS65_LH_BFX2 U8473 ( .A(n31973), .Z(n31972) );
  HS65_LH_BFX2 U8474 ( .A(n31974), .Z(n31973) );
  HS65_LH_BFX2 U8475 ( .A(n31975), .Z(n31974) );
  HS65_LH_BFX2 U8476 ( .A(n31976), .Z(n31975) );
  HS65_LH_BFX2 U8477 ( .A(n31977), .Z(n31976) );
  HS65_LH_BFX2 U8478 ( .A(n31978), .Z(n31977) );
  HS65_LH_BFX2 U8479 ( .A(n31979), .Z(n31978) );
  HS65_LH_BFX2 U8480 ( .A(n31980), .Z(n31979) );
  HS65_LH_BFX2 U8481 ( .A(n31981), .Z(n31980) );
  HS65_LH_BFX2 U8482 ( .A(n31982), .Z(n31981) );
  HS65_LH_BFX2 U8483 ( .A(n31983), .Z(n31982) );
  HS65_LH_BFX2 U8484 ( .A(n31984), .Z(n31983) );
  HS65_LH_BFX2 U8485 ( .A(n31985), .Z(n31984) );
  HS65_LH_BFX2 U8486 ( .A(n31986), .Z(n31985) );
  HS65_LH_BFX2 U8487 ( .A(n31987), .Z(n31986) );
  HS65_LH_BFX2 U8488 ( .A(n31988), .Z(n31987) );
  HS65_LH_BFX2 U8490 ( .A(n31989), .Z(n31988) );
  HS65_LH_BFX2 U8493 ( .A(n31990), .Z(n31989) );
  HS65_LH_BFX2 U8494 ( .A(n31991), .Z(n31990) );
  HS65_LH_BFX2 U8496 ( .A(n31992), .Z(n31991) );
  HS65_LH_BFX2 U8497 ( .A(n14222), .Z(n31992) );
  HS65_LH_BFX2 U8499 ( .A(n32005), .Z(n31993) );
  HS65_LH_BFX2 U8500 ( .A(n31995), .Z(n31994) );
  HS65_LH_BFX2 U8502 ( .A(n31996), .Z(n31995) );
  HS65_LH_BFX2 U8503 ( .A(n31997), .Z(n31996) );
  HS65_LH_BFX2 U8505 ( .A(n31998), .Z(n31997) );
  HS65_LH_BFX2 U8507 ( .A(n31999), .Z(n31998) );
  HS65_LH_BFX2 U8508 ( .A(n32000), .Z(n31999) );
  HS65_LH_BFX2 U8510 ( .A(n32001), .Z(n32000) );
  HS65_LH_BFX2 U8511 ( .A(n32002), .Z(n32001) );
  HS65_LH_BFX2 U8513 ( .A(n32003), .Z(n32002) );
  HS65_LH_BFX2 U8514 ( .A(n32004), .Z(n32003) );
  HS65_LH_BFX2 U8516 ( .A(n31993), .Z(n32004) );
  HS65_LH_BFX2 U8517 ( .A(n32006), .Z(n32005) );
  HS65_LH_BFX2 U8519 ( .A(n32007), .Z(n32006) );
  HS65_LH_BFX2 U8520 ( .A(n32008), .Z(n32007) );
  HS65_LH_BFX2 U8522 ( .A(n32009), .Z(n32008) );
  HS65_LH_BFX2 U8523 ( .A(n32010), .Z(n32009) );
  HS65_LH_BFX2 U8525 ( .A(n32011), .Z(n32010) );
  HS65_LH_BFX2 U8526 ( .A(n32012), .Z(n32011) );
  HS65_LH_BFX2 U8528 ( .A(n32013), .Z(n32012) );
  HS65_LH_BFX2 U8529 ( .A(n14215), .Z(n32013) );
  HS65_LH_BFX2 U8531 ( .A(n32015), .Z(n32014) );
  HS65_LH_BFX2 U8532 ( .A(n32016), .Z(n32015) );
  HS65_LH_BFX2 U8534 ( .A(n32017), .Z(n32016) );
  HS65_LH_BFX2 U8535 ( .A(n32018), .Z(n32017) );
  HS65_LH_BFX2 U8537 ( .A(n32019), .Z(n32018) );
  HS65_LH_BFX2 U8538 ( .A(n32020), .Z(n32019) );
  HS65_LH_BFX2 U8540 ( .A(n32021), .Z(n32020) );
  HS65_LH_BFX2 U8541 ( .A(n32022), .Z(n32021) );
  HS65_LH_BFX2 U8543 ( .A(n32023), .Z(n32022) );
  HS65_LH_BFX2 U8545 ( .A(n32024), .Z(n32023) );
  HS65_LH_BFX2 U8595 ( .A(n32025), .Z(n32024) );
  HS65_LH_BFX2 U8597 ( .A(n32026), .Z(n32025) );
  HS65_LH_BFX2 U8599 ( .A(n32027), .Z(n32026) );
  HS65_LH_BFX2 U8601 ( .A(n32028), .Z(n32027) );
  HS65_LH_BFX2 U8603 ( .A(n32029), .Z(n32028) );
  HS65_LH_BFX2 U8605 ( .A(n32030), .Z(n32029) );
  HS65_LH_BFX2 U8607 ( .A(n32031), .Z(n32030) );
  HS65_LH_BFX2 U8609 ( .A(n32032), .Z(n32031) );
  HS65_LH_BFX2 U8611 ( .A(n32033), .Z(n32032) );
  HS65_LH_BFX2 U8613 ( .A(n32034), .Z(n32033) );
  HS65_LH_BFX2 U8615 ( .A(n32035), .Z(n32034) );
  HS65_LH_BFX2 U8617 ( .A(n17259), .Z(n32035) );
  HS65_LH_BFX2 U8619 ( .A(n32037), .Z(n32036) );
  HS65_LH_BFX2 U8621 ( .A(n32038), .Z(n32037) );
  HS65_LH_BFX2 U8623 ( .A(n32039), .Z(n32038) );
  HS65_LH_BFX2 U8625 ( .A(n32040), .Z(n32039) );
  HS65_LH_BFX2 U8627 ( .A(n32041), .Z(n32040) );
  HS65_LH_BFX2 U8629 ( .A(n32042), .Z(n32041) );
  HS65_LH_BFX2 U8631 ( .A(n32043), .Z(n32042) );
  HS65_LH_BFX2 U8655 ( .A(n32044), .Z(n32043) );
  HS65_LH_BFX2 U8656 ( .A(n32045), .Z(n32044) );
  HS65_LH_BFX2 U8657 ( .A(n32046), .Z(n32045) );
  HS65_LH_BFX2 U8658 ( .A(n32047), .Z(n32046) );
  HS65_LH_BFX2 U8659 ( .A(n32048), .Z(n32047) );
  HS65_LH_BFX2 U8660 ( .A(n32049), .Z(n32048) );
  HS65_LH_BFX2 U8661 ( .A(n32050), .Z(n32049) );
  HS65_LH_BFX2 U8662 ( .A(n32051), .Z(n32050) );
  HS65_LH_BFX2 U8663 ( .A(n32052), .Z(n32051) );
  HS65_LH_BFX2 U8664 ( .A(n32053), .Z(n32052) );
  HS65_LH_BFX2 U8665 ( .A(n32054), .Z(n32053) );
  HS65_LH_BFX2 U8666 ( .A(n32055), .Z(n32054) );
  HS65_LH_BFX2 U8667 ( .A(n32056), .Z(n32055) );
  HS65_LH_BFX2 U8668 ( .A(n32504), .Z(n32056) );
  HS65_LH_BFX2 U8669 ( .A(n32058), .Z(n32057) );
  HS65_LH_BFX2 U8670 ( .A(n32059), .Z(n32058) );
  HS65_LH_BFX2 U8671 ( .A(n32060), .Z(n32059) );
  HS65_LH_BFX2 U8672 ( .A(n32061), .Z(n32060) );
  HS65_LH_BFX2 U8673 ( .A(n32062), .Z(n32061) );
  HS65_LH_BFX2 U8674 ( .A(n32063), .Z(n32062) );
  HS65_LH_BFX2 U8675 ( .A(n32064), .Z(n32063) );
  HS65_LH_BFX2 U8676 ( .A(n32065), .Z(n32064) );
  HS65_LH_BFX2 U8677 ( .A(n32066), .Z(n32065) );
  HS65_LH_BFX2 U8678 ( .A(n32067), .Z(n32066) );
  HS65_LH_BFX2 U8679 ( .A(n32068), .Z(n32067) );
  HS65_LH_BFX2 U8680 ( .A(n32069), .Z(n32068) );
  HS65_LH_BFX2 U8681 ( .A(n32070), .Z(n32069) );
  HS65_LH_BFX2 U8683 ( .A(n32071), .Z(n32070) );
  HS65_LH_BFX2 U8684 ( .A(n32072), .Z(n32071) );
  HS65_LH_BFX2 U8686 ( .A(n32073), .Z(n32072) );
  HS65_LH_BFX2 U8687 ( .A(n32074), .Z(n32073) );
  HS65_LH_BFX2 U8689 ( .A(n32075), .Z(n32074) );
  HS65_LH_BFX2 U8690 ( .A(n32076), .Z(n32075) );
  HS65_LH_BFX2 U8692 ( .A(n32077), .Z(n32076) );
  HS65_LH_BFX2 U8693 ( .A(n32078), .Z(n32077) );
  HS65_LH_BFX2 U8695 ( .A(n17258), .Z(n32078) );
  HS65_LH_BFX2 U8696 ( .A(n32080), .Z(n32079) );
  HS65_LH_BFX2 U8698 ( .A(n32081), .Z(n32080) );
  HS65_LH_BFX2 U8699 ( .A(n32082), .Z(n32081) );
  HS65_LH_BFX2 U8701 ( .A(n32083), .Z(n32082) );
  HS65_LH_BFX2 U8702 ( .A(n32084), .Z(n32083) );
  HS65_LH_BFX2 U8704 ( .A(n32085), .Z(n32084) );
  HS65_LH_BFX2 U8705 ( .A(n32086), .Z(n32085) );
  HS65_LH_BFX2 U8707 ( .A(n32087), .Z(n32086) );
  HS65_LH_BFX2 U8708 ( .A(n32088), .Z(n32087) );
  HS65_LH_BFX2 U8710 ( .A(n32089), .Z(n32088) );
  HS65_LH_BFX2 U8711 ( .A(n32090), .Z(n32089) );
  HS65_LH_BFX2 U8713 ( .A(n32091), .Z(n32090) );
  HS65_LH_BFX2 U8714 ( .A(n32092), .Z(n32091) );
  HS65_LH_BFX2 U8716 ( .A(n32093), .Z(n32092) );
  HS65_LH_BFX2 U8717 ( .A(n32094), .Z(n32093) );
  HS65_LH_BFX2 U8719 ( .A(n32095), .Z(n32094) );
  HS65_LH_BFX2 U8720 ( .A(n32097), .Z(n32095) );
  HS65_LH_BFX2 U8722 ( .A(n14250), .Z(n32096) );
  HS65_LH_BFX2 U8723 ( .A(n15574), .Z(n32097) );
  HS65_LH_IVX2 U8725 ( .A(n32102), .Z(n32098) );
  HS65_LH_IVX2 U8727 ( .A(n32098), .Z(n32099) );
  HS65_LH_IVX2 U8728 ( .A(n17331), .Z(n32100) );
  HS65_LH_IVX2 U8730 ( .A(n32100), .Z(n32101) );
  HS65_LH_BFX2 U8731 ( .A(n32103), .Z(n32102) );
  HS65_LH_BFX2 U8733 ( .A(n32104), .Z(n32103) );
  HS65_LH_BFX2 U8735 ( .A(n32105), .Z(n32104) );
  HS65_LH_BFX2 U8737 ( .A(n32106), .Z(n32105) );
  HS65_LH_BFX2 U8762 ( .A(n32107), .Z(n32106) );
  HS65_LH_BFX2 U8763 ( .A(n32108), .Z(n32107) );
  HS65_LH_BFX2 U8764 ( .A(n32109), .Z(n32108) );
  HS65_LH_BFX2 U8765 ( .A(n32110), .Z(n32109) );
  HS65_LH_BFX2 U8766 ( .A(n32111), .Z(n32110) );
  HS65_LH_BFX2 U8767 ( .A(n32112), .Z(n32111) );
  HS65_LH_BFX2 U8768 ( .A(n32113), .Z(n32112) );
  HS65_LH_BFX2 U8769 ( .A(n32114), .Z(n32113) );
  HS65_LH_BFX2 U8770 ( .A(n32115), .Z(n32114) );
  HS65_LH_BFX2 U8771 ( .A(n32116), .Z(n32115) );
  HS65_LH_BFX2 U8772 ( .A(n32117), .Z(n32116) );
  HS65_LH_BFX2 U8773 ( .A(n32118), .Z(n32117) );
  HS65_LH_BFX2 U8774 ( .A(n14513), .Z(n32118) );
  HS65_LH_IVX2 U8775 ( .A(n32121), .Z(n32119) );
  HS65_LH_IVX2 U8776 ( .A(n32119), .Z(n32120) );
  HS65_LH_BFX2 U8777 ( .A(n32122), .Z(n32121) );
  HS65_LH_BFX2 U8778 ( .A(n32123), .Z(n32122) );
  HS65_LH_BFX2 U8779 ( .A(n32124), .Z(n32123) );
  HS65_LH_BFX2 U8780 ( .A(n32125), .Z(n32124) );
  HS65_LH_BFX2 U8781 ( .A(n32126), .Z(n32125) );
  HS65_LH_BFX2 U8782 ( .A(n32127), .Z(n32126) );
  HS65_LH_BFX2 U8783 ( .A(n32128), .Z(n32127) );
  HS65_LH_BFX2 U8784 ( .A(n32129), .Z(n32128) );
  HS65_LH_BFX2 U8785 ( .A(n32130), .Z(n32129) );
  HS65_LH_BFX2 U8786 ( .A(n32131), .Z(n32130) );
  HS65_LH_BFX2 U8790 ( .A(n32132), .Z(n32131) );
  HS65_LH_BFX2 U8792 ( .A(n32133), .Z(n32132) );
  HS65_LH_BFX2 U8793 ( .A(n40558), .Z(n32133) );
  HS65_LH_BFX2 U8795 ( .A(n32135), .Z(n32134) );
  HS65_LH_BFX2 U8796 ( .A(n32136), .Z(n32135) );
  HS65_LH_BFX2 U8798 ( .A(n17341), .Z(n32136) );
  HS65_LH_BFX2 U8799 ( .A(n32138), .Z(n32137) );
  HS65_LH_BFX2 U8801 ( .A(n32139), .Z(n32138) );
  HS65_LH_BFX2 U8802 ( .A(n32140), .Z(n32139) );
  HS65_LH_BFX2 U8804 ( .A(n32141), .Z(n32140) );
  HS65_LH_BFX2 U8805 ( .A(n32142), .Z(n32141) );
  HS65_LH_BFX2 U8807 ( .A(n32143), .Z(n32142) );
  HS65_LH_BFX2 U8808 ( .A(n32144), .Z(n32143) );
  HS65_LH_BFX2 U8810 ( .A(n32145), .Z(n32144) );
  HS65_LH_BFX2 U8811 ( .A(n32146), .Z(n32145) );
  HS65_LH_BFX2 U8813 ( .A(n32147), .Z(n32146) );
  HS65_LH_BFX2 U8814 ( .A(n32148), .Z(n32147) );
  HS65_LH_BFX2 U8816 ( .A(n32149), .Z(n32148) );
  HS65_LH_BFX2 U8817 ( .A(n32150), .Z(n32149) );
  HS65_LH_BFX2 U8819 ( .A(n32151), .Z(n32150) );
  HS65_LH_BFX2 U8820 ( .A(n32154), .Z(n32151) );
  HS65_LH_BFX2 U8822 ( .A(n32153), .Z(n32152) );
  HS65_LH_BFX2 U8823 ( .A(n14477), .Z(n32153) );
  HS65_LH_BFX2 U8825 ( .A(n15573), .Z(n32154) );
  HS65_LH_IVX2 U8826 ( .A(n32161), .Z(n32155) );
  HS65_LH_IVX2 U8828 ( .A(n32155), .Z(n32156) );
  HS65_LH_BFX2 U8829 ( .A(n32159), .Z(n32157) );
  HS65_LH_BFX2 U8831 ( .A(n32160), .Z(n32158) );
  HS65_LH_BFX2 U8832 ( .A(n32162), .Z(n32159) );
  HS65_LH_BFX2 U8834 ( .A(n32163), .Z(n32160) );
  HS65_LH_BFX2 U8835 ( .A(n32164), .Z(n32161) );
  HS65_LH_BFX2 U8837 ( .A(n32165), .Z(n32162) );
  HS65_LH_BFX2 U8838 ( .A(n32166), .Z(n32163) );
  HS65_LH_BFX2 U8840 ( .A(n32167), .Z(n32164) );
  HS65_LH_BFX2 U8842 ( .A(n32168), .Z(n32165) );
  HS65_LH_BFX2 U8844 ( .A(n32169), .Z(n32166) );
  HS65_LH_BFX2 U8846 ( .A(n32170), .Z(n32167) );
  HS65_LH_BFX2 U8871 ( .A(n32171), .Z(n32168) );
  HS65_LH_BFX2 U8872 ( .A(n32172), .Z(n32169) );
  HS65_LH_BFX2 U8873 ( .A(n32173), .Z(n32170) );
  HS65_LH_BFX2 U8874 ( .A(n32174), .Z(n32171) );
  HS65_LH_BFX2 U8875 ( .A(n32175), .Z(n32172) );
  HS65_LH_BFX2 U8876 ( .A(n32176), .Z(n32173) );
  HS65_LH_BFX2 U8877 ( .A(n32177), .Z(n32174) );
  HS65_LH_BFX2 U8878 ( .A(n32178), .Z(n32175) );
  HS65_LH_BFX2 U8879 ( .A(n32179), .Z(n32176) );
  HS65_LH_BFX2 U8880 ( .A(n32180), .Z(n32177) );
  HS65_LH_BFX2 U8881 ( .A(n32181), .Z(n32178) );
  HS65_LH_BFX2 U8882 ( .A(n32182), .Z(n32179) );
  HS65_LH_BFX2 U8883 ( .A(n32183), .Z(n32180) );
  HS65_LH_BFX2 U8884 ( .A(n32184), .Z(n32181) );
  HS65_LH_BFX2 U8885 ( .A(n32185), .Z(n32182) );
  HS65_LH_BFX2 U8886 ( .A(n32186), .Z(n32183) );
  HS65_LH_BFX2 U8887 ( .A(n32187), .Z(n32184) );
  HS65_LH_BFX2 U8888 ( .A(n32188), .Z(n32185) );
  HS65_LH_BFX2 U8889 ( .A(n32189), .Z(n32186) );
  HS65_LH_BFX2 U8890 ( .A(n32190), .Z(n32187) );
  HS65_LH_BFX2 U8891 ( .A(n32191), .Z(n32188) );
  HS65_LH_BFX2 U8892 ( .A(n32192), .Z(n32189) );
  HS65_LH_BFX2 U8899 ( .A(n32193), .Z(n32190) );
  HS65_LH_BFX2 U8901 ( .A(n32194), .Z(n32191) );
  HS65_LH_BFX2 U8902 ( .A(n32195), .Z(n32192) );
  HS65_LH_BFX2 U8904 ( .A(n32196), .Z(n32193) );
  HS65_LH_BFX2 U8905 ( .A(n32197), .Z(n32194) );
  HS65_LH_BFX2 U8907 ( .A(n32198), .Z(n32195) );
  HS65_LH_BFX2 U8908 ( .A(n32199), .Z(n32196) );
  HS65_LH_BFX2 U8910 ( .A(n32200), .Z(n32197) );
  HS65_LH_BFX2 U8911 ( .A(n32201), .Z(n32198) );
  HS65_LH_BFX2 U8913 ( .A(n15558), .Z(n32199) );
  HS65_LH_BFX2 U8914 ( .A(n32202), .Z(n32200) );
  HS65_LH_BFX2 U8916 ( .A(n32203), .Z(n32201) );
  HS65_LH_BFX2 U8917 ( .A(n32204), .Z(n32202) );
  HS65_LH_BFX2 U8919 ( .A(n32205), .Z(n32203) );
  HS65_LH_BFX2 U8920 ( .A(n32206), .Z(n32204) );
  HS65_LH_BFX2 U8922 ( .A(n32207), .Z(n32205) );
  HS65_LH_BFX2 U8923 ( .A(n32208), .Z(n32206) );
  HS65_LH_BFX2 U8925 ( .A(n32209), .Z(n32207) );
  HS65_LH_BFX2 U8926 ( .A(n14381), .Z(n32208) );
  HS65_LH_BFX2 U8928 ( .A(n32210), .Z(n32209) );
  HS65_LH_BFX2 U8929 ( .A(n17975), .Z(n32210) );
  HS65_LH_IVX2 U8931 ( .A(n32215), .Z(n32211) );
  HS65_LH_IVX2 U8932 ( .A(n32211), .Z(n32212) );
  HS65_LH_IVX2 U8934 ( .A(n32231), .Z(n32213) );
  HS65_LH_IVX2 U8935 ( .A(n32213), .Z(n32214) );
  HS65_LH_BFX2 U8937 ( .A(n32216), .Z(n32215) );
  HS65_LH_BFX2 U8938 ( .A(n32217), .Z(n32216) );
  HS65_LH_BFX2 U8940 ( .A(n32218), .Z(n32217) );
  HS65_LH_BFX2 U8941 ( .A(n32219), .Z(n32218) );
  HS65_LH_BFX2 U8943 ( .A(n32220), .Z(n32219) );
  HS65_LH_BFX2 U8944 ( .A(n32221), .Z(n32220) );
  HS65_LH_BFX2 U8946 ( .A(n32222), .Z(n32221) );
  HS65_LH_BFX2 U8948 ( .A(n32223), .Z(n32222) );
  HS65_LH_BFX2 U8950 ( .A(n32224), .Z(n32223) );
  HS65_LH_BFX2 U8952 ( .A(n32225), .Z(n32224) );
  HS65_LH_BFX2 U8954 ( .A(n32226), .Z(n32225) );
  HS65_LH_BFX2 U8959 ( .A(n32227), .Z(n32226) );
  HS65_LH_BFX2 U8960 ( .A(n32228), .Z(n32227) );
  HS65_LH_BFX2 U8961 ( .A(n32229), .Z(n32228) );
  HS65_LH_BFX2 U8962 ( .A(n32230), .Z(n32229) );
  HS65_LH_BFX2 U8963 ( .A(n14251), .Z(n32230) );
  HS65_LH_BFX2 U8964 ( .A(n32232), .Z(n32231) );
  HS65_LH_BFX2 U8965 ( .A(n17332), .Z(n32232) );
  HS65_LH_IVX2 U8966 ( .A(n32237), .Z(n32233) );
  HS65_LH_IVX2 U8967 ( .A(n32233), .Z(n32234) );
  HS65_LH_IVX2 U8968 ( .A(n17329), .Z(n32235) );
  HS65_LH_IVX2 U8969 ( .A(n32235), .Z(n32236) );
  HS65_LH_BFX2 U8970 ( .A(n32238), .Z(n32237) );
  HS65_LH_BFX2 U8971 ( .A(n32239), .Z(n32238) );
  HS65_LH_BFX2 U8972 ( .A(n32240), .Z(n32239) );
  HS65_LH_BFX2 U8973 ( .A(n32241), .Z(n32240) );
  HS65_LH_BFX2 U8974 ( .A(n32242), .Z(n32241) );
  HS65_LH_BFX2 U8975 ( .A(n32243), .Z(n32242) );
  HS65_LH_BFX2 U8976 ( .A(n32244), .Z(n32243) );
  HS65_LH_BFX2 U8977 ( .A(n32245), .Z(n32244) );
  HS65_LH_BFX2 U8978 ( .A(n32246), .Z(n32245) );
  HS65_LH_BFX2 U8979 ( .A(n32247), .Z(n32246) );
  HS65_LH_BFX2 U8980 ( .A(n32248), .Z(n32247) );
  HS65_LH_BFX2 U8981 ( .A(n32249), .Z(n32248) );
  HS65_LH_BFX2 U8982 ( .A(n32250), .Z(n32249) );
  HS65_LH_BFX2 U8983 ( .A(n32251), .Z(n32250) );
  HS65_LH_BFX2 U8984 ( .A(n32252), .Z(n32251) );
  HS65_LH_BFX2 U8985 ( .A(n32253), .Z(n32252) );
  HS65_LH_BFX2 U8986 ( .A(n32254), .Z(n32253) );
  HS65_LH_BFX2 U8987 ( .A(n14252), .Z(n32254) );
  HS65_LH_IVX2 U8988 ( .A(n32259), .Z(n32255) );
  HS65_LH_IVX2 U8989 ( .A(n32255), .Z(n32256) );
  HS65_LH_IVX2 U8990 ( .A(n17340), .Z(n32257) );
  HS65_LH_IVX2 U8991 ( .A(n32257), .Z(n32258) );
  HS65_LH_BFX2 U8992 ( .A(n32260), .Z(n32259) );
  HS65_LH_BFX2 U8993 ( .A(n32261), .Z(n32260) );
  HS65_LH_BFX2 U8994 ( .A(n32262), .Z(n32261) );
  HS65_LH_BFX2 U8995 ( .A(n32263), .Z(n32262) );
  HS65_LH_BFX2 U8996 ( .A(n32264), .Z(n32263) );
  HS65_LH_BFX2 U8997 ( .A(n32265), .Z(n32264) );
  HS65_LH_BFX2 U8999 ( .A(n32266), .Z(n32265) );
  HS65_LH_BFX2 U9001 ( .A(n32267), .Z(n32266) );
  HS65_LH_BFX2 U9003 ( .A(n32268), .Z(n32267) );
  HS65_LH_BFX2 U9005 ( .A(n32269), .Z(n32268) );
  HS65_LH_BFX2 U9007 ( .A(n32270), .Z(n32269) );
  HS65_LH_BFX2 U9009 ( .A(n32271), .Z(n32270) );
  HS65_LH_BFX2 U9011 ( .A(n32272), .Z(n32271) );
  HS65_LH_BFX2 U9013 ( .A(n32273), .Z(n32272) );
  HS65_LH_BFX2 U9015 ( .A(n32274), .Z(n32273) );
  HS65_LH_BFX2 U9017 ( .A(n32275), .Z(n32274) );
  HS65_LH_BFX2 U9020 ( .A(n32276), .Z(n32275) );
  HS65_LH_BFX2 U9021 ( .A(n14253), .Z(n32276) );
  HS65_LH_BFX2 U9071 ( .A(n32279), .Z(n32277) );
  HS65_LH_IVX2 U9073 ( .A(n32282), .Z(n32278) );
  HS65_LH_IVX2 U9075 ( .A(n32278), .Z(n32279) );
  HS65_LH_IVX2 U9077 ( .A(n17333), .Z(n32280) );
  HS65_LH_IVX2 U9079 ( .A(n32280), .Z(n32281) );
  HS65_LH_BFX2 U9081 ( .A(n32283), .Z(n32282) );
  HS65_LH_BFX2 U9083 ( .A(n32284), .Z(n32283) );
  HS65_LH_BFX2 U9085 ( .A(n32285), .Z(n32284) );
  HS65_LH_BFX2 U9087 ( .A(n32286), .Z(n32285) );
  HS65_LH_BFX2 U9089 ( .A(n32287), .Z(n32286) );
  HS65_LH_BFX2 U9091 ( .A(n32288), .Z(n32287) );
  HS65_LH_BFX2 U9093 ( .A(n32289), .Z(n32288) );
  HS65_LH_BFX2 U9095 ( .A(n32290), .Z(n32289) );
  HS65_LH_BFX2 U9097 ( .A(n32291), .Z(n32290) );
  HS65_LH_BFX2 U9099 ( .A(n32292), .Z(n32291) );
  HS65_LH_BFX2 U9101 ( .A(n32293), .Z(n32292) );
  HS65_LH_BFX2 U9103 ( .A(n32294), .Z(n32293) );
  HS65_LH_BFX2 U9109 ( .A(n32295), .Z(n32294) );
  HS65_LH_BFX2 U9110 ( .A(n32296), .Z(n32295) );
  HS65_LH_BFX2 U9112 ( .A(n32297), .Z(n32296) );
  HS65_LH_BFX2 U9114 ( .A(n32298), .Z(n32297) );
  HS65_LH_BFX2 U9117 ( .A(n32299), .Z(n32298) );
  HS65_LH_BFX2 U9119 ( .A(n14254), .Z(n32299) );
  HS65_LH_BFX2 U9121 ( .A(n32302), .Z(n32300) );
  HS65_LH_IVX2 U9123 ( .A(n32305), .Z(n32301) );
  HS65_LH_IVX2 U9164 ( .A(n32301), .Z(n32302) );
  HS65_LH_IVX2 U9165 ( .A(n17338), .Z(n32303) );
  HS65_LH_IVX2 U9167 ( .A(n32303), .Z(n32304) );
  HS65_LH_BFX2 U9169 ( .A(n32306), .Z(n32305) );
  HS65_LH_BFX2 U9171 ( .A(n32307), .Z(n32306) );
  HS65_LH_BFX2 U9173 ( .A(n32308), .Z(n32307) );
  HS65_LH_BFX2 U9175 ( .A(n32309), .Z(n32308) );
  HS65_LH_BFX2 U9177 ( .A(n32310), .Z(n32309) );
  HS65_LH_BFX2 U9179 ( .A(n32311), .Z(n32310) );
  HS65_LH_BFX2 U9181 ( .A(n32312), .Z(n32311) );
  HS65_LH_BFX2 U9183 ( .A(n32313), .Z(n32312) );
  HS65_LH_BFX2 U9185 ( .A(n32314), .Z(n32313) );
  HS65_LH_BFX2 U9187 ( .A(n32315), .Z(n32314) );
  HS65_LH_BFX2 U9189 ( .A(n32316), .Z(n32315) );
  HS65_LH_BFX2 U9191 ( .A(n32317), .Z(n32316) );
  HS65_LH_BFX2 U9193 ( .A(n32318), .Z(n32317) );
  HS65_LH_BFX2 U9195 ( .A(n32319), .Z(n32318) );
  HS65_LH_BFX2 U9197 ( .A(n32320), .Z(n32319) );
  HS65_LH_BFX2 U9222 ( .A(n32321), .Z(n32320) );
  HS65_LH_BFX2 U9223 ( .A(n32322), .Z(n32321) );
  HS65_LH_BFX2 U9224 ( .A(n14243), .Z(n32322) );
  HS65_LH_BFX2 U9225 ( .A(n32324), .Z(n32323) );
  HS65_LH_BFX2 U9226 ( .A(n32325), .Z(n32324) );
  HS65_LH_BFX2 U9227 ( .A(n32326), .Z(n32325) );
  HS65_LH_BFX2 U9228 ( .A(n32327), .Z(n32326) );
  HS65_LH_BFX2 U9229 ( .A(n32328), .Z(n32327) );
  HS65_LH_BFX2 U9230 ( .A(n32329), .Z(n32328) );
  HS65_LH_BFX2 U9231 ( .A(n32330), .Z(n32329) );
  HS65_LH_BFX2 U9232 ( .A(n32331), .Z(n32330) );
  HS65_LH_BFX2 U9233 ( .A(n32332), .Z(n32331) );
  HS65_LH_BFX2 U9234 ( .A(n32333), .Z(n32332) );
  HS65_LH_BFX2 U9235 ( .A(n32334), .Z(n32333) );
  HS65_LH_BFX2 U9236 ( .A(n32335), .Z(n32334) );
  HS65_LH_BFX2 U9237 ( .A(n32336), .Z(n32335) );
  HS65_LH_BFX2 U9238 ( .A(n32338), .Z(n32336) );
  HS65_LH_BFX2 U9250 ( .A(n15211), .Z(n32337) );
  HS65_LH_BFX2 U9252 ( .A(n32339), .Z(n32338) );
  HS65_LH_BFX2 U9253 ( .A(n32340), .Z(n32339) );
  HS65_LH_BFX2 U9255 ( .A(n38578), .Z(n32340) );
  HS65_LH_BFX2 U9256 ( .A(n33012), .Z(n32341) );
  HS65_LH_BFX2 U9258 ( .A(n32345), .Z(n32342) );
  HS65_LH_BFX2 U9259 ( .A(n32347), .Z(n32343) );
  HS65_LH_IVX2 U9261 ( .A(n32355), .Z(n32344) );
  HS65_LH_IVX2 U9262 ( .A(n32344), .Z(n32345) );
  HS65_LH_IVX2 U9264 ( .A(n32357), .Z(n32346) );
  HS65_LH_IVX2 U9265 ( .A(n32346), .Z(n32347) );
  HS65_LH_BFX2 U9267 ( .A(n32351), .Z(n32348) );
  HS65_LH_BFX2 U9268 ( .A(n32359), .Z(n32349) );
  HS65_LH_IVX2 U9270 ( .A(n32361), .Z(n32350) );
  HS65_LH_IVX2 U9271 ( .A(n32350), .Z(n32351) );
  HS65_LH_BFX2 U9273 ( .A(n17758), .Z(n32352) );
  HS65_LH_BFX2 U9274 ( .A(n17606), .Z(n32353) );
  HS65_LH_IVX2 U9276 ( .A(n32364), .Z(n32354) );
  HS65_LH_IVX2 U9277 ( .A(n32354), .Z(n32355) );
  HS65_LH_IVX2 U9279 ( .A(n32366), .Z(n32356) );
  HS65_LH_IVX2 U9280 ( .A(n32356), .Z(n32357) );
  HS65_LH_IVX2 U9282 ( .A(n32368), .Z(n32358) );
  HS65_LH_IVX2 U9283 ( .A(n32358), .Z(n32359) );
  HS65_LH_IVX2 U9285 ( .A(n32370), .Z(n32360) );
  HS65_LH_IVX2 U9286 ( .A(n32360), .Z(n32361) );
  HS65_LH_BFX2 U9288 ( .A(n32352), .Z(n32362) );
  HS65_LH_IVX2 U9289 ( .A(n32379), .Z(n32363) );
  HS65_LH_IVX2 U9291 ( .A(n32363), .Z(n32364) );
  HS65_LH_IVX2 U9292 ( .A(n32373), .Z(n32365) );
  HS65_LH_IVX2 U9294 ( .A(n32365), .Z(n32366) );
  HS65_LH_IVX2 U9295 ( .A(n32375), .Z(n32367) );
  HS65_LH_IVX2 U9297 ( .A(n32367), .Z(n32368) );
  HS65_LH_IVX2 U9298 ( .A(n32377), .Z(n32369) );
  HS65_LH_IVX2 U9300 ( .A(n32369), .Z(n32370) );
  HS65_LH_BFX2 U9302 ( .A(n32362), .Z(n32371) );
  HS65_LH_IVX2 U9304 ( .A(n32383), .Z(n32372) );
  HS65_LH_IVX2 U9306 ( .A(n32372), .Z(n32373) );
  HS65_LH_IVX2 U9356 ( .A(n32385), .Z(n32374) );
  HS65_LH_IVX2 U9357 ( .A(n32374), .Z(n32375) );
  HS65_LH_IVX2 U9359 ( .A(n32389), .Z(n32376) );
  HS65_LH_IVX2 U9360 ( .A(n32376), .Z(n32377) );
  HS65_LH_BFX2 U9362 ( .A(n32371), .Z(n32378) );
  HS65_LH_BFX2 U9363 ( .A(n32381), .Z(n32379) );
  HS65_LH_IVX2 U9365 ( .A(n32388), .Z(n32380) );
  HS65_LH_IVX2 U9366 ( .A(n32380), .Z(n32381) );
  HS65_LH_IVX2 U9368 ( .A(n32393), .Z(n32382) );
  HS65_LH_IVX2 U9369 ( .A(n32382), .Z(n32383) );
  HS65_LH_IVX2 U9371 ( .A(n32391), .Z(n32384) );
  HS65_LH_IVX2 U9372 ( .A(n32384), .Z(n32385) );
  HS65_LH_BFX2 U9374 ( .A(n32378), .Z(n32386) );
  HS65_LH_IVX2 U9375 ( .A(n32398), .Z(n32387) );
  HS65_LH_IVX2 U9377 ( .A(n32387), .Z(n32388) );
  HS65_LH_BFX2 U9378 ( .A(n32394), .Z(n32389) );
  HS65_LH_IVX2 U9380 ( .A(n32400), .Z(n32390) );
  HS65_LH_IVX2 U9381 ( .A(n32390), .Z(n32391) );
  HS65_LH_BFX2 U9383 ( .A(n32386), .Z(n32392) );
  HS65_LH_BFX2 U9384 ( .A(n32396), .Z(n32393) );
  HS65_LH_BFX2 U9386 ( .A(n32402), .Z(n32394) );
  HS65_LH_IVX2 U9387 ( .A(n32404), .Z(n32395) );
  HS65_LH_IVX2 U9389 ( .A(n32395), .Z(n32396) );
  HS65_LH_IVX2 U9390 ( .A(n32406), .Z(n32397) );
  HS65_LH_IVX2 U9392 ( .A(n32397), .Z(n32398) );
  HS65_LH_IVX2 U9393 ( .A(n32408), .Z(n32399) );
  HS65_LH_IVX2 U9395 ( .A(n32399), .Z(n32400) );
  HS65_LH_BFX2 U9396 ( .A(n32392), .Z(n32401) );
  HS65_LH_BFX2 U9398 ( .A(n32410), .Z(n32402) );
  HS65_LH_IVX2 U9399 ( .A(n32412), .Z(n32403) );
  HS65_LH_IVX2 U9401 ( .A(n32403), .Z(n32404) );
  HS65_LH_IVX2 U9402 ( .A(n32414), .Z(n32405) );
  HS65_LH_IVX2 U9404 ( .A(n32405), .Z(n32406) );
  HS65_LH_IVX2 U9405 ( .A(n32416), .Z(n32407) );
  HS65_LH_IVX2 U9407 ( .A(n32407), .Z(n32408) );
  HS65_LH_BFX2 U9408 ( .A(n32401), .Z(n32409) );
  HS65_LH_BFX2 U9410 ( .A(n32418), .Z(n32410) );
  HS65_LH_IVX2 U9439 ( .A(n32420), .Z(n32411) );
  HS65_LH_IVX2 U9440 ( .A(n32411), .Z(n32412) );
  HS65_LH_IVX2 U9464 ( .A(n32422), .Z(n32413) );
  HS65_LH_IVX2 U9466 ( .A(n32413), .Z(n32414) );
  HS65_LH_IVX2 U9467 ( .A(n32424), .Z(n32415) );
  HS65_LH_IVX2 U9469 ( .A(n32415), .Z(n32416) );
  HS65_LH_BFX2 U9470 ( .A(n32409), .Z(n32417) );
  HS65_LH_BFX2 U9472 ( .A(n32426), .Z(n32418) );
  HS65_LH_IVX2 U9473 ( .A(n32428), .Z(n32419) );
  HS65_LH_IVX2 U9475 ( .A(n32419), .Z(n32420) );
  HS65_LH_IVX2 U9476 ( .A(n32433), .Z(n32421) );
  HS65_LH_IVX2 U9478 ( .A(n32421), .Z(n32422) );
  HS65_LH_IVX2 U9479 ( .A(n32999), .Z(n32423) );
  HS65_LH_IVX2 U9481 ( .A(n32423), .Z(n32424) );
  HS65_LH_BFX2 U9482 ( .A(n32417), .Z(n32425) );
  HS65_LH_BFX2 U9484 ( .A(n32997), .Z(n32426) );
  HS65_LH_IVX2 U9485 ( .A(n33001), .Z(n32427) );
  HS65_LH_IVX2 U9487 ( .A(n32427), .Z(n32428) );
  HS65_LH_IVX2 U9488 ( .A(n17336), .Z(n32429) );
  HS65_LH_IVX2 U9490 ( .A(n32429), .Z(n32430) );
  HS65_LH_BFX2 U9491 ( .A(n32425), .Z(n32431) );
  HS65_LH_IVX2 U9493 ( .A(n32434), .Z(n32432) );
  HS65_LH_IVX2 U9494 ( .A(n32432), .Z(n32433) );
  HS65_LH_BFX2 U9496 ( .A(n32435), .Z(n32434) );
  HS65_LH_BFX2 U9497 ( .A(n32436), .Z(n32435) );
  HS65_LH_BFX2 U9500 ( .A(n32437), .Z(n32436) );
  HS65_LH_BFX2 U9502 ( .A(n32438), .Z(n32437) );
  HS65_LH_BFX2 U9503 ( .A(n32439), .Z(n32438) );
  HS65_LH_BFX2 U9505 ( .A(n32440), .Z(n32439) );
  HS65_LH_BFX2 U9506 ( .A(n14514), .Z(n32440) );
  HS65_LH_BFX2 U9508 ( .A(n32448), .Z(n32441) );
  HS65_LH_IVX2 U9509 ( .A(n32450), .Z(n32442) );
  HS65_LH_IVX2 U9511 ( .A(n32442), .Z(n32443) );
  HS65_LH_BFX2 U9512 ( .A(n32451), .Z(n32444) );
  HS65_LH_BFX2 U9514 ( .A(n15183), .Z(n32445) );
  HS65_LH_BFX2 U9516 ( .A(n2726), .Z(n32446) );
  HS65_LH_IVX2 U9518 ( .A(n32453), .Z(n32447) );
  HS65_LH_IVX2 U9520 ( .A(n32447), .Z(n32448) );
  HS65_LH_IVX2 U9522 ( .A(n34397), .Z(n32449) );
  HS65_LH_IVX2 U9527 ( .A(n32449), .Z(n32450) );
  HS65_LH_BFX2 U9528 ( .A(n32452), .Z(n32451) );
  HS65_LH_BFX2 U9529 ( .A(n32454), .Z(n32452) );
  HS65_LH_BFX2 U9530 ( .A(n32455), .Z(n32453) );
  HS65_LH_BFX2 U9531 ( .A(n32456), .Z(n32454) );
  HS65_LH_BFX2 U9532 ( .A(n32457), .Z(n32455) );
  HS65_LH_BFX2 U9533 ( .A(n32458), .Z(n32456) );
  HS65_LH_BFX2 U9534 ( .A(n32459), .Z(n32457) );
  HS65_LH_BFX2 U9535 ( .A(n32460), .Z(n32458) );
  HS65_LH_BFX2 U9536 ( .A(n32461), .Z(n32459) );
  HS65_LH_BFX2 U9537 ( .A(n32462), .Z(n32460) );
  HS65_LH_BFX2 U9538 ( .A(n32463), .Z(n32461) );
  HS65_LH_BFX2 U9539 ( .A(n32464), .Z(n32462) );
  HS65_LH_BFX2 U9540 ( .A(n32465), .Z(n32463) );
  HS65_LH_BFX2 U9541 ( .A(n32466), .Z(n32464) );
  HS65_LH_BFX2 U9542 ( .A(n32467), .Z(n32465) );
  HS65_LH_BFX2 U9543 ( .A(n32468), .Z(n32466) );
  HS65_LH_BFX2 U9544 ( .A(n32446), .Z(n32467) );
  HS65_LH_BFX2 U9545 ( .A(n2727), .Z(n32468) );
  HS65_LH_BFX2 U9546 ( .A(n32470), .Z(n32469) );
  HS65_LH_BFX2 U9547 ( .A(n32471), .Z(n32470) );
  HS65_LH_BFX2 U9548 ( .A(n32472), .Z(n32471) );
  HS65_LH_BFX2 U9549 ( .A(n32473), .Z(n32472) );
  HS65_LH_BFX2 U9550 ( .A(n32474), .Z(n32473) );
  HS65_LH_BFX2 U9551 ( .A(n32475), .Z(n32474) );
  HS65_LH_BFX2 U9552 ( .A(n32476), .Z(n32475) );
  HS65_LH_BFX2 U9553 ( .A(n32477), .Z(n32476) );
  HS65_LH_BFX2 U9554 ( .A(n32478), .Z(n32477) );
  HS65_LH_BFX2 U9555 ( .A(n32479), .Z(n32478) );
  HS65_LH_BFX2 U9557 ( .A(n32480), .Z(n32479) );
  HS65_LH_BFX2 U9559 ( .A(n32481), .Z(n32480) );
  HS65_LH_BFX2 U9561 ( .A(n32482), .Z(n32481) );
  HS65_LH_BFX2 U9563 ( .A(n32483), .Z(n32482) );
  HS65_LH_BFX2 U9565 ( .A(n32484), .Z(n32483) );
  HS65_LH_BFX2 U9567 ( .A(n32485), .Z(n32484) );
  HS65_LH_BFX2 U9569 ( .A(n32486), .Z(n32485) );
  HS65_LH_BFX2 U9571 ( .A(n15570), .Z(n32486) );
  HS65_LH_BFX2 U9573 ( .A(n32488), .Z(n32487) );
  HS65_LH_BFX2 U9575 ( .A(n32489), .Z(n32488) );
  HS65_LH_BFX2 U9577 ( .A(n32490), .Z(n32489) );
  HS65_LH_BFX2 U9579 ( .A(n32491), .Z(n32490) );
  HS65_LH_BFX2 U9581 ( .A(n32492), .Z(n32491) );
  HS65_LH_BFX2 U9583 ( .A(n32493), .Z(n32492) );
  HS65_LH_BFX2 U9585 ( .A(n32494), .Z(n32493) );
  HS65_LH_BFX2 U9587 ( .A(n32495), .Z(n32494) );
  HS65_LH_BFX2 U9639 ( .A(n32496), .Z(n32495) );
  HS65_LH_BFX2 U9641 ( .A(n32497), .Z(n32496) );
  HS65_LH_BFX2 U9643 ( .A(n32498), .Z(n32497) );
  HS65_LH_BFX2 U9645 ( .A(n32499), .Z(n32498) );
  HS65_LH_BFX2 U9647 ( .A(n32500), .Z(n32499) );
  HS65_LH_BFX2 U9649 ( .A(n32501), .Z(n32500) );
  HS65_LH_BFX2 U9651 ( .A(n32502), .Z(n32501) );
  HS65_LH_BFX2 U9653 ( .A(n32503), .Z(n32502) );
  HS65_LH_BFX2 U9656 ( .A(n15569), .Z(n32503) );
  HS65_LH_BFX2 U9657 ( .A(n17257), .Z(n32504) );
  HS65_LH_BFX2 U9661 ( .A(n32508), .Z(n32505) );
  HS65_LH_BFX2 U9663 ( .A(n15542), .Z(n32506) );
  HS65_LH_IVX2 U9665 ( .A(n32513), .Z(n32507) );
  HS65_LH_IVX2 U9667 ( .A(n32507), .Z(n32508) );
  HS65_LH_BFX2 U9669 ( .A(n17850), .Z(n32509) );
  HS65_LH_BFX2 U9671 ( .A(n32509), .Z(n32510) );
  HS65_LH_IVX2 U9673 ( .A(n32510), .Z(n32511) );
  HS65_LH_IVX2 U9698 ( .A(n32511), .Z(n32512) );
  HS65_LH_BFX2 U9699 ( .A(n17851), .Z(n32513) );
  HS65_LH_BFX2 U9700 ( .A(n40992), .Z(n32514) );
  HS65_LH_BFX2 U9701 ( .A(n32519), .Z(n32515) );
  HS65_LH_IVX2 U9702 ( .A(n32524), .Z(n32516) );
  HS65_LH_IVX2 U9703 ( .A(n32516), .Z(n32517) );
  HS65_LH_IVX2 U9704 ( .A(n32522), .Z(n32518) );
  HS65_LH_IVX2 U9705 ( .A(n32518), .Z(n32519) );
  HS65_LH_BFX2 U9725 ( .A(n17871), .Z(n32520) );
  HS65_LH_IVX2 U9727 ( .A(n32530), .Z(n32521) );
  HS65_LH_IVX2 U9729 ( .A(n32521), .Z(n32522) );
  HS65_LH_BFX2 U9730 ( .A(n32520), .Z(n32523) );
  HS65_LH_BFX2 U9732 ( .A(n32527), .Z(n32524) );
  HS65_LH_BFX2 U9733 ( .A(n15124), .Z(n32525) );
  HS65_LH_BFX2 U9735 ( .A(n32523), .Z(n32526) );
  HS65_LH_BFX2 U9737 ( .A(n32529), .Z(n32527) );
  HS65_LH_BFX2 U9738 ( .A(n32526), .Z(n32528) );
  HS65_LH_BFX2 U9740 ( .A(n32532), .Z(n32529) );
  HS65_LH_BFX2 U9741 ( .A(n32533), .Z(n32530) );
  HS65_LH_BFX2 U9743 ( .A(n32528), .Z(n32531) );
  HS65_LH_BFX2 U9744 ( .A(n32535), .Z(n32532) );
  HS65_LH_BFX2 U9746 ( .A(n32536), .Z(n32533) );
  HS65_LH_BFX2 U9747 ( .A(n32531), .Z(n32534) );
  HS65_LH_BFX2 U9749 ( .A(n32540), .Z(n32535) );
  HS65_LH_BFX2 U9750 ( .A(n32539), .Z(n32536) );
  HS65_LH_BFX2 U9752 ( .A(n32534), .Z(n32537) );
  HS65_LH_IVX2 U9753 ( .A(n32543), .Z(n32538) );
  HS65_LH_IVX2 U9755 ( .A(n32538), .Z(n32539) );
  HS65_LH_BFX2 U9756 ( .A(n32542), .Z(n32540) );
  HS65_LH_BFX2 U9758 ( .A(n32537), .Z(n32541) );
  HS65_LH_BFX2 U9759 ( .A(n32545), .Z(n32542) );
  HS65_LH_BFX2 U9761 ( .A(n32546), .Z(n32543) );
  HS65_LH_BFX2 U9762 ( .A(n32541), .Z(n32544) );
  HS65_LH_BFX2 U9764 ( .A(n32548), .Z(n32545) );
  HS65_LH_BFX2 U9765 ( .A(n32549), .Z(n32546) );
  HS65_LH_BFX2 U9767 ( .A(n32544), .Z(n32547) );
  HS65_LH_BFX2 U9768 ( .A(n32551), .Z(n32548) );
  HS65_LH_BFX2 U9770 ( .A(n32552), .Z(n32549) );
  HS65_LH_BFX2 U9771 ( .A(n32547), .Z(n32550) );
  HS65_LH_BFX2 U9773 ( .A(n32554), .Z(n32551) );
  HS65_LH_BFX2 U9774 ( .A(n32555), .Z(n32552) );
  HS65_LH_BFX2 U9776 ( .A(n32550), .Z(n32553) );
  HS65_LH_BFX2 U9777 ( .A(n32557), .Z(n32554) );
  HS65_LH_BFX2 U9779 ( .A(n32558), .Z(n32555) );
  HS65_LH_BFX2 U9781 ( .A(n32553), .Z(n32556) );
  HS65_LH_BFX2 U9783 ( .A(n32560), .Z(n32557) );
  HS65_LH_BFX2 U9813 ( .A(n32561), .Z(n32558) );
  HS65_LH_BFX2 U9815 ( .A(n32556), .Z(n32559) );
  HS65_LH_BFX2 U9818 ( .A(n32514), .Z(n32560) );
  HS65_LH_OAI112X1 U9821 ( .A(n15121), .B(n15120), .C(n15111), .D(n15119), .Z(
        n40992) );
  HS65_LH_BFX2 U9823 ( .A(n32563), .Z(n32561) );
  HS65_LH_BFX2 U9825 ( .A(n32559), .Z(n32562) );
  HS65_LH_BFX2 U9827 ( .A(n32567), .Z(n32563) );
  HS65_LH_BFX2 U9829 ( .A(n32562), .Z(n32564) );
  HS65_LH_IVX2 U9831 ( .A(n32569), .Z(n32565) );
  HS65_LH_IVX2 U9833 ( .A(n32565), .Z(n32566) );
  HS65_LH_BFX2 U9835 ( .A(n32568), .Z(n32567) );
  HS65_LH_BFX2 U9837 ( .A(n32570), .Z(n32568) );
  HS65_LH_BFX2 U9839 ( .A(n32571), .Z(n32569) );
  HS65_LH_BFX2 U9841 ( .A(n32525), .Z(n32570) );
  HS65_LH_BFX2 U9843 ( .A(n32572), .Z(n32571) );
  HS65_LH_BFX2 U9845 ( .A(n32573), .Z(n32572) );
  HS65_LH_BFX2 U9847 ( .A(n32564), .Z(n32573) );
  HS65_LH_BFX2 U9849 ( .A(n32576), .Z(n32574) );
  HS65_LH_IVX2 U9853 ( .A(n32580), .Z(n32575) );
  HS65_LH_IVX2 U9854 ( .A(n32575), .Z(n32576) );
  HS65_LH_BFX2 U9855 ( .A(n32579), .Z(n32577) );
  HS65_LH_BFX2 U9856 ( .A(n33591), .Z(n32578) );
  HS65_LH_BFX2 U9857 ( .A(n32581), .Z(n32579) );
  HS65_LH_BFX2 U9858 ( .A(n32582), .Z(n32580) );
  HS65_LH_BFX2 U9859 ( .A(n32583), .Z(n32581) );
  HS65_LH_BFX2 U9860 ( .A(n32584), .Z(n32582) );
  HS65_LH_BFX2 U9861 ( .A(n32585), .Z(n32583) );
  HS65_LH_BFX2 U9862 ( .A(n32586), .Z(n32584) );
  HS65_LH_BFX2 U9863 ( .A(n32587), .Z(n32585) );
  HS65_LH_BFX2 U9864 ( .A(n32588), .Z(n32586) );
  HS65_LH_BFX2 U9865 ( .A(n32589), .Z(n32587) );
  HS65_LH_BFX2 U9866 ( .A(n32590), .Z(n32588) );
  HS65_LH_BFX2 U9867 ( .A(n32591), .Z(n32589) );
  HS65_LH_BFX2 U9868 ( .A(n32592), .Z(n32590) );
  HS65_LH_BFX2 U9869 ( .A(n32593), .Z(n32591) );
  HS65_LH_BFX2 U9870 ( .A(n32594), .Z(n32592) );
  HS65_LH_BFX2 U9871 ( .A(n32595), .Z(n32593) );
  HS65_LH_BFX2 U9872 ( .A(n32596), .Z(n32594) );
  HS65_LH_BFX2 U9873 ( .A(n32597), .Z(n32595) );
  HS65_LH_BFX2 U9874 ( .A(n32598), .Z(n32596) );
  HS65_LH_BFX2 U9875 ( .A(n32599), .Z(n32597) );
  HS65_LH_BFX2 U9876 ( .A(n32600), .Z(n32598) );
  HS65_LH_BFX2 U9897 ( .A(n32601), .Z(n32599) );
  HS65_LH_BFX2 U9898 ( .A(n32602), .Z(n32600) );
  HS65_LH_BFX2 U9899 ( .A(n32603), .Z(n32601) );
  HS65_LH_BFX2 U9900 ( .A(n32604), .Z(n32602) );
  HS65_LH_BFX2 U9901 ( .A(n32605), .Z(n32603) );
  HS65_LH_BFX2 U9902 ( .A(n32606), .Z(n32604) );
  HS65_LH_BFX2 U9903 ( .A(n1518), .Z(n32605) );
  HS65_LH_BFX2 U9904 ( .A(n1519), .Z(n32606) );
  HS65_LH_BFX2 U9905 ( .A(n32608), .Z(n32607) );
  HS65_LH_BFX2 U9906 ( .A(n32609), .Z(n32608) );
  HS65_LH_BFX2 U9907 ( .A(n32610), .Z(n32609) );
  HS65_LH_BFX2 U9908 ( .A(n32611), .Z(n32610) );
  HS65_LH_BFX2 U9909 ( .A(n32612), .Z(n32611) );
  HS65_LH_BFX2 U9910 ( .A(n32613), .Z(n32612) );
  HS65_LH_BFX2 U9911 ( .A(n32614), .Z(n32613) );
  HS65_LH_BFX2 U9921 ( .A(n32615), .Z(n32614) );
  HS65_LH_BFX2 U9923 ( .A(n32616), .Z(n32615) );
  HS65_LH_BFX2 U9925 ( .A(n32617), .Z(n32616) );
  HS65_LH_BFX2 U9927 ( .A(n32618), .Z(n32617) );
  HS65_LH_BFX2 U9929 ( .A(n32619), .Z(n32618) );
  HS65_LH_BFX2 U9931 ( .A(n32620), .Z(n32619) );
  HS65_LH_BFX2 U9933 ( .A(n32621), .Z(n32620) );
  HS65_LH_BFX2 U9935 ( .A(n32622), .Z(n32621) );
  HS65_LH_BFX2 U9937 ( .A(n32623), .Z(n32622) );
  HS65_LH_BFX2 U9939 ( .A(n32624), .Z(n32623) );
  HS65_LH_BFX2 U9941 ( .A(n15567), .Z(n32624) );
  HS65_LH_BFX2 U9943 ( .A(n17248), .Z(n32625) );
  HS65_LH_IVX2 U9945 ( .A(n32637), .Z(n32626) );
  HS65_LH_IVX2 U9947 ( .A(n32626), .Z(n32627) );
  HS65_LH_BFX2 U9949 ( .A(n32631), .Z(n32628) );
  HS65_LH_BFX2 U9951 ( .A(n17601), .Z(n32629) );
  HS65_LH_IVX2 U9953 ( .A(n32634), .Z(n32630) );
  HS65_LH_IVX2 U9955 ( .A(n32630), .Z(n32631) );
  HS65_LH_BFX2 U9957 ( .A(n17887), .Z(n32632) );
  HS65_LH_IVX2 U9959 ( .A(n32640), .Z(n32633) );
  HS65_LH_IVX2 U9984 ( .A(n32633), .Z(n32634) );
  HS65_LH_BFX2 U9986 ( .A(n32632), .Z(n32635) );
  HS65_LH_BFX2 U9987 ( .A(n17310), .Z(n32636) );
  HS65_LH_BFX2 U9988 ( .A(n32642), .Z(n32637) );
  HS65_LH_BFX2 U9989 ( .A(n32635), .Z(n32638) );
  HS65_LH_IVX2 U9990 ( .A(n32645), .Z(n32639) );
  HS65_LH_IVX2 U9991 ( .A(n32639), .Z(n32640) );
  HS65_LH_IVX2 U9992 ( .A(n32647), .Z(n32641) );
  HS65_LH_IVX2 U9993 ( .A(n32641), .Z(n32642) );
  HS65_LH_BFX2 U9994 ( .A(n32638), .Z(n32643) );
  HS65_LH_IVX2 U9995 ( .A(n32650), .Z(n32644) );
  HS65_LH_IVX2 U9996 ( .A(n32644), .Z(n32645) );
  HS65_LH_IVX2 U9997 ( .A(n32652), .Z(n32646) );
  HS65_LH_IVX2 U9998 ( .A(n32646), .Z(n32647) );
  HS65_LH_BFX2 U9999 ( .A(n32643), .Z(n32648) );
  HS65_LH_IVX2 U10000 ( .A(n32655), .Z(n32649) );
  HS65_LH_IVX2 U10001 ( .A(n32649), .Z(n32650) );
  HS65_LH_IVX2 U10007 ( .A(n32657), .Z(n32651) );
  HS65_LH_IVX2 U10009 ( .A(n32651), .Z(n32652) );
  HS65_LH_BFX2 U10011 ( .A(n32648), .Z(n32653) );
  HS65_LH_IVX2 U10013 ( .A(n32660), .Z(n32654) );
  HS65_LH_IVX2 U10015 ( .A(n32654), .Z(n32655) );
  HS65_LH_IVX2 U10017 ( .A(n32662), .Z(n32656) );
  HS65_LH_IVX2 U10019 ( .A(n32656), .Z(n32657) );
  HS65_LH_BFX2 U10021 ( .A(n32653), .Z(n32658) );
  HS65_LH_IVX2 U10023 ( .A(n32665), .Z(n32659) );
  HS65_LH_IVX2 U10025 ( .A(n32659), .Z(n32660) );
  HS65_LH_IVX2 U10027 ( .A(n32667), .Z(n32661) );
  HS65_LH_IVX2 U10029 ( .A(n32661), .Z(n32662) );
  HS65_LH_BFX2 U10031 ( .A(n32658), .Z(n32663) );
  HS65_LH_IVX2 U10032 ( .A(n32670), .Z(n32664) );
  HS65_LH_IVX2 U10051 ( .A(n32664), .Z(n32665) );
  HS65_LH_IVX2 U10053 ( .A(n32672), .Z(n32666) );
  HS65_LH_IVX2 U10055 ( .A(n32666), .Z(n32667) );
  HS65_LH_BFX2 U10057 ( .A(n32663), .Z(n32668) );
  HS65_LH_IVX2 U10059 ( .A(n32675), .Z(n32669) );
  HS65_LH_IVX2 U10061 ( .A(n32669), .Z(n32670) );
  HS65_LH_IVX2 U10063 ( .A(n32677), .Z(n32671) );
  HS65_LH_IVX2 U10065 ( .A(n32671), .Z(n32672) );
  HS65_LH_BFX2 U10067 ( .A(n32668), .Z(n32673) );
  HS65_LH_IVX2 U10068 ( .A(n32680), .Z(n32674) );
  HS65_LH_IVX2 U10069 ( .A(n32674), .Z(n32675) );
  HS65_LH_IVX2 U10071 ( .A(n32682), .Z(n32676) );
  HS65_LH_IVX2 U10073 ( .A(n32676), .Z(n32677) );
  HS65_LH_BFX2 U10123 ( .A(n32673), .Z(n32678) );
  HS65_LH_IVX2 U10126 ( .A(n32685), .Z(n32679) );
  HS65_LH_IVX2 U10129 ( .A(n32679), .Z(n32680) );
  HS65_LH_IVX2 U10132 ( .A(n32687), .Z(n32681) );
  HS65_LH_IVX2 U10135 ( .A(n32681), .Z(n32682) );
  HS65_LH_BFX2 U10138 ( .A(n32678), .Z(n32683) );
  HS65_LH_IVX2 U10141 ( .A(n32692), .Z(n32684) );
  HS65_LH_IVX2 U10144 ( .A(n32684), .Z(n32685) );
  HS65_LH_IVX2 U10147 ( .A(n32690), .Z(n32686) );
  HS65_LH_IVX2 U10150 ( .A(n32686), .Z(n32687) );
  HS65_LH_BFX2 U10153 ( .A(n32683), .Z(n32688) );
  HS65_LH_IVX2 U10156 ( .A(n32695), .Z(n32689) );
  HS65_LH_IVX2 U10159 ( .A(n32689), .Z(n32690) );
  HS65_LH_BFX2 U10162 ( .A(n32688), .Z(n32691) );
  HS65_LH_BFX2 U10165 ( .A(n32698), .Z(n32692) );
  HS65_LH_BFX2 U10168 ( .A(n32691), .Z(n32693) );
  HS65_LH_IVX2 U10171 ( .A(n15557), .Z(n32694) );
  HS65_LH_IVX2 U10174 ( .A(n32694), .Z(n32695) );
  HS65_LH_IVX2 U10178 ( .A(n32701), .Z(n32696) );
  HS65_LH_IVX2 U10180 ( .A(n32696), .Z(n32697) );
  HS65_LH_BFX2 U10181 ( .A(n32700), .Z(n32698) );
  HS65_LH_IVX2 U10192 ( .A(n32702), .Z(n32699) );
  HS65_LH_IVX2 U10193 ( .A(n32699), .Z(n32700) );
  HS65_LH_BFX2 U10194 ( .A(n32703), .Z(n32701) );
  HS65_LH_BFX2 U10195 ( .A(n32704), .Z(n32702) );
  HS65_LH_BFX2 U10196 ( .A(n32705), .Z(n32703) );
  HS65_LH_BFX2 U10197 ( .A(n32706), .Z(n32704) );
  HS65_LH_BFX2 U10198 ( .A(n32707), .Z(n32705) );
  HS65_LH_BFX2 U10199 ( .A(n32708), .Z(n32706) );
  HS65_LH_BFX2 U10200 ( .A(n32709), .Z(n32707) );
  HS65_LH_BFX2 U10201 ( .A(n17886), .Z(n32708) );
  HS65_LH_BFX2 U10202 ( .A(n32693), .Z(n32709) );
  HS65_LH_BFX2 U10203 ( .A(n32713), .Z(n32710) );
  HS65_LH_BFX2 U10204 ( .A(n32714), .Z(n32711) );
  HS65_LH_BFX2 U10205 ( .A(n17882), .Z(n32712) );
  HS65_LH_BFX2 U10206 ( .A(n32716), .Z(n32713) );
  HS65_LH_BFX2 U10207 ( .A(n32717), .Z(n32714) );
  HS65_LH_BFX2 U10208 ( .A(n32712), .Z(n32715) );
  HS65_LH_BFX2 U10209 ( .A(n32719), .Z(n32716) );
  HS65_LH_BFX2 U10210 ( .A(n32720), .Z(n32717) );
  HS65_LH_BFX2 U10211 ( .A(n32715), .Z(n32718) );
  HS65_LH_BFX2 U10212 ( .A(n32722), .Z(n32719) );
  HS65_LH_BFX2 U10213 ( .A(n32723), .Z(n32720) );
  HS65_LH_BFX2 U10214 ( .A(n32718), .Z(n32721) );
  HS65_LH_BFX2 U10215 ( .A(n32725), .Z(n32722) );
  HS65_LH_BFX2 U10216 ( .A(n32726), .Z(n32723) );
  HS65_LH_BFX2 U10217 ( .A(n32721), .Z(n32724) );
  HS65_LH_BFX2 U10218 ( .A(n32728), .Z(n32725) );
  HS65_LH_BFX2 U10220 ( .A(n32729), .Z(n32726) );
  HS65_LH_BFX2 U10221 ( .A(n32724), .Z(n32727) );
  HS65_LH_BFX2 U10223 ( .A(n32731), .Z(n32728) );
  HS65_LH_BFX2 U10224 ( .A(n32732), .Z(n32729) );
  HS65_LH_BFX2 U10226 ( .A(n32727), .Z(n32730) );
  HS65_LH_BFX2 U10227 ( .A(n32734), .Z(n32731) );
  HS65_LH_BFX2 U10229 ( .A(n32735), .Z(n32732) );
  HS65_LH_BFX2 U10230 ( .A(n32730), .Z(n32733) );
  HS65_LH_BFX2 U10232 ( .A(n32737), .Z(n32734) );
  HS65_LH_BFX2 U10233 ( .A(n32738), .Z(n32735) );
  HS65_LH_BFX2 U10235 ( .A(n32733), .Z(n32736) );
  HS65_LH_BFX2 U10236 ( .A(n32740), .Z(n32737) );
  HS65_LH_BFX2 U10238 ( .A(n32741), .Z(n32738) );
  HS65_LH_BFX2 U10239 ( .A(n32736), .Z(n32739) );
  HS65_LH_BFX2 U10241 ( .A(n32743), .Z(n32740) );
  HS65_LH_BFX2 U10242 ( .A(n32744), .Z(n32741) );
  HS65_LH_BFX2 U10244 ( .A(n32739), .Z(n32742) );
  HS65_LH_BFX2 U10245 ( .A(n32746), .Z(n32743) );
  HS65_LH_BFX2 U10247 ( .A(n32747), .Z(n32744) );
  HS65_LH_BFX2 U10248 ( .A(n32742), .Z(n32745) );
  HS65_LH_BFX2 U10250 ( .A(n32752), .Z(n32746) );
  HS65_LH_BFX2 U10251 ( .A(n32750), .Z(n32747) );
  HS65_LH_IVX2 U10253 ( .A(n32756), .Z(n32749) );
  HS65_LH_IVX2 U10255 ( .A(n32749), .Z(n32750) );
  HS65_LH_BFX2 U10256 ( .A(n32745), .Z(n32751) );
  HS65_LH_BFX2 U10258 ( .A(n32754), .Z(n32752) );
  HS65_LH_IVX2 U10259 ( .A(n15559), .Z(n32753) );
  HS65_LH_IVX2 U10261 ( .A(n32753), .Z(n32754) );
  HS65_LH_IVX2 U10262 ( .A(n32760), .Z(n32755) );
  HS65_LH_IVX2 U10264 ( .A(n32755), .Z(n32756) );
  HS65_LH_BFX2 U10265 ( .A(n32751), .Z(n32757) );
  HS65_LH_BFX2 U10267 ( .A(n32757), .Z(n32758) );
  HS65_LH_BFX2 U10269 ( .A(n17603), .Z(n32759) );
  HS65_LH_BFX2 U10271 ( .A(n32762), .Z(n32760) );
  HS65_LH_BFX2 U10273 ( .A(n32758), .Z(n32761) );
  HS65_LH_BFX2 U10275 ( .A(n32764), .Z(n32762) );
  HS65_LH_BFX2 U10311 ( .A(n32761), .Z(n32763) );
  HS65_LH_BFX2 U10312 ( .A(n32769), .Z(n32764) );
  HS65_LH_BFX2 U10313 ( .A(n32763), .Z(n32765) );
  HS65_LH_BFX2 U10314 ( .A(n32765), .Z(n32766) );
  HS65_LH_BFX2 U10315 ( .A(n15054), .Z(n32767) );
  HS65_LH_BFX2 U10316 ( .A(n32766), .Z(n32768) );
  HS65_LH_BFX2 U10317 ( .A(n32767), .Z(n32769) );
  HS65_LH_IVX2 U10318 ( .A(n32768), .Z(n32770) );
  HS65_LH_IVX2 U10319 ( .A(n32770), .Z(n32771) );
  HS65_LH_BFX2 U10320 ( .A(n32774), .Z(n32772) );
  HS65_LH_BFX2 U10321 ( .A(n17982), .Z(n32773) );
  HS65_LH_BFX2 U10322 ( .A(n32776), .Z(n32774) );
  HS65_LH_BFX2 U10323 ( .A(n32773), .Z(n32775) );
  HS65_LH_BFX2 U10324 ( .A(n32778), .Z(n32776) );
  HS65_LH_BFX2 U10325 ( .A(n32775), .Z(n32777) );
  HS65_LH_BFX2 U10327 ( .A(n32781), .Z(n32778) );
  HS65_LH_BFX2 U10329 ( .A(n32777), .Z(n32779) );
  HS65_LH_IVX2 U10331 ( .A(n32783), .Z(n32780) );
  HS65_LH_IVX2 U10332 ( .A(n32780), .Z(n32781) );
  HS65_LH_BFX2 U10333 ( .A(n32779), .Z(n32782) );
  HS65_LH_BFX2 U10336 ( .A(n32785), .Z(n32783) );
  HS65_LH_BFX2 U10338 ( .A(n32782), .Z(n32784) );
  HS65_LH_BFX2 U10339 ( .A(n32787), .Z(n32785) );
  HS65_LH_BFX2 U10344 ( .A(n32784), .Z(n32786) );
  HS65_LH_BFX2 U10348 ( .A(n32789), .Z(n32787) );
  HS65_LH_BFX2 U10349 ( .A(n32786), .Z(n32788) );
  HS65_LH_BFX2 U10351 ( .A(n32791), .Z(n32789) );
  HS65_LH_BFX2 U10952 ( .A(n32788), .Z(n32790) );
  HS65_LH_BFX2 U10957 ( .A(n32793), .Z(n32791) );
  HS65_LH_BFX2 U10961 ( .A(n32790), .Z(n32792) );
  HS65_LH_BFX2 U10965 ( .A(n32795), .Z(n32793) );
  HS65_LH_BFX2 U10969 ( .A(n32792), .Z(n32794) );
  HS65_LH_BFX2 U10973 ( .A(n32797), .Z(n32795) );
  HS65_LH_BFX2 U10977 ( .A(n32794), .Z(n32796) );
  HS65_LH_BFX2 U10981 ( .A(n32799), .Z(n32797) );
  HS65_LH_BFX2 U10985 ( .A(n32796), .Z(n32798) );
  HS65_LH_BFX2 U10989 ( .A(n32801), .Z(n32799) );
  HS65_LH_BFX2 U10993 ( .A(n32798), .Z(n32800) );
  HS65_LH_BFX2 U10997 ( .A(n32803), .Z(n32801) );
  HS65_LH_BFX2 U11001 ( .A(n32800), .Z(n32802) );
  HS65_LH_BFX2 U11005 ( .A(n32807), .Z(n32803) );
  HS65_LH_BFX2 U11009 ( .A(n32802), .Z(n32804) );
  HS65_LH_IVX2 U11013 ( .A(n32808), .Z(n32805) );
  HS65_LH_IVX2 U11017 ( .A(n32805), .Z(n32806) );
  HS65_LH_BFX2 U11021 ( .A(n15552), .Z(n32807) );
  HS65_LH_BFX2 U11172 ( .A(n32809), .Z(n32808) );
  HS65_LH_BFX2 U11174 ( .A(n32810), .Z(n32809) );
  HS65_LH_BFX2 U11175 ( .A(n32811), .Z(n32810) );
  HS65_LH_BFX2 U11177 ( .A(n32804), .Z(n32811) );
  HS65_LH_IVX2 U11178 ( .A(n33598), .Z(n32812) );
  HS65_LH_IVX2 U11180 ( .A(n32812), .Z(n32813) );
  HS65_LH_BFX2 U11181 ( .A(n32816), .Z(n32814) );
  HS65_LH_BFX2 U11183 ( .A(n1564), .Z(n32815) );
  HS65_LH_BFX2 U11184 ( .A(n32818), .Z(n32816) );
  HS65_LH_BFX2 U11186 ( .A(n32815), .Z(n32817) );
  HS65_LH_BFX2 U11188 ( .A(n32820), .Z(n32818) );
  HS65_LH_BFX2 U11189 ( .A(n32817), .Z(n32819) );
  HS65_LH_BFX2 U11191 ( .A(n32822), .Z(n32820) );
  HS65_LH_BFX2 U11192 ( .A(n32819), .Z(n32821) );
  HS65_LH_BFX2 U11194 ( .A(n32824), .Z(n32822) );
  HS65_LH_BFX2 U11195 ( .A(n32821), .Z(n32823) );
  HS65_LH_BFX2 U11197 ( .A(n32826), .Z(n32824) );
  HS65_LH_BFX2 U11198 ( .A(n32823), .Z(n32825) );
  HS65_LH_BFX2 U11199 ( .A(n32828), .Z(n32826) );
  HS65_LH_BFX2 U11201 ( .A(n32825), .Z(n32827) );
  HS65_LH_BFX2 U11202 ( .A(n32830), .Z(n32828) );
  HS65_LH_BFX2 U11203 ( .A(n32827), .Z(n32829) );
  HS65_LH_BFX2 U11205 ( .A(n32832), .Z(n32830) );
  HS65_LH_BFX2 U11206 ( .A(n32829), .Z(n32831) );
  HS65_LH_BFX2 U11207 ( .A(n32834), .Z(n32832) );
  HS65_LH_BFX2 U11209 ( .A(n32831), .Z(n32833) );
  HS65_LH_BFX2 U11210 ( .A(n32836), .Z(n32834) );
  HS65_LH_BFX2 U11211 ( .A(n32833), .Z(n32835) );
  HS65_LH_BFX2 U11213 ( .A(n32838), .Z(n32836) );
  HS65_LH_BFX2 U11214 ( .A(n32835), .Z(n32837) );
  HS65_LH_BFX2 U11215 ( .A(n32841), .Z(n32838) );
  HS65_LH_BFX2 U11217 ( .A(n32837), .Z(n32839) );
  HS65_LH_IVX2 U11218 ( .A(n32845), .Z(n32840) );
  HS65_LH_IVX2 U11219 ( .A(n32840), .Z(n32841) );
  HS65_LH_BFX2 U11221 ( .A(n32839), .Z(n32842) );
  HS65_LH_BFX2 U11222 ( .A(n16760), .Z(n32843) );
  HS65_LH_IVX2 U11223 ( .A(n1565), .Z(n32844) );
  HS65_LH_IVX2 U11225 ( .A(n32844), .Z(n32845) );
  HS65_LH_IVX2 U11226 ( .A(n32842), .Z(n32846) );
  HS65_LH_IVX2 U11227 ( .A(n32846), .Z(n32847) );
  HS65_LH_BFX2 U11229 ( .A(n32853), .Z(n32848) );
  HS65_LH_BFX2 U11230 ( .A(n32880), .Z(n32849) );
  HS65_LH_BFX2 U11231 ( .A(n17942), .Z(n32850) );
  HS65_LH_BFX2 U11233 ( .A(n17255), .Z(n32851) );
  HS65_LH_IVX2 U11234 ( .A(n32856), .Z(n32852) );
  HS65_LH_IVX2 U11235 ( .A(n32852), .Z(n32853) );
  HS65_LH_BFX2 U11236 ( .A(n15551), .Z(n32854) );
  HS65_LH_BFX2 U11237 ( .A(n32854), .Z(n32855) );
  HS65_LH_BFX2 U11239 ( .A(n32858), .Z(n32856) );
  HS65_LH_BFX2 U11240 ( .A(n32855), .Z(n32857) );
  HS65_LH_BFX2 U11241 ( .A(n32860), .Z(n32858) );
  HS65_LH_BFX2 U11242 ( .A(n32857), .Z(n32859) );
  HS65_LH_BFX2 U11255 ( .A(n32862), .Z(n32860) );
  HS65_LH_BFX2 U11258 ( .A(n32859), .Z(n32861) );
  HS65_LH_BFX2 U11261 ( .A(n32864), .Z(n32862) );
  HS65_LH_BFX2 U11264 ( .A(n32861), .Z(n32863) );
  HS65_LH_BFX2 U11267 ( .A(n32866), .Z(n32864) );
  HS65_LH_BFX2 U11270 ( .A(n32863), .Z(n32865) );
  HS65_LH_BFX2 U11273 ( .A(n32868), .Z(n32866) );
  HS65_LH_BFX2 U11275 ( .A(n32865), .Z(n32867) );
  HS65_LH_BFX2 U11277 ( .A(n32870), .Z(n32868) );
  HS65_LH_BFX2 U11279 ( .A(n32867), .Z(n32869) );
  HS65_LH_BFX2 U11284 ( .A(n32872), .Z(n32870) );
  HS65_LH_BFX2 U11287 ( .A(n32869), .Z(n32871) );
  HS65_LH_BFX2 U11289 ( .A(n32874), .Z(n32872) );
  HS65_LH_BFX2 U11291 ( .A(n32871), .Z(n32873) );
  HS65_LH_BFX2 U11293 ( .A(n32876), .Z(n32874) );
  HS65_LH_BFX2 U11295 ( .A(n32873), .Z(n32875) );
  HS65_LH_BFX2 U11297 ( .A(n32878), .Z(n32876) );
  HS65_LH_BFX2 U11299 ( .A(n32875), .Z(n32877) );
  HS65_LH_BFX2 U11301 ( .A(n32881), .Z(n32878) );
  HS65_LH_IVX2 U11303 ( .A(n32877), .Z(n32879) );
  HS65_LH_IVX2 U11305 ( .A(n32879), .Z(n32880) );
  HS65_LH_BFX2 U11307 ( .A(n32882), .Z(n32881) );
  HS65_LH_BFX2 U11309 ( .A(n32883), .Z(n32882) );
  HS65_LH_BFX2 U11311 ( .A(n32884), .Z(n32883) );
  HS65_LH_BFX2 U11313 ( .A(n32885), .Z(n32884) );
  HS65_LH_BFX2 U11315 ( .A(n32886), .Z(n32885) );
  HS65_LH_BFX2 U11317 ( .A(n32850), .Z(n32886) );
  HS65_LH_BFX2 U11327 ( .A(n32894), .Z(n32887) );
  HS65_LH_BFX2 U11328 ( .A(n32891), .Z(n32888) );
  HS65_LH_BFX2 U11329 ( .A(n32893), .Z(n32889) );
  HS65_LH_IVX2 U11330 ( .A(n32898), .Z(n32890) );
  HS65_LH_IVX2 U11331 ( .A(n32890), .Z(n32891) );
  HS65_LH_IVX2 U11332 ( .A(n32896), .Z(n32892) );
  HS65_LH_IVX2 U11333 ( .A(n32892), .Z(n32893) );
  HS65_LH_BFX2 U11334 ( .A(n32897), .Z(n32894) );
  HS65_LH_IVX2 U11335 ( .A(n33594), .Z(n32895) );
  HS65_LH_IVX2 U11336 ( .A(n32895), .Z(n32896) );
  HS65_LH_BFX2 U11337 ( .A(n32899), .Z(n32897) );
  HS65_LH_BFX2 U11338 ( .A(n32900), .Z(n32898) );
  HS65_LH_BFX2 U11339 ( .A(n32901), .Z(n32899) );
  HS65_LH_BFX2 U11340 ( .A(n32902), .Z(n32900) );
  HS65_LH_BFX2 U11341 ( .A(n32903), .Z(n32901) );
  HS65_LH_BFX2 U11342 ( .A(n32904), .Z(n32902) );
  HS65_LH_BFX2 U11343 ( .A(n32905), .Z(n32903) );
  HS65_LH_BFX2 U11344 ( .A(n32906), .Z(n32904) );
  HS65_LH_BFX2 U11345 ( .A(n32907), .Z(n32905) );
  HS65_LH_BFX2 U11346 ( .A(n32908), .Z(n32906) );
  HS65_LH_BFX2 U11347 ( .A(n32909), .Z(n32907) );
  HS65_LH_BFX2 U11348 ( .A(n32910), .Z(n32908) );
  HS65_LH_BFX2 U11349 ( .A(n32911), .Z(n32909) );
  HS65_LH_BFX2 U11350 ( .A(n32912), .Z(n32910) );
  HS65_LH_BFX2 U11352 ( .A(n32913), .Z(n32911) );
  HS65_LH_BFX2 U11552 ( .A(n32914), .Z(n32912) );
  HS65_LH_BFX2 U11558 ( .A(n32915), .Z(n32913) );
  HS65_LH_BFX2 U11564 ( .A(n32916), .Z(n32914) );
  HS65_LH_BFX2 U11572 ( .A(n32917), .Z(n32915) );
  HS65_LH_BFX2 U11577 ( .A(n32918), .Z(n32916) );
  HS65_LH_BFX2 U11585 ( .A(n32919), .Z(n32917) );
  HS65_LH_BFX2 U11592 ( .A(n32920), .Z(n32918) );
  HS65_LH_BFX2 U11599 ( .A(n32921), .Z(n32919) );
  HS65_LH_BFX2 U11604 ( .A(n32922), .Z(n32920) );
  HS65_LH_BFX2 U11612 ( .A(n32923), .Z(n32921) );
  HS65_LH_BFX2 U11619 ( .A(n32924), .Z(n32922) );
  HS65_LH_BFX2 U11626 ( .A(n1587), .Z(n32923) );
  HS65_LH_BFX2 U11631 ( .A(n1588), .Z(n32924) );
  HS65_LH_AND2ABX9 U11639 ( .A(n14919), .B(n17474), .Z(n14930) );
  HS65_LH_BFX2 U11646 ( .A(n32927), .Z(n32925) );
  HS65_LH_BFX2 U11651 ( .A(n15548), .Z(n32926) );
  HS65_LH_BFX2 U11659 ( .A(n32929), .Z(n32927) );
  HS65_LH_BFX2 U11666 ( .A(n32926), .Z(n32928) );
  HS65_LH_BFX2 U11673 ( .A(n32931), .Z(n32929) );
  HS65_LH_BFX2 U11712 ( .A(n32932), .Z(n32930) );
  HS65_LH_BFX2 U11713 ( .A(n32933), .Z(n32931) );
  HS65_LH_BFX2 U11714 ( .A(n32934), .Z(n32932) );
  HS65_LH_BFX2 U11715 ( .A(n32935), .Z(n32933) );
  HS65_LH_BFX2 U11716 ( .A(n32936), .Z(n32934) );
  HS65_LH_BFX2 U11717 ( .A(n32937), .Z(n32935) );
  HS65_LH_BFX2 U11718 ( .A(n32938), .Z(n32936) );
  HS65_LH_BFX2 U11719 ( .A(n32939), .Z(n32937) );
  HS65_LH_BFX2 U11720 ( .A(n32940), .Z(n32938) );
  HS65_LH_BFX2 U11721 ( .A(n32941), .Z(n32939) );
  HS65_LH_BFX2 U11722 ( .A(n32942), .Z(n32940) );
  HS65_LH_BFX2 U11723 ( .A(n32943), .Z(n32941) );
  HS65_LH_BFX2 U11724 ( .A(n32944), .Z(n32942) );
  HS65_LH_BFX2 U11725 ( .A(n32945), .Z(n32943) );
  HS65_LH_BFX2 U11726 ( .A(n32946), .Z(n32944) );
  HS65_LH_BFX2 U11727 ( .A(n32947), .Z(n32945) );
  HS65_LH_BFX2 U11728 ( .A(n32948), .Z(n32946) );
  HS65_LH_BFX2 U11729 ( .A(n32949), .Z(n32947) );
  HS65_LH_BFX2 U11730 ( .A(n32950), .Z(n32948) );
  HS65_LH_BFX2 U11731 ( .A(n32951), .Z(n32949) );
  HS65_LH_BFX2 U11732 ( .A(n32952), .Z(n32950) );
  HS65_LH_BFX2 U11733 ( .A(n32953), .Z(n32951) );
  HS65_LH_BFX2 U11734 ( .A(n32954), .Z(n32952) );
  HS65_LH_BFX2 U11735 ( .A(n32955), .Z(n32953) );
  HS65_LH_BFX2 U11736 ( .A(n32956), .Z(n32954) );
  HS65_LH_BFX2 U11737 ( .A(n32957), .Z(n32955) );
  HS65_LH_BFX2 U11738 ( .A(n32928), .Z(n32956) );
  HS65_LH_BFX2 U11739 ( .A(n32958), .Z(n32957) );
  HS65_LH_BFX2 U11740 ( .A(n32959), .Z(n32958) );
  HS65_LH_BFX2 U11741 ( .A(n32960), .Z(n32959) );
  HS65_LH_BFX2 U11742 ( .A(n32961), .Z(n32960) );
  HS65_LH_BFX2 U11743 ( .A(n17948), .Z(n32961) );
  HS65_LH_BFX2 U11744 ( .A(n32969), .Z(n32962) );
  HS65_LH_BFX2 U11745 ( .A(n32970), .Z(n32963) );
  HS65_LH_BFX2 U11746 ( .A(n32966), .Z(n32964) );
  HS65_LH_IVX2 U11747 ( .A(n33596), .Z(n32965) );
  HS65_LH_IVX2 U11748 ( .A(n32965), .Z(n32966) );
  HS65_LH_BFX2 U11749 ( .A(n1611), .Z(n32967) );
  HS65_LH_IVX2 U11750 ( .A(n32972), .Z(n32968) );
  HS65_LH_IVX2 U11751 ( .A(n32968), .Z(n32969) );
  HS65_LH_BFX2 U11752 ( .A(n32971), .Z(n32970) );
  HS65_LH_BFX2 U11753 ( .A(n32973), .Z(n32971) );
  HS65_LH_BFX2 U11754 ( .A(n32974), .Z(n32972) );
  HS65_LH_BFX2 U11755 ( .A(n32975), .Z(n32973) );
  HS65_LH_BFX2 U11756 ( .A(n32976), .Z(n32974) );
  HS65_LH_BFX2 U11757 ( .A(n32977), .Z(n32975) );
  HS65_LH_BFX2 U11758 ( .A(n32978), .Z(n32976) );
  HS65_LH_BFX2 U11759 ( .A(n32979), .Z(n32977) );
  HS65_LH_BFX2 U11760 ( .A(n32980), .Z(n32978) );
  HS65_LH_BFX2 U11761 ( .A(n32981), .Z(n32979) );
  HS65_LH_BFX2 U11762 ( .A(n32982), .Z(n32980) );
  HS65_LH_BFX2 U11763 ( .A(n32983), .Z(n32981) );
  HS65_LH_BFX2 U11764 ( .A(n32984), .Z(n32982) );
  HS65_LH_BFX2 U11765 ( .A(n32985), .Z(n32983) );
  HS65_LH_BFX2 U11766 ( .A(n32986), .Z(n32984) );
  HS65_LH_BFX2 U11767 ( .A(n32987), .Z(n32985) );
  HS65_LH_BFX2 U11768 ( .A(n32988), .Z(n32986) );
  HS65_LH_BFX2 U11769 ( .A(n32989), .Z(n32987) );
  HS65_LH_BFX2 U11770 ( .A(n32990), .Z(n32988) );
  HS65_LH_BFX2 U11771 ( .A(n32991), .Z(n32989) );
  HS65_LH_BFX2 U11772 ( .A(n32992), .Z(n32990) );
  HS65_LH_BFX2 U11773 ( .A(n32993), .Z(n32991) );
  HS65_LH_BFX2 U11774 ( .A(n32994), .Z(n32992) );
  HS65_LH_BFX2 U11775 ( .A(n32995), .Z(n32993) );
  HS65_LH_BFX2 U11776 ( .A(n32996), .Z(n32994) );
  HS65_LH_BFX2 U11777 ( .A(n1610), .Z(n32995) );
  HS65_LH_BFX2 U11778 ( .A(n32967), .Z(n32996) );
  HS65_LH_BFX2 U11779 ( .A(n33000), .Z(n32997) );
  HS65_LH_BFX2 U11780 ( .A(n32431), .Z(n32998) );
  HS65_LH_BFX2 U11781 ( .A(n15536), .Z(n32999) );
  HS65_LH_BFX2 U11782 ( .A(n33003), .Z(n33000) );
  HS65_LH_BFX2 U11783 ( .A(n33004), .Z(n33001) );
  HS65_LH_BFX2 U11784 ( .A(n32998), .Z(n33002) );
  HS65_LH_BFX2 U11785 ( .A(n33006), .Z(n33003) );
  HS65_LH_BFX2 U11786 ( .A(n33007), .Z(n33004) );
  HS65_LH_BFX2 U11787 ( .A(n33002), .Z(n33005) );
  HS65_LH_BFX2 U11788 ( .A(n17757), .Z(n33006) );
  HS65_LH_BFX2 U11789 ( .A(n33010), .Z(n33007) );
  HS65_LH_BFX2 U11790 ( .A(n33005), .Z(n33008) );
  HS65_LH_IVX2 U11791 ( .A(n17756), .Z(n33009) );
  HS65_LH_IVX2 U11792 ( .A(n33009), .Z(n33010) );
  HS65_LH_IVX2 U11793 ( .A(n33008), .Z(n33011) );
  HS65_LH_IVX2 U11794 ( .A(n33011), .Z(n33012) );
  HS65_LH_BFX2 U11795 ( .A(n33016), .Z(n33013) );
  HS65_LH_BFX2 U11796 ( .A(n15554), .Z(n33014) );
  HS65_LH_IVX2 U11797 ( .A(n33019), .Z(n33015) );
  HS65_LH_IVX2 U11798 ( .A(n33015), .Z(n33016) );
  HS65_LH_BFX2 U11799 ( .A(n33014), .Z(n33017) );
  HS65_LH_IVX2 U11800 ( .A(n33022), .Z(n33018) );
  HS65_LH_IVX2 U11801 ( .A(n33018), .Z(n33019) );
  HS65_LH_BFX2 U11802 ( .A(n33021), .Z(n33020) );
  HS65_LH_BFX2 U11803 ( .A(n33023), .Z(n33021) );
  HS65_LH_BFX2 U11804 ( .A(n33024), .Z(n33022) );
  HS65_LH_BFX2 U11805 ( .A(n33025), .Z(n33023) );
  HS65_LH_BFX2 U11806 ( .A(n33026), .Z(n33024) );
  HS65_LH_BFX2 U11807 ( .A(n33027), .Z(n33025) );
  HS65_LH_BFX2 U11808 ( .A(n33028), .Z(n33026) );
  HS65_LH_BFX2 U11809 ( .A(n33029), .Z(n33027) );
  HS65_LH_BFX2 U11810 ( .A(n33030), .Z(n33028) );
  HS65_LH_BFX2 U11811 ( .A(n33031), .Z(n33029) );
  HS65_LH_BFX2 U11812 ( .A(n33032), .Z(n33030) );
  HS65_LH_BFX2 U11813 ( .A(n33033), .Z(n33031) );
  HS65_LH_BFX2 U11814 ( .A(n33034), .Z(n33032) );
  HS65_LH_BFX2 U11815 ( .A(n33035), .Z(n33033) );
  HS65_LH_BFX2 U11816 ( .A(n33036), .Z(n33034) );
  HS65_LH_BFX2 U11817 ( .A(n33037), .Z(n33035) );
  HS65_LH_BFX2 U11818 ( .A(n33038), .Z(n33036) );
  HS65_LH_BFX2 U11819 ( .A(n33039), .Z(n33037) );
  HS65_LH_BFX2 U11820 ( .A(n33040), .Z(n33038) );
  HS65_LH_BFX2 U11821 ( .A(n33041), .Z(n33039) );
  HS65_LH_BFX2 U11822 ( .A(n33042), .Z(n33040) );
  HS65_LH_BFX2 U11823 ( .A(n33043), .Z(n33041) );
  HS65_LH_BFX2 U11824 ( .A(n33044), .Z(n33042) );
  HS65_LH_BFX2 U11825 ( .A(n33017), .Z(n33043) );
  HS65_LH_BFX2 U11826 ( .A(n33046), .Z(n33044) );
  HS65_LH_BFX2 U11827 ( .A(n17246), .Z(n33045) );
  HS65_LH_BFX2 U11828 ( .A(n33047), .Z(n33046) );
  HS65_LH_BFX2 U11829 ( .A(n33048), .Z(n33047) );
  HS65_LH_BFX2 U11830 ( .A(n33049), .Z(n33048) );
  HS65_LH_BFX2 U11831 ( .A(n33050), .Z(n33049) );
  HS65_LH_BFX2 U11832 ( .A(n33051), .Z(n33050) );
  HS65_LH_BFX2 U11833 ( .A(n17979), .Z(n33051) );
  HS65_LH_BFX2 U11834 ( .A(n33053), .Z(n33052) );
  HS65_LH_BFX2 U11835 ( .A(n33054), .Z(n33053) );
  HS65_LH_BFX2 U11836 ( .A(n33055), .Z(n33054) );
  HS65_LH_BFX2 U11837 ( .A(n33056), .Z(n33055) );
  HS65_LH_BFX2 U11838 ( .A(n33057), .Z(n33056) );
  HS65_LH_BFX2 U11839 ( .A(n33058), .Z(n33057) );
  HS65_LH_BFX2 U11840 ( .A(n33059), .Z(n33058) );
  HS65_LH_BFX2 U11841 ( .A(n33060), .Z(n33059) );
  HS65_LH_BFX2 U11842 ( .A(n33061), .Z(n33060) );
  HS65_LH_BFX2 U11843 ( .A(n33062), .Z(n33061) );
  HS65_LH_BFX2 U11844 ( .A(n33063), .Z(n33062) );
  HS65_LH_BFX2 U11845 ( .A(n33064), .Z(n33063) );
  HS65_LH_BFX2 U11846 ( .A(n33065), .Z(n33064) );
  HS65_LH_BFX2 U11847 ( .A(n33066), .Z(n33065) );
  HS65_LH_BFX2 U11848 ( .A(n15426), .Z(n33066) );
  HS65_LH_BFX2 U11849 ( .A(n33068), .Z(n33067) );
  HS65_LH_BFX2 U11850 ( .A(n33640), .Z(n33068) );
  HS65_LH_BFX2 U11851 ( .A(n17602), .Z(n33069) );
  HS65_LH_BFX2 U11852 ( .A(n33069), .Z(n33070) );
  HS65_LH_BFX2 U11853 ( .A(n33076), .Z(n33071) );
  HS65_LH_IVX2 U11854 ( .A(n33106), .Z(n33072) );
  HS65_LH_IVX2 U11855 ( .A(n33072), .Z(n33073) );
  HS65_LH_BFX2 U11856 ( .A(n33078), .Z(n33074) );
  HS65_LH_IVX2 U11857 ( .A(n33092), .Z(n33075) );
  HS65_LH_IVX2 U11858 ( .A(n33075), .Z(n33076) );
  HS65_LH_IVX2 U11859 ( .A(n33094), .Z(n33077) );
  HS65_LH_IVX2 U11860 ( .A(n33077), .Z(n33078) );
  HS65_LH_BFX2 U11861 ( .A(n33095), .Z(n33079) );
  HS65_LH_BFX2 U11862 ( .A(n33084), .Z(n33080) );
  HS65_LH_BFX2 U11863 ( .A(n33086), .Z(n33081) );
  HS65_LH_BFX2 U11864 ( .A(n33089), .Z(n33082) );
  HS65_LH_IVX2 U11865 ( .A(n33098), .Z(n33083) );
  HS65_LH_IVX2 U11866 ( .A(n33083), .Z(n33084) );
  HS65_LH_IVX2 U11867 ( .A(n33101), .Z(n33085) );
  HS65_LH_IVX2 U11868 ( .A(n33085), .Z(n33086) );
  HS65_LH_BFX2 U11869 ( .A(n33103), .Z(n33087) );
  HS65_LH_IVX2 U11870 ( .A(n33105), .Z(n33088) );
  HS65_LH_IVX2 U11871 ( .A(n33088), .Z(n33089) );
  HS65_LH_BFX2 U11872 ( .A(n33099), .Z(n33090) );
  HS65_LH_IVX2 U11873 ( .A(n33108), .Z(n33091) );
  HS65_LH_IVX2 U11874 ( .A(n33091), .Z(n33092) );
  HS65_LH_IVX2 U11875 ( .A(n33112), .Z(n33093) );
  HS65_LH_IVX2 U11876 ( .A(n33093), .Z(n33094) );
  HS65_LH_BFX2 U11877 ( .A(n33109), .Z(n33095) );
  HS65_LH_BFX2 U11878 ( .A(n17824), .Z(n33096) );
  HS65_LH_IVX2 U11879 ( .A(n33114), .Z(n33097) );
  HS65_LH_IVX2 U11880 ( .A(n33097), .Z(n33098) );
  HS65_LH_BFX2 U11881 ( .A(n33110), .Z(n33099) );
  HS65_LH_IVX2 U11882 ( .A(n17825), .Z(n33100) );
  HS65_LH_IVX2 U11883 ( .A(n33100), .Z(n33101) );
  HS65_LH_IVX2 U11884 ( .A(n33115), .Z(n33102) );
  HS65_LH_IVX2 U11885 ( .A(n33102), .Z(n33103) );
  HS65_LH_IVX2 U11886 ( .A(n33117), .Z(n33104) );
  HS65_LH_IVX2 U11887 ( .A(n33104), .Z(n33105) );
  HS65_LH_BFX2 U11888 ( .A(n33111), .Z(n33106) );
  HS65_LH_IVX2 U11889 ( .A(n33120), .Z(n33107) );
  HS65_LH_IVX2 U11890 ( .A(n33107), .Z(n33108) );
  HS65_LH_BFX2 U11891 ( .A(n33113), .Z(n33109) );
  HS65_LH_BFX2 U11892 ( .A(n33116), .Z(n33110) );
  HS65_LH_BFX2 U11893 ( .A(n33118), .Z(n33111) );
  HS65_LH_BFX2 U11894 ( .A(n33119), .Z(n33112) );
  HS65_LH_BFX2 U11895 ( .A(n33121), .Z(n33113) );
  HS65_LH_BFX2 U11896 ( .A(n33122), .Z(n33114) );
  HS65_LH_BFX2 U11897 ( .A(n34013), .Z(n33115) );
  HS65_LH_BFX2 U11898 ( .A(n33123), .Z(n33116) );
  HS65_LH_BFX2 U11899 ( .A(n33124), .Z(n33117) );
  HS65_LH_BFX2 U11900 ( .A(n33125), .Z(n33118) );
  HS65_LH_BFX2 U11901 ( .A(n33126), .Z(n33119) );
  HS65_LH_BFX2 U11902 ( .A(n33127), .Z(n33120) );
  HS65_LH_BFX2 U11903 ( .A(n33128), .Z(n33121) );
  HS65_LH_BFX2 U11904 ( .A(n33129), .Z(n33122) );
  HS65_LH_BFX2 U11905 ( .A(n33130), .Z(n33123) );
  HS65_LH_BFX2 U11906 ( .A(n33131), .Z(n33124) );
  HS65_LH_BFX2 U11907 ( .A(n33132), .Z(n33125) );
  HS65_LH_BFX2 U11908 ( .A(n33133), .Z(n33126) );
  HS65_LH_BFX2 U11909 ( .A(n33134), .Z(n33127) );
  HS65_LH_BFX2 U11910 ( .A(n33647), .Z(n33128) );
  HS65_LH_BFX2 U11911 ( .A(n33135), .Z(n33129) );
  HS65_LH_BFX2 U11912 ( .A(n33136), .Z(n33130) );
  HS65_LH_BFX2 U11913 ( .A(n33137), .Z(n33131) );
  HS65_LH_BFX2 U11914 ( .A(n33138), .Z(n33132) );
  HS65_LH_BFX2 U11915 ( .A(n33139), .Z(n33133) );
  HS65_LH_BFX2 U11916 ( .A(n33140), .Z(n33134) );
  HS65_LH_BFX2 U11917 ( .A(n33141), .Z(n33135) );
  HS65_LH_BFX2 U11918 ( .A(n33142), .Z(n33136) );
  HS65_LH_BFX2 U11919 ( .A(n33143), .Z(n33137) );
  HS65_LH_BFX2 U11920 ( .A(n33648), .Z(n33138) );
  HS65_LH_BFX2 U11921 ( .A(n33144), .Z(n33139) );
  HS65_LH_BFX2 U11922 ( .A(n33145), .Z(n33140) );
  HS65_LH_BFX2 U11923 ( .A(n33146), .Z(n33141) );
  HS65_LH_BFX2 U11924 ( .A(n33147), .Z(n33142) );
  HS65_LH_BFX2 U11925 ( .A(n33148), .Z(n33143) );
  HS65_LH_BFX2 U11926 ( .A(n33149), .Z(n33144) );
  HS65_LH_BFX2 U11927 ( .A(n33150), .Z(n33145) );
  HS65_LH_BFX2 U11928 ( .A(n33151), .Z(n33146) );
  HS65_LH_BFX2 U11929 ( .A(n33152), .Z(n33147) );
  HS65_LH_BFX2 U11930 ( .A(n33153), .Z(n33148) );
  HS65_LH_BFX2 U11932 ( .A(n33154), .Z(n33149) );
  HS65_LH_BFX2 U11933 ( .A(n33510), .Z(n33150) );
  HS65_LH_BFX2 U11934 ( .A(n33155), .Z(n33151) );
  HS65_LH_BFX2 U11935 ( .A(n33156), .Z(n33152) );
  HS65_LH_BFX2 U11936 ( .A(n33157), .Z(n33153) );
  HS65_LH_BFX2 U11937 ( .A(n33158), .Z(n33154) );
  HS65_LH_BFX2 U11938 ( .A(n33159), .Z(n33155) );
  HS65_LH_BFX2 U11939 ( .A(n33160), .Z(n33156) );
  HS65_LH_BFX2 U11940 ( .A(n33161), .Z(n33157) );
  HS65_LH_BFX2 U11941 ( .A(n33162), .Z(n33158) );
  HS65_LH_BFX2 U11942 ( .A(n33511), .Z(n33159) );
  HS65_LH_BFX2 U11944 ( .A(n33163), .Z(n33160) );
  HS65_LH_BFX2 U11945 ( .A(n33164), .Z(n33161) );
  HS65_LH_BFX2 U11946 ( .A(n33165), .Z(n33162) );
  HS65_LH_BFX2 U11947 ( .A(n33166), .Z(n33163) );
  HS65_LH_BFX2 U11948 ( .A(n33167), .Z(n33164) );
  HS65_LH_BFX2 U11949 ( .A(n33168), .Z(n33165) );
  HS65_LH_BFX2 U11950 ( .A(n33169), .Z(n33166) );
  HS65_LH_BFX2 U11951 ( .A(n33170), .Z(n33167) );
  HS65_LH_BFX2 U11952 ( .A(n17818), .Z(n33168) );
  HS65_LH_BFX2 U11953 ( .A(n33171), .Z(n33169) );
  HS65_LH_BFX2 U11954 ( .A(n33172), .Z(n33170) );
  HS65_LH_BFX2 U11955 ( .A(n33173), .Z(n33171) );
  HS65_LH_BFX2 U11956 ( .A(n33174), .Z(n33172) );
  HS65_LH_BFX2 U11957 ( .A(n33175), .Z(n33173) );
  HS65_LH_BFX2 U11958 ( .A(n17817), .Z(n33174) );
  HS65_LH_BFX2 U11959 ( .A(n33176), .Z(n33175) );
  HS65_LH_BFX2 U11960 ( .A(n17816), .Z(n33176) );
  HS65_LH_BFX2 U11961 ( .A(n33182), .Z(n33177) );
  HS65_LH_BFX2 U11962 ( .A(n1633), .Z(n33178) );
  HS65_LH_BFX2 U11963 ( .A(n33181), .Z(n33179) );
  HS65_LH_IVX2 U11964 ( .A(n33601), .Z(n33180) );
  HS65_LH_IVX2 U11965 ( .A(n33180), .Z(n33181) );
  HS65_LH_BFX2 U11966 ( .A(n33184), .Z(n33182) );
  HS65_LH_BFX2 U11967 ( .A(n33178), .Z(n33183) );
  HS65_LH_BFX2 U11968 ( .A(n33186), .Z(n33184) );
  HS65_LH_BFX2 U11969 ( .A(n33183), .Z(n33185) );
  HS65_LH_BFX2 U11970 ( .A(n33188), .Z(n33186) );
  HS65_LH_BFX2 U11971 ( .A(n33185), .Z(n33187) );
  HS65_LH_BFX2 U11972 ( .A(n33190), .Z(n33188) );
  HS65_LH_BFX2 U11973 ( .A(n33187), .Z(n33189) );
  HS65_LH_BFX2 U11974 ( .A(n33192), .Z(n33190) );
  HS65_LH_BFX2 U11975 ( .A(n33189), .Z(n33191) );
  HS65_LH_BFX2 U11976 ( .A(n33194), .Z(n33192) );
  HS65_LH_BFX2 U11977 ( .A(n33191), .Z(n33193) );
  HS65_LH_BFX2 U11978 ( .A(n33196), .Z(n33194) );
  HS65_LH_BFX2 U11979 ( .A(n33193), .Z(n33195) );
  HS65_LH_BFX2 U11980 ( .A(n33198), .Z(n33196) );
  HS65_LH_BFX2 U11981 ( .A(n33195), .Z(n33197) );
  HS65_LH_BFX2 U11982 ( .A(n33200), .Z(n33198) );
  HS65_LH_BFX2 U11983 ( .A(n33197), .Z(n33199) );
  HS65_LH_BFX2 U11984 ( .A(n33203), .Z(n33200) );
  HS65_LH_BFX2 U11985 ( .A(n33199), .Z(n33201) );
  HS65_LH_IVX2 U11986 ( .A(n33208), .Z(n33202) );
  HS65_LH_IVX2 U11987 ( .A(n33202), .Z(n33203) );
  HS65_LH_BFX2 U11988 ( .A(n33201), .Z(n33204) );
  HS65_LH_IVX2 U11989 ( .A(n33211), .Z(n33205) );
  HS65_LH_IVX2 U11990 ( .A(n33205), .Z(n33206) );
  HS65_LH_IVX2 U11991 ( .A(n33210), .Z(n33207) );
  HS65_LH_IVX2 U11992 ( .A(n33207), .Z(n33208) );
  HS65_LH_IVX2 U11993 ( .A(n1634), .Z(n33209) );
  HS65_LH_IVX2 U11994 ( .A(n33209), .Z(n33210) );
  HS65_LH_BFX2 U11995 ( .A(n33212), .Z(n33211) );
  HS65_LH_BFX2 U11996 ( .A(n33204), .Z(n33212) );
  HS65_LH_BFX2 U11997 ( .A(n33214), .Z(n33213) );
  HS65_LH_BFX2 U11998 ( .A(n33215), .Z(n33214) );
  HS65_LH_BFX2 U11999 ( .A(n33216), .Z(n33215) );
  HS65_LH_BFX2 U12000 ( .A(n33217), .Z(n33216) );
  HS65_LH_BFX2 U12001 ( .A(n33218), .Z(n33217) );
  HS65_LH_BFX2 U12002 ( .A(n33219), .Z(n33218) );
  HS65_LH_BFX2 U12003 ( .A(n33220), .Z(n33219) );
  HS65_LH_BFX2 U12004 ( .A(n33221), .Z(n33220) );
  HS65_LH_BFX2 U12005 ( .A(n33222), .Z(n33221) );
  HS65_LH_BFX2 U12006 ( .A(n33223), .Z(n33222) );
  HS65_LH_BFX2 U12007 ( .A(n33224), .Z(n33223) );
  HS65_LH_BFX2 U12008 ( .A(n33225), .Z(n33224) );
  HS65_LH_BFX2 U12009 ( .A(n33226), .Z(n33225) );
  HS65_LH_BFX2 U12010 ( .A(n15719), .Z(n33226) );
  HS65_LH_BFX2 U12011 ( .A(n15392), .Z(n33227) );
  HS65_LH_BFX2 U12012 ( .A(n33230), .Z(n33228) );
  HS65_LH_BFX2 U12013 ( .A(n15544), .Z(n33229) );
  HS65_LH_BFX2 U12014 ( .A(n33251), .Z(n33230) );
  HS65_LH_BFX2 U12015 ( .A(n33229), .Z(n33231) );
  HS65_LH_BFX2 U12016 ( .A(n17966), .Z(n33232) );
  HS65_LH_BFX2 U12017 ( .A(n33231), .Z(n33233) );
  HS65_LH_BFX2 U12018 ( .A(n33232), .Z(n33234) );
  HS65_LH_BFX2 U12019 ( .A(n33233), .Z(n33235) );
  HS65_LH_BFX2 U12020 ( .A(n33234), .Z(n33236) );
  HS65_LH_BFX2 U12021 ( .A(n33235), .Z(n33237) );
  HS65_LH_BFX2 U12022 ( .A(n33236), .Z(n33238) );
  HS65_LH_BFX2 U12023 ( .A(n33237), .Z(n33239) );
  HS65_LH_BFX2 U12024 ( .A(n33238), .Z(n33240) );
  HS65_LH_BFX2 U12025 ( .A(n33239), .Z(n33241) );
  HS65_LH_BFX2 U12026 ( .A(n33240), .Z(n33242) );
  HS65_LH_BFX2 U12027 ( .A(n33241), .Z(n33243) );
  HS65_LH_BFX2 U12028 ( .A(n33242), .Z(n33244) );
  HS65_LH_BFX2 U12029 ( .A(n33243), .Z(n33245) );
  HS65_LH_BFX2 U12030 ( .A(n33244), .Z(n33246) );
  HS65_LH_BFX2 U12031 ( .A(n33245), .Z(n33247) );
  HS65_LH_BFX2 U12032 ( .A(n33246), .Z(n33248) );
  HS65_LH_BFX2 U12033 ( .A(n33247), .Z(n33249) );
  HS65_LH_IVX2 U12034 ( .A(n33256), .Z(n33250) );
  HS65_LH_IVX2 U12035 ( .A(n33250), .Z(n33251) );
  HS65_LH_BFX2 U12036 ( .A(n33249), .Z(n33252) );
  HS65_LH_IVX2 U12037 ( .A(n14448), .Z(n33253) );
  HS65_LH_IVX2 U12038 ( .A(n33253), .Z(n33254) );
  HS65_LH_IVX2 U12039 ( .A(n33261), .Z(n33255) );
  HS65_LH_IVX2 U12040 ( .A(n33255), .Z(n33256) );
  HS65_LH_BFX2 U12041 ( .A(n33252), .Z(n33257) );
  HS65_LH_IVX2 U12042 ( .A(n33264), .Z(n33258) );
  HS65_LH_IVX2 U12043 ( .A(n33258), .Z(n33259) );
  HS65_LH_IVX2 U12044 ( .A(n33263), .Z(n33260) );
  HS65_LH_IVX2 U12045 ( .A(n33260), .Z(n33261) );
  HS65_LH_IVX2 U12046 ( .A(n33265), .Z(n33262) );
  HS65_LH_IVX2 U12047 ( .A(n33262), .Z(n33263) );
  HS65_LH_BFX2 U12048 ( .A(n33257), .Z(n33264) );
  HS65_LH_BFX2 U12049 ( .A(n33266), .Z(n33265) );
  HS65_LH_BFX2 U12050 ( .A(n33267), .Z(n33266) );
  HS65_LH_BFX2 U12051 ( .A(n33268), .Z(n33267) );
  HS65_LH_BFX2 U12052 ( .A(n33269), .Z(n33268) );
  HS65_LH_BFX2 U12053 ( .A(n33270), .Z(n33269) );
  HS65_LH_BFX2 U12055 ( .A(n33248), .Z(n33270) );
  HS65_LH_BFX2 U12056 ( .A(n33273), .Z(n33271) );
  HS65_LH_BFX2 U12057 ( .A(n33274), .Z(n33272) );
  HS65_LH_BFX2 U12058 ( .A(n33275), .Z(n33273) );
  HS65_LH_BFX2 U12059 ( .A(n33276), .Z(n33274) );
  HS65_LH_BFX2 U12060 ( .A(n33277), .Z(n33275) );
  HS65_LH_BFX2 U12061 ( .A(n33278), .Z(n33276) );
  HS65_LH_BFX2 U12062 ( .A(n33279), .Z(n33277) );
  HS65_LH_BFX2 U12063 ( .A(n33280), .Z(n33278) );
  HS65_LH_BFX2 U12064 ( .A(n33281), .Z(n33279) );
  HS65_LH_BFX2 U12065 ( .A(n33282), .Z(n33280) );
  HS65_LH_BFX2 U12066 ( .A(n33283), .Z(n33281) );
  HS65_LH_BFX2 U12067 ( .A(n33284), .Z(n33282) );
  HS65_LH_BFX2 U12068 ( .A(n33285), .Z(n33283) );
  HS65_LH_BFX2 U12069 ( .A(n33286), .Z(n33284) );
  HS65_LH_BFX2 U12070 ( .A(n33287), .Z(n33285) );
  HS65_LH_BFX2 U12071 ( .A(n33288), .Z(n33286) );
  HS65_LH_BFX2 U12072 ( .A(n33289), .Z(n33287) );
  HS65_LH_BFX2 U12073 ( .A(n33290), .Z(n33288) );
  HS65_LH_BFX2 U12074 ( .A(n33291), .Z(n33289) );
  HS65_LH_BFX2 U12075 ( .A(n33292), .Z(n33290) );
  HS65_LH_BFX2 U12076 ( .A(n33293), .Z(n33291) );
  HS65_LH_BFX2 U12077 ( .A(n33294), .Z(n33292) );
  HS65_LH_BFX2 U12078 ( .A(n33295), .Z(n33293) );
  HS65_LH_BFX2 U12079 ( .A(n33296), .Z(n33294) );
  HS65_LH_BFX2 U12080 ( .A(n33297), .Z(n33295) );
  HS65_LH_BFX2 U12081 ( .A(n33298), .Z(n33296) );
  HS65_LH_BFX2 U12082 ( .A(n33299), .Z(n33297) );
  HS65_LH_BFX2 U12083 ( .A(n33300), .Z(n33298) );
  HS65_LH_BFX2 U12084 ( .A(n33301), .Z(n33299) );
  HS65_LH_BFX2 U12085 ( .A(n1725), .Z(n33300) );
  HS65_LH_BFX2 U12086 ( .A(n1726), .Z(n33301) );
  HS65_LH_BFX2 U12087 ( .A(n33307), .Z(n33302) );
  HS65_LH_BFX2 U12088 ( .A(n2597), .Z(n33303) );
  HS65_LH_BFX2 U12089 ( .A(n36170), .Z(n33304) );
  HS65_LH_BFX2 U12090 ( .A(n15870), .Z(n33305) );
  HS65_LH_BFX2 U12091 ( .A(n33303), .Z(n33306) );
  HS65_LH_BFX2 U12092 ( .A(n33309), .Z(n33307) );
  HS65_LH_BFX2 U12093 ( .A(n33306), .Z(n33308) );
  HS65_LH_BFX2 U12094 ( .A(n33311), .Z(n33309) );
  HS65_LH_BFX2 U12095 ( .A(n33308), .Z(n33310) );
  HS65_LH_BFX2 U12096 ( .A(n33313), .Z(n33311) );
  HS65_LH_BFX2 U12097 ( .A(n33310), .Z(n33312) );
  HS65_LH_BFX2 U12098 ( .A(n33315), .Z(n33313) );
  HS65_LH_BFX2 U12099 ( .A(n33312), .Z(n33314) );
  HS65_LH_BFX2 U12100 ( .A(n33317), .Z(n33315) );
  HS65_LH_BFX2 U12101 ( .A(n33314), .Z(n33316) );
  HS65_LH_BFX2 U12102 ( .A(n33319), .Z(n33317) );
  HS65_LH_BFX2 U12103 ( .A(n33316), .Z(n33318) );
  HS65_LH_BFX2 U12104 ( .A(n33321), .Z(n33319) );
  HS65_LH_BFX2 U12105 ( .A(n33318), .Z(n33320) );
  HS65_LH_BFX2 U12106 ( .A(n33323), .Z(n33321) );
  HS65_LH_BFX2 U12107 ( .A(n33320), .Z(n33322) );
  HS65_LH_BFX2 U12108 ( .A(n33325), .Z(n33323) );
  HS65_LH_BFX2 U12109 ( .A(n33322), .Z(n33324) );
  HS65_LH_BFX2 U12110 ( .A(n33328), .Z(n33325) );
  HS65_LH_BFX2 U12111 ( .A(n33324), .Z(n33326) );
  HS65_LH_IVX2 U12112 ( .A(n2598), .Z(n33327) );
  HS65_LH_IVX2 U12113 ( .A(n33327), .Z(n33328) );
  HS65_LH_BFX2 U12114 ( .A(n33326), .Z(n33329) );
  HS65_LH_IVX2 U12115 ( .A(n33332), .Z(n33330) );
  HS65_LH_IVX2 U12116 ( .A(n33330), .Z(n33331) );
  HS65_LH_BFX2 U12117 ( .A(n33329), .Z(n33332) );
  HS65_LH_BFX2 U12118 ( .A(n33335), .Z(n33333) );
  HS65_LH_IVX2 U12119 ( .A(n33338), .Z(n33334) );
  HS65_LH_IVX2 U12120 ( .A(n33334), .Z(n33335) );
  HS65_LH_BFX2 U12121 ( .A(n2621), .Z(n33336) );
  HS65_LH_BFX2 U12122 ( .A(n33336), .Z(n33337) );
  HS65_LH_BFX2 U12123 ( .A(n33340), .Z(n33338) );
  HS65_LH_BFX2 U12124 ( .A(n33337), .Z(n33339) );
  HS65_LH_BFX2 U12125 ( .A(n33342), .Z(n33340) );
  HS65_LH_BFX2 U12126 ( .A(n33339), .Z(n33341) );
  HS65_LH_BFX2 U12127 ( .A(n33344), .Z(n33342) );
  HS65_LH_BFX2 U12128 ( .A(n33341), .Z(n33343) );
  HS65_LH_BFX2 U12129 ( .A(n33346), .Z(n33344) );
  HS65_LH_BFX2 U12130 ( .A(n33343), .Z(n33345) );
  HS65_LH_BFX2 U12131 ( .A(n33348), .Z(n33346) );
  HS65_LH_BFX2 U12132 ( .A(n33345), .Z(n33347) );
  HS65_LH_BFX2 U12133 ( .A(n33350), .Z(n33348) );
  HS65_LH_BFX2 U12134 ( .A(n33347), .Z(n33349) );
  HS65_LH_BFX2 U12135 ( .A(n33352), .Z(n33350) );
  HS65_LH_BFX2 U12136 ( .A(n33349), .Z(n33351) );
  HS65_LH_BFX2 U12137 ( .A(n33354), .Z(n33352) );
  HS65_LH_BFX2 U12138 ( .A(n33351), .Z(n33353) );
  HS65_LH_BFX2 U12139 ( .A(n33356), .Z(n33354) );
  HS65_LH_BFX2 U12140 ( .A(n33353), .Z(n33355) );
  HS65_LH_BFX2 U12141 ( .A(n33358), .Z(n33356) );
  HS65_LH_BFX2 U12142 ( .A(n33355), .Z(n33357) );
  HS65_LH_BFX2 U12143 ( .A(n33360), .Z(n33358) );
  HS65_LH_BFX2 U12144 ( .A(n33357), .Z(n33359) );
  HS65_LH_BFX2 U12145 ( .A(n33364), .Z(n33360) );
  HS65_LH_BFX2 U12146 ( .A(n33359), .Z(n33361) );
  HS65_LH_IVX2 U12147 ( .A(n33361), .Z(n33362) );
  HS65_LH_IVX2 U12148 ( .A(n33362), .Z(n33363) );
  HS65_LH_BFX2 U12149 ( .A(n2622), .Z(n33364) );
  HS65_LH_IVX2 U12150 ( .A(n33603), .Z(n33365) );
  HS65_LH_IVX2 U12151 ( .A(n33365), .Z(n33366) );
  HS65_LH_BFX2 U12152 ( .A(n33369), .Z(n33367) );
  HS65_LH_BFX2 U12153 ( .A(n1656), .Z(n33368) );
  HS65_LH_BFX2 U12154 ( .A(n33371), .Z(n33369) );
  HS65_LH_BFX2 U12155 ( .A(n33368), .Z(n33370) );
  HS65_LH_BFX2 U12156 ( .A(n33373), .Z(n33371) );
  HS65_LH_BFX2 U12157 ( .A(n33370), .Z(n33372) );
  HS65_LH_BFX2 U12158 ( .A(n33375), .Z(n33373) );
  HS65_LH_BFX2 U12159 ( .A(n33372), .Z(n33374) );
  HS65_LH_BFX2 U12160 ( .A(n33377), .Z(n33375) );
  HS65_LH_BFX2 U12161 ( .A(n33374), .Z(n33376) );
  HS65_LH_BFX2 U12162 ( .A(n33379), .Z(n33377) );
  HS65_LH_BFX2 U12163 ( .A(n33376), .Z(n33378) );
  HS65_LH_BFX2 U12164 ( .A(n33381), .Z(n33379) );
  HS65_LH_BFX2 U12165 ( .A(n33378), .Z(n33380) );
  HS65_LH_BFX2 U12166 ( .A(n33383), .Z(n33381) );
  HS65_LH_BFX2 U12167 ( .A(n33380), .Z(n33382) );
  HS65_LH_BFX2 U12168 ( .A(n33385), .Z(n33383) );
  HS65_LH_BFX2 U12169 ( .A(n33382), .Z(n33384) );
  HS65_LH_BFX2 U12170 ( .A(n33387), .Z(n33385) );
  HS65_LH_BFX2 U12171 ( .A(n33384), .Z(n33386) );
  HS65_LH_BFX2 U12172 ( .A(n33389), .Z(n33387) );
  HS65_LH_BFX2 U12173 ( .A(n33386), .Z(n33388) );
  HS65_LH_BFX2 U12174 ( .A(n33392), .Z(n33389) );
  HS65_LH_BFX2 U12175 ( .A(n33388), .Z(n33390) );
  HS65_LH_IVX2 U12176 ( .A(n33397), .Z(n33391) );
  HS65_LH_IVX2 U12177 ( .A(n33391), .Z(n33392) );
  HS65_LH_BFX2 U12178 ( .A(n33390), .Z(n33393) );
  HS65_LH_IVX2 U12179 ( .A(n33393), .Z(n33394) );
  HS65_LH_IVX2 U12180 ( .A(n33394), .Z(n33395) );
  HS65_LH_IVX2 U12181 ( .A(n33399), .Z(n33396) );
  HS65_LH_IVX2 U12182 ( .A(n33396), .Z(n33397) );
  HS65_LH_IVX2 U12183 ( .A(n1657), .Z(n33398) );
  HS65_LH_IVX2 U12184 ( .A(n33398), .Z(n33399) );
  HS65_LH_BFX2 U12185 ( .A(n33405), .Z(n33400) );
  HS65_LH_BFX2 U12186 ( .A(n1679), .Z(n33401) );
  HS65_LH_BFX2 U12187 ( .A(n33404), .Z(n33402) );
  HS65_LH_IVX2 U12188 ( .A(n33412), .Z(n33403) );
  HS65_LH_IVX2 U12189 ( .A(n33403), .Z(n33404) );
  HS65_LH_BFX2 U12190 ( .A(n33413), .Z(n33405) );
  HS65_LH_BFX2 U12191 ( .A(n33401), .Z(n33406) );
  HS65_LH_IVX2 U12192 ( .A(n33430), .Z(n33407) );
  HS65_LH_IVX2 U12193 ( .A(n33407), .Z(n33408) );
  HS65_LH_IVX2 U12194 ( .A(n33415), .Z(n33409) );
  HS65_LH_IVX2 U12195 ( .A(n33409), .Z(n33410) );
  HS65_LH_IVX2 U12196 ( .A(n33606), .Z(n33411) );
  HS65_LH_IVX2 U12197 ( .A(n33411), .Z(n33412) );
  HS65_LH_BFX2 U12198 ( .A(n33414), .Z(n33413) );
  HS65_LH_BFX2 U12199 ( .A(n33416), .Z(n33414) );
  HS65_LH_BFX2 U12200 ( .A(n33417), .Z(n33415) );
  HS65_LH_BFX2 U12201 ( .A(n33418), .Z(n33416) );
  HS65_LH_BFX2 U12202 ( .A(n33419), .Z(n33417) );
  HS65_LH_BFX2 U12203 ( .A(n33420), .Z(n33418) );
  HS65_LH_BFX2 U12204 ( .A(n33421), .Z(n33419) );
  HS65_LH_BFX2 U12205 ( .A(n33422), .Z(n33420) );
  HS65_LH_BFX2 U12206 ( .A(n33423), .Z(n33421) );
  HS65_LH_BFX2 U12207 ( .A(n33424), .Z(n33422) );
  HS65_LH_BFX2 U12208 ( .A(n33425), .Z(n33423) );
  HS65_LH_BFX2 U12209 ( .A(n33426), .Z(n33424) );
  HS65_LH_BFX2 U12210 ( .A(n33427), .Z(n33425) );
  HS65_LH_BFX2 U12211 ( .A(n33428), .Z(n33426) );
  HS65_LH_BFX2 U12212 ( .A(n33434), .Z(n33427) );
  HS65_LH_BFX2 U12213 ( .A(n33429), .Z(n33428) );
  HS65_LH_BFX2 U12214 ( .A(n33431), .Z(n33429) );
  HS65_LH_BFX2 U12215 ( .A(n33432), .Z(n33430) );
  HS65_LH_BFX2 U12216 ( .A(n33433), .Z(n33431) );
  HS65_LH_BFX2 U12219 ( .A(n16662), .Z(n33432) );
  HS65_LH_BFX2 U12220 ( .A(n33435), .Z(n33433) );
  HS65_LH_BFX2 U12221 ( .A(n33406), .Z(n33434) );
  HS65_LH_BFX2 U12222 ( .A(n1680), .Z(n33435) );
  HS65_LH_BFX2 U12223 ( .A(n33441), .Z(n33436) );
  HS65_LH_BFX2 U12224 ( .A(n1702), .Z(n33437) );
  HS65_LH_BFX2 U12225 ( .A(n33440), .Z(n33438) );
  HS65_LH_IVX2 U12226 ( .A(n33827), .Z(n33439) );
  HS65_LH_IVX2 U12227 ( .A(n33439), .Z(n33440) );
  HS65_LH_BFX2 U12228 ( .A(n33443), .Z(n33441) );
  HS65_LH_BFX2 U12229 ( .A(n33437), .Z(n33442) );
  HS65_LH_BFX2 U12230 ( .A(n33445), .Z(n33443) );
  HS65_LH_BFX2 U12231 ( .A(n33442), .Z(n33444) );
  HS65_LH_BFX2 U12232 ( .A(n33447), .Z(n33445) );
  HS65_LH_BFX2 U12233 ( .A(n33444), .Z(n33446) );
  HS65_LH_BFX2 U12234 ( .A(n33449), .Z(n33447) );
  HS65_LH_BFX2 U12235 ( .A(n33446), .Z(n33448) );
  HS65_LH_BFX2 U12241 ( .A(n33451), .Z(n33449) );
  HS65_LH_BFX2 U12242 ( .A(n33448), .Z(n33450) );
  HS65_LH_BFX2 U12243 ( .A(n33453), .Z(n33451) );
  HS65_LH_BFX2 U12244 ( .A(n33450), .Z(n33452) );
  HS65_LH_BFX2 U12245 ( .A(n33455), .Z(n33453) );
  HS65_LH_BFX2 U12246 ( .A(n33452), .Z(n33454) );
  HS65_LH_BFX2 U12247 ( .A(n33457), .Z(n33455) );
  HS65_LH_BFX2 U12248 ( .A(n33454), .Z(n33456) );
  HS65_LH_BFX2 U12249 ( .A(n33459), .Z(n33457) );
  HS65_LH_BFX2 U12250 ( .A(n33456), .Z(n33458) );
  HS65_LH_BFX2 U12251 ( .A(n33461), .Z(n33459) );
  HS65_LH_BFX2 U12252 ( .A(n33458), .Z(n33460) );
  HS65_LH_BFX2 U12253 ( .A(n33464), .Z(n33461) );
  HS65_LH_BFX2 U12254 ( .A(n33460), .Z(n33462) );
  HS65_LH_IVX2 U12255 ( .A(n33469), .Z(n33463) );
  HS65_LH_IVX2 U12263 ( .A(n33463), .Z(n33464) );
  HS65_LH_BFX2 U12264 ( .A(n33462), .Z(n33465) );
  HS65_LH_IVX2 U12265 ( .A(n33465), .Z(n33466) );
  HS65_LH_IVX2 U12266 ( .A(n33466), .Z(n33467) );
  HS65_LH_IVX2 U12267 ( .A(n33470), .Z(n33468) );
  HS65_LH_IVX2 U12268 ( .A(n33468), .Z(n33469) );
  HS65_LH_BFX2 U12269 ( .A(n1703), .Z(n33470) );
  HS65_LH_BFX2 U12270 ( .A(n33477), .Z(n33471) );
  HS65_LH_BFX2 U12271 ( .A(n33474), .Z(n33472) );
  HS65_LH_BFX2 U12272 ( .A(n15550), .Z(n33473) );
  HS65_LH_BFX2 U12273 ( .A(n33476), .Z(n33474) );
  HS65_LH_BFX2 U12274 ( .A(n33473), .Z(n33475) );
  HS65_LH_BFX2 U12285 ( .A(n33478), .Z(n33476) );
  HS65_LH_BFX2 U12286 ( .A(n33479), .Z(n33477) );
  HS65_LH_BFX2 U12287 ( .A(n33480), .Z(n33478) );
  HS65_LH_BFX2 U12288 ( .A(n33481), .Z(n33479) );
  HS65_LH_BFX2 U12289 ( .A(n33482), .Z(n33480) );
  HS65_LH_BFX2 U12290 ( .A(n33483), .Z(n33481) );
  HS65_LH_BFX2 U12291 ( .A(n33484), .Z(n33482) );
  HS65_LH_BFX2 U12292 ( .A(n33485), .Z(n33483) );
  HS65_LH_BFX2 U12293 ( .A(n33486), .Z(n33484) );
  HS65_LH_BFX2 U12294 ( .A(n33487), .Z(n33485) );
  HS65_LH_BFX2 U12307 ( .A(n33488), .Z(n33486) );
  HS65_LH_BFX2 U12308 ( .A(n33489), .Z(n33487) );
  HS65_LH_BFX2 U12309 ( .A(n33490), .Z(n33488) );
  HS65_LH_BFX2 U12310 ( .A(n33491), .Z(n33489) );
  HS65_LH_BFX2 U12311 ( .A(n33492), .Z(n33490) );
  HS65_LH_BFX2 U12312 ( .A(n33493), .Z(n33491) );
  HS65_LH_BFX2 U12313 ( .A(n33494), .Z(n33492) );
  HS65_LH_BFX2 U12329 ( .A(n33495), .Z(n33493) );
  HS65_LH_BFX2 U12330 ( .A(n33496), .Z(n33494) );
  HS65_LH_BFX2 U12331 ( .A(n33497), .Z(n33495) );
  HS65_LH_BFX2 U12332 ( .A(n33498), .Z(n33496) );
  HS65_LH_BFX2 U12333 ( .A(n33499), .Z(n33497) );
  HS65_LH_BFX2 U12351 ( .A(n33500), .Z(n33498) );
  HS65_LH_BFX2 U12352 ( .A(n33503), .Z(n33499) );
  HS65_LH_BFX2 U12417 ( .A(n33502), .Z(n33500) );
  HS65_LH_BFX2 U12421 ( .A(n14789), .Z(n33501) );
  HS65_LH_BFX2 U12423 ( .A(n33504), .Z(n33502) );
  HS65_LH_BFX2 U12427 ( .A(n33475), .Z(n33503) );
  HS65_LH_BFX2 U12431 ( .A(n33506), .Z(n33504) );
  HS65_LH_BFX2 U12435 ( .A(n17470), .Z(n33505) );
  HS65_LH_BFX2 U12439 ( .A(n33507), .Z(n33506) );
  HS65_LH_BFX2 U12722 ( .A(n33508), .Z(n33507) );
  HS65_LH_BFX2 U12724 ( .A(n33509), .Z(n33508) );
  HS65_LH_BFX2 U12726 ( .A(n17921), .Z(n33509) );
  HS65_LH_BFX2 U12728 ( .A(n17820), .Z(n33510) );
  HS65_LH_BFX2 U12730 ( .A(n17819), .Z(n33511) );
  HS65_LH_IVX2 U12732 ( .A(n17251), .Z(n33512) );
  HS65_LH_IVX2 U12765 ( .A(n33512), .Z(n33513) );
  HS65_LH_BFX2 U12769 ( .A(n17869), .Z(n33514) );
  HS65_LH_BFX2 U12771 ( .A(n33514), .Z(n33515) );
  HS65_LH_IVX2 U12773 ( .A(n33520), .Z(n33516) );
  HS65_LH_IVX2 U12775 ( .A(n33516), .Z(n33517) );
  HS65_LH_IVX2 U12777 ( .A(n33521), .Z(n33518) );
  HS65_LH_IVX2 U12779 ( .A(n33518), .Z(n33519) );
  HS65_LH_BFX2 U12783 ( .A(n33522), .Z(n33520) );
  HS65_LH_BFX2 U12785 ( .A(n33523), .Z(n33521) );
  HS65_LH_BFX2 U12812 ( .A(n33524), .Z(n33522) );
  HS65_LH_BFX2 U12814 ( .A(n33525), .Z(n33523) );
  HS65_LH_BFX2 U12818 ( .A(n33526), .Z(n33524) );
  HS65_LH_BFX2 U12820 ( .A(n33527), .Z(n33525) );
  HS65_LH_BFX2 U12822 ( .A(n33528), .Z(n33526) );
  HS65_LH_BFX2 U12824 ( .A(n33529), .Z(n33527) );
  HS65_LH_BFX2 U12826 ( .A(n33530), .Z(n33528) );
  HS65_LH_BFX2 U12828 ( .A(n33531), .Z(n33529) );
  HS65_LH_BFX2 U12830 ( .A(n33532), .Z(n33530) );
  HS65_LH_BFX2 U12832 ( .A(n33533), .Z(n33531) );
  HS65_LH_BFX2 U12834 ( .A(n33534), .Z(n33532) );
  HS65_LH_BFX2 U12855 ( .A(n33535), .Z(n33533) );
  HS65_LH_BFX2 U12857 ( .A(n33536), .Z(n33534) );
  HS65_LH_BFX2 U12859 ( .A(n33537), .Z(n33535) );
  HS65_LH_BFX2 U12861 ( .A(n33538), .Z(n33536) );
  HS65_LH_BFX2 U12863 ( .A(n33539), .Z(n33537) );
  HS65_LH_BFX2 U12865 ( .A(n33540), .Z(n33538) );
  HS65_LH_BFX2 U12867 ( .A(n33541), .Z(n33539) );
  HS65_LH_BFX2 U12869 ( .A(n33542), .Z(n33540) );
  HS65_LH_BFX2 U12871 ( .A(n33543), .Z(n33541) );
  HS65_LH_BFX2 U12873 ( .A(n33544), .Z(n33542) );
  HS65_LH_BFX2 U12875 ( .A(n33545), .Z(n33543) );
  HS65_LH_BFX2 U12877 ( .A(n33546), .Z(n33544) );
  HS65_LH_BFX2 U12879 ( .A(n33547), .Z(n33545) );
  HS65_LH_BFX2 U12881 ( .A(n15545), .Z(n33546) );
  HS65_LH_BFX2 U12883 ( .A(n33548), .Z(n33547) );
  HS65_LH_BFX2 U12885 ( .A(n33549), .Z(n33548) );
  HS65_LH_BFX2 U12902 ( .A(n33550), .Z(n33549) );
  HS65_LH_BFX2 U12904 ( .A(n33551), .Z(n33550) );
  HS65_LH_BFX2 U12906 ( .A(n33515), .Z(n33551) );
  HS65_LH_BFX2 U12908 ( .A(n17987), .Z(n33552) );
  HS65_LH_BFX2 U12910 ( .A(n33555), .Z(n33553) );
  HS65_LH_BFX2 U12912 ( .A(n17928), .Z(n33554) );
  HS65_LH_BFX2 U12914 ( .A(n33559), .Z(n33555) );
  HS65_LH_BFX2 U12916 ( .A(n33554), .Z(n33556) );
  HS65_LH_IVX2 U12918 ( .A(n33561), .Z(n33557) );
  HS65_LH_IVX2 U12920 ( .A(n33557), .Z(n33558) );
  HS65_LH_BFX2 U12922 ( .A(n33560), .Z(n33559) );
  HS65_LH_BFX2 U12924 ( .A(n33562), .Z(n33560) );
  HS65_LH_BFX2 U12926 ( .A(n33563), .Z(n33561) );
  HS65_LH_BFX2 U12928 ( .A(n33564), .Z(n33562) );
  HS65_LH_BFX2 U12930 ( .A(n33565), .Z(n33563) );
  HS65_LH_BFX2 U12932 ( .A(n33566), .Z(n33564) );
  HS65_LH_BFX2 U12934 ( .A(n33567), .Z(n33565) );
  HS65_LH_BFX2 U12936 ( .A(n33568), .Z(n33566) );
  HS65_LH_BFX2 U12945 ( .A(n33569), .Z(n33567) );
  HS65_LH_BFX2 U12947 ( .A(n33570), .Z(n33568) );
  HS65_LH_BFX2 U12949 ( .A(n33571), .Z(n33569) );
  HS65_LH_BFX2 U12951 ( .A(n33572), .Z(n33570) );
  HS65_LH_BFX2 U12953 ( .A(n33573), .Z(n33571) );
  HS65_LH_BFX2 U12955 ( .A(n33574), .Z(n33572) );
  HS65_LH_BFX2 U12957 ( .A(n33575), .Z(n33573) );
  HS65_LH_BFX2 U12959 ( .A(n33576), .Z(n33574) );
  HS65_LH_BFX2 U12961 ( .A(n33577), .Z(n33575) );
  HS65_LH_BFX2 U12963 ( .A(n33578), .Z(n33576) );
  HS65_LH_BFX2 U12965 ( .A(n33579), .Z(n33577) );
  HS65_LH_BFX2 U12967 ( .A(n33580), .Z(n33578) );
  HS65_LH_BFX2 U12969 ( .A(n33581), .Z(n33579) );
  HS65_LH_BFX2 U12971 ( .A(n33582), .Z(n33580) );
  HS65_LH_BFX2 U12973 ( .A(n33583), .Z(n33581) );
  HS65_LH_BFX2 U12975 ( .A(n33584), .Z(n33582) );
  HS65_LH_BFX2 U12977 ( .A(n33585), .Z(n33583) );
  HS65_LH_BFX2 U12979 ( .A(n15540), .Z(n33584) );
  HS65_LH_BFX2 U12981 ( .A(n33586), .Z(n33585) );
  HS65_LH_BFX2 U12983 ( .A(n33587), .Z(n33586) );
  HS65_LH_BFX2 U12985 ( .A(n33588), .Z(n33587) );
  HS65_LH_BFX2 U12992 ( .A(n33589), .Z(n33588) );
  HS65_LH_BFX2 U12994 ( .A(n33590), .Z(n33589) );
  HS65_LH_BFX2 U12996 ( .A(n33556), .Z(n33590) );
  HS65_LH_BFX2 U12998 ( .A(n33592), .Z(n33591) );
  HS65_LH_BFX2 U13000 ( .A(n33593), .Z(n33592) );
  HS65_LH_BFX2 U13002 ( .A(n17983), .Z(n33593) );
  HS65_LH_BFX2 U13004 ( .A(n33595), .Z(n33594) );
  HS65_LH_BFX2 U13006 ( .A(n17949), .Z(n33595) );
  HS65_LH_BFX2 U13008 ( .A(n33597), .Z(n33596) );
  HS65_LH_BFX2 U13010 ( .A(n17980), .Z(n33597) );
  HS65_LH_BFX2 U13012 ( .A(n33599), .Z(n33598) );
  HS65_LH_BFX2 U13014 ( .A(n33600), .Z(n33599) );
  HS65_LH_BFX2 U13016 ( .A(n17943), .Z(n33600) );
  HS65_LH_BFX2 U13018 ( .A(n33602), .Z(n33601) );
  HS65_LH_BFX2 U13020 ( .A(n17968), .Z(n33602) );
  HS65_LH_BFX2 U13022 ( .A(n33604), .Z(n33603) );
  HS65_LH_BFX2 U13024 ( .A(n33605), .Z(n33604) );
  HS65_LH_BFX2 U13026 ( .A(n17922), .Z(n33605) );
  HS65_LH_BFX2 U13028 ( .A(n33607), .Z(n33606) );
  HS65_LH_BFX2 U13030 ( .A(n17897), .Z(n33607) );
  HS65_LH_IVX2 U13035 ( .A(n33612), .Z(n33608) );
  HS65_LH_IVX2 U13037 ( .A(n33608), .Z(n33609) );
  HS65_LH_BFX2 U13039 ( .A(n33611), .Z(n33610) );
  HS65_LH_BFX2 U13041 ( .A(n33613), .Z(n33611) );
  HS65_LH_BFX2 U13043 ( .A(n33614), .Z(n33612) );
  HS65_LH_BFX2 U13045 ( .A(n33615), .Z(n33613) );
  HS65_LH_BFX2 U13047 ( .A(n33616), .Z(n33614) );
  HS65_LH_BFX2 U13049 ( .A(n33617), .Z(n33615) );
  HS65_LH_BFX2 U13051 ( .A(n33618), .Z(n33616) );
  HS65_LH_BFX2 U13053 ( .A(n33619), .Z(n33617) );
  HS65_LH_BFX2 U13055 ( .A(n33620), .Z(n33618) );
  HS65_LH_BFX2 U13057 ( .A(n33621), .Z(n33619) );
  HS65_LH_BFX2 U13059 ( .A(n33622), .Z(n33620) );
  HS65_LH_BFX2 U13061 ( .A(n33623), .Z(n33621) );
  HS65_LH_BFX2 U13063 ( .A(n33624), .Z(n33622) );
  HS65_LH_BFX2 U13065 ( .A(n33625), .Z(n33623) );
  HS65_LH_BFX2 U13067 ( .A(n33626), .Z(n33624) );
  HS65_LH_BFX2 U13069 ( .A(n33627), .Z(n33625) );
  HS65_LH_BFX2 U13071 ( .A(n33628), .Z(n33626) );
  HS65_LH_BFX2 U13073 ( .A(n33629), .Z(n33627) );
  HS65_LH_BFX2 U13075 ( .A(n33630), .Z(n33628) );
  HS65_LH_BFX2 U13287 ( .A(n33631), .Z(n33629) );
  HS65_LH_BFX2 U14059 ( .A(n33632), .Z(n33630) );
  HS65_LH_BFX2 U14102 ( .A(n33633), .Z(n33631) );
  HS65_LH_BFX2 U14104 ( .A(n33634), .Z(n33632) );
  HS65_LH_BFX2 U14106 ( .A(n33635), .Z(n33633) );
  HS65_LH_BFX2 U14108 ( .A(n33636), .Z(n33634) );
  HS65_LH_BFX2 U14110 ( .A(n33637), .Z(n33635) );
  HS65_LH_BFX2 U14149 ( .A(n33638), .Z(n33636) );
  HS65_LH_BFX2 U14151 ( .A(n33639), .Z(n33637) );
  HS65_LH_BFX2 U14153 ( .A(n15546), .Z(n33638) );
  HS65_LH_BFX2 U14155 ( .A(n33641), .Z(n33639) );
  HS65_LH_BFX2 U14157 ( .A(n33643), .Z(n33640) );
  HS65_LH_BFX2 U14159 ( .A(n33642), .Z(n33641) );
  HS65_LH_BFX2 U14161 ( .A(n33644), .Z(n33642) );
  HS65_LH_BFX2 U14163 ( .A(n33070), .Z(n33643) );
  HS65_LH_BFX2 U14165 ( .A(n33645), .Z(n33644) );
  HS65_LH_BFX2 U14167 ( .A(n33646), .Z(n33645) );
  HS65_LH_BFX2 U14169 ( .A(n17945), .Z(n33646) );
  HS65_LH_BFX2 U14171 ( .A(n17823), .Z(n33647) );
  HS65_LH_BFX2 U14173 ( .A(n17821), .Z(n33648) );
  HS65_LH_BFX2 U14175 ( .A(n33650), .Z(n33649) );
  HS65_LH_BFX2 U14177 ( .A(n33651), .Z(n33650) );
  HS65_LH_BFX2 U14179 ( .A(n33652), .Z(n33651) );
  HS65_LH_BFX2 U14181 ( .A(n17888), .Z(n33652) );
  HS65_LH_BFX2 U14183 ( .A(\u_DataPath/dataOut_exe_i [30]), .Z(n33653) );
  HS65_LH_BFX2 U14185 ( .A(\u_DataPath/dataOut_exe_i [29]), .Z(n33654) );
  HS65_LH_BFX2 U14187 ( .A(n33689), .Z(n33655) );
  HS65_LH_BFX2 U14192 ( .A(n33658), .Z(n33656) );
  HS65_LH_IVX2 U14194 ( .A(n33661), .Z(n33657) );
  HS65_LH_IVX2 U14196 ( .A(n33657), .Z(n33658) );
  HS65_LH_BFX2 U14198 ( .A(n15549), .Z(n33659) );
  HS65_LH_IVX2 U14200 ( .A(n33664), .Z(n33660) );
  HS65_LH_IVX2 U14202 ( .A(n33660), .Z(n33661) );
  HS65_LH_BFX2 U14204 ( .A(n33659), .Z(n33662) );
  HS65_LH_BFX2 U14206 ( .A(n33662), .Z(n33663) );
  HS65_LH_BFX2 U14208 ( .A(n33666), .Z(n33664) );
  HS65_LH_BFX2 U14210 ( .A(n33663), .Z(n33665) );
  HS65_LH_BFX2 U14212 ( .A(n33668), .Z(n33666) );
  HS65_LH_BFX2 U14214 ( .A(n33665), .Z(n33667) );
  HS65_LH_BFX2 U14216 ( .A(n33670), .Z(n33668) );
  HS65_LH_BFX2 U14218 ( .A(n33667), .Z(n33669) );
  HS65_LH_BFX2 U14220 ( .A(n33672), .Z(n33670) );
  HS65_LH_BFX2 U14222 ( .A(n33669), .Z(n33671) );
  HS65_LH_BFX2 U14224 ( .A(n33674), .Z(n33672) );
  HS65_LH_BFX2 U14226 ( .A(n33671), .Z(n33673) );
  HS65_LH_BFX2 U14228 ( .A(n33676), .Z(n33674) );
  HS65_LH_BFX2 U14230 ( .A(n33673), .Z(n33675) );
  HS65_LH_BFX2 U14232 ( .A(n33678), .Z(n33676) );
  HS65_LH_BFX2 U14239 ( .A(n33675), .Z(n33677) );
  HS65_LH_BFX2 U14241 ( .A(n33680), .Z(n33678) );
  HS65_LH_BFX2 U14243 ( .A(n33677), .Z(n33679) );
  HS65_LH_BFX2 U14245 ( .A(n33682), .Z(n33680) );
  HS65_LH_BFX2 U14247 ( .A(n33679), .Z(n33681) );
  HS65_LH_BFX2 U14249 ( .A(n33684), .Z(n33682) );
  HS65_LH_BFX2 U14251 ( .A(n33681), .Z(n33683) );
  HS65_LH_BFX2 U14253 ( .A(n33686), .Z(n33684) );
  HS65_LH_BFX2 U14255 ( .A(n33683), .Z(n33685) );
  HS65_LH_BFX2 U14257 ( .A(n33690), .Z(n33686) );
  HS65_LH_BFX2 U14259 ( .A(n14961), .Z(n33687) );
  HS65_LH_IVX2 U14261 ( .A(n33685), .Z(n33688) );
  HS65_LH_IVX2 U14263 ( .A(n33688), .Z(n33689) );
  HS65_LH_BFX2 U14265 ( .A(n33692), .Z(n33690) );
  HS65_LH_IVX2 U14267 ( .A(n33694), .Z(n33691) );
  HS65_LH_IVX2 U14269 ( .A(n33691), .Z(n33692) );
  HS65_LH_BFX2 U14271 ( .A(n15202), .Z(n33693) );
  HS65_LH_BFX2 U14273 ( .A(n33695), .Z(n33694) );
  HS65_LH_BFX2 U14275 ( .A(n33696), .Z(n33695) );
  HS65_LH_BFX2 U14277 ( .A(n33697), .Z(n33696) );
  HS65_LH_BFX2 U14282 ( .A(n17896), .Z(n33697) );
  HS65_LH_BFX2 U14284 ( .A(n15541), .Z(n33698) );
  HS65_LH_BFX2 U14286 ( .A(n33701), .Z(n33699) );
  HS65_LH_BFX2 U14288 ( .A(n33698), .Z(n33700) );
  HS65_LH_BFX2 U14290 ( .A(n33703), .Z(n33701) );
  HS65_LH_BFX2 U14292 ( .A(n33700), .Z(n33702) );
  HS65_LH_BFX2 U14294 ( .A(n33705), .Z(n33703) );
  HS65_LH_BFX2 U14296 ( .A(n33702), .Z(n33704) );
  HS65_LH_BFX2 U14298 ( .A(n33707), .Z(n33705) );
  HS65_LH_BFX2 U14300 ( .A(n33704), .Z(n33706) );
  HS65_LH_BFX2 U14302 ( .A(n33709), .Z(n33707) );
  HS65_LH_BFX2 U14304 ( .A(n33706), .Z(n33708) );
  HS65_LH_BFX2 U14306 ( .A(n33711), .Z(n33709) );
  HS65_LH_BFX2 U14308 ( .A(n33708), .Z(n33710) );
  HS65_LH_BFX2 U14310 ( .A(n33713), .Z(n33711) );
  HS65_LH_BFX2 U14312 ( .A(n33710), .Z(n33712) );
  HS65_LH_BFX2 U14314 ( .A(n33715), .Z(n33713) );
  HS65_LH_BFX2 U14316 ( .A(n33712), .Z(n33714) );
  HS65_LH_BFX2 U14318 ( .A(n33717), .Z(n33715) );
  HS65_LH_BFX2 U14320 ( .A(n33714), .Z(n33716) );
  HS65_LH_BFX2 U14322 ( .A(n33719), .Z(n33717) );
  HS65_LH_BFX2 U14330 ( .A(n33716), .Z(n33718) );
  HS65_LH_BFX2 U14335 ( .A(n33721), .Z(n33719) );
  HS65_LH_BFX2 U14336 ( .A(n33718), .Z(n33720) );
  HS65_LH_BFX2 U14344 ( .A(n33723), .Z(n33721) );
  HS65_LH_BFX2 U14345 ( .A(n33720), .Z(n33722) );
  HS65_LH_BFX2 U14346 ( .A(n33725), .Z(n33723) );
  HS65_LH_BFX2 U14354 ( .A(n33722), .Z(n33724) );
  HS65_LH_BFX2 U14355 ( .A(n33727), .Z(n33725) );
  HS65_LH_BFX2 U14356 ( .A(n33724), .Z(n33726) );
  HS65_LH_BFX2 U14363 ( .A(n33730), .Z(n33727) );
  HS65_LH_BFX2 U14364 ( .A(n14940), .Z(n33728) );
  HS65_LH_IVX2 U14365 ( .A(n33733), .Z(n33729) );
  HS65_LH_IVX2 U14372 ( .A(n33729), .Z(n33730) );
  HS65_LH_IVX2 U14373 ( .A(n33726), .Z(n33731) );
  HS65_LH_IVX2 U14374 ( .A(n33731), .Z(n33732) );
  HS65_LH_BFX2 U14381 ( .A(n33734), .Z(n33733) );
  HS65_LH_BFX2 U14382 ( .A(n33735), .Z(n33734) );
  HS65_LH_BFX2 U14389 ( .A(n33736), .Z(n33735) );
  HS65_LH_BFX2 U14396 ( .A(n33737), .Z(n33736) );
  HS65_LH_BFX2 U14399 ( .A(n17899), .Z(n33737) );
  HS65_LH_BFX2 U14403 ( .A(n33739), .Z(n33738) );
  HS65_LH_BFX2 U14409 ( .A(n33740), .Z(n33739) );
  HS65_LH_BFX2 U14412 ( .A(n33741), .Z(n33740) );
  HS65_LH_BFX2 U14416 ( .A(n33742), .Z(n33741) );
  HS65_LH_BFX2 U14418 ( .A(n17883), .Z(n33742) );
  HS65_LH_BFX2 U14421 ( .A(n33744), .Z(n33743) );
  HS65_LH_BFX2 U14424 ( .A(n33745), .Z(n33744) );
  HS65_LH_BFX2 U14426 ( .A(n33746), .Z(n33745) );
  HS65_LH_BFX2 U14428 ( .A(n33747), .Z(n33746) );
  HS65_LH_BFX2 U14430 ( .A(n17873), .Z(n33747) );
  HS65_LH_IVX2 U14432 ( .A(n17265), .Z(n33748) );
  HS65_LH_IVX2 U14435 ( .A(n33748), .Z(n33749) );
  HS65_LH_BFX2 U14439 ( .A(n33751), .Z(n33750) );
  HS65_LH_BFX2 U14452 ( .A(n26577), .Z(n33751) );
  HS65_LH_BFX2 U14465 ( .A(n33753), .Z(n33752) );
  HS65_LH_BFX2 U14478 ( .A(n33754), .Z(n33753) );
  HS65_LH_BFX2 U14491 ( .A(n33755), .Z(n33754) );
  HS65_LH_BFX2 U14504 ( .A(n33756), .Z(n33755) );
  HS65_LH_BFX2 U14517 ( .A(n17933), .Z(n33756) );
  HS65_LH_BFX2 U14530 ( .A(n33758), .Z(n33757) );
  HS65_LH_BFX2 U14543 ( .A(n33759), .Z(n33758) );
  HS65_LH_BFX2 U14555 ( .A(n14802), .Z(n33759) );
  HS65_LH_BFX2 U14566 ( .A(n33761), .Z(n33760) );
  HS65_LH_BFX2 U14579 ( .A(n33762), .Z(n33761) );
  HS65_LH_BFX2 U14592 ( .A(n33763), .Z(n33762) );
  HS65_LH_BFX2 U14605 ( .A(n33764), .Z(n33763) );
  HS65_LH_BFX2 U14618 ( .A(n17976), .Z(n33764) );
  HS65_LH_BFX2 U14630 ( .A(n33766), .Z(n33765) );
  HS65_LH_BFX2 U14641 ( .A(n33767), .Z(n33766) );
  HS65_LH_BFX2 U14654 ( .A(n33768), .Z(n33767) );
  HS65_LH_BFX2 U14667 ( .A(n33769), .Z(n33768) );
  HS65_LH_BFX2 U14692 ( .A(n17907), .Z(n33769) );
  HS65_LH_BFX2 U14724 ( .A(n14213), .Z(n33770) );
  HS65_LH_BFX2 U14799 ( .A(\u_DataPath/dataOut_exe_i [27]), .Z(n33771) );
  HS65_LH_BFX2 U14830 ( .A(n33773), .Z(n33772) );
  HS65_LH_BFX2 U14882 ( .A(n33774), .Z(n33773) );
  HS65_LH_BFX2 U14886 ( .A(n14747), .Z(n33774) );
  HS65_LH_BFX2 U14888 ( .A(n14452), .Z(n33775) );
  HS65_LH_BFX2 U14928 ( .A(\u_DataPath/dataOut_exe_i [26]), .Z(n33776) );
  HS65_LH_BFX2 U14932 ( .A(n33778), .Z(n33777) );
  HS65_LH_BFX2 U14939 ( .A(n33779), .Z(n33778) );
  HS65_LH_BFX2 U14950 ( .A(n33780), .Z(n33779) );
  HS65_LH_BFX2 U14965 ( .A(n33781), .Z(n33780) );
  HS65_LH_BFX2 U15004 ( .A(n33782), .Z(n33781) );
  HS65_LH_BFX2 U15025 ( .A(n17893), .Z(n33782) );
  HS65_LH_BFX2 U15112 ( .A(n33784), .Z(n33783) );
  HS65_LH_BFX2 U15113 ( .A(n26759), .Z(n33784) );
  HS65_LH_BFX2 U15114 ( .A(\u_DataPath/dataOut_exe_i [28]), .Z(n33785) );
  HS65_LH_BFX2 U15170 ( .A(n15537), .Z(n33786) );
  HS65_LH_BFX2 U15311 ( .A(n33789), .Z(n33787) );
  HS65_LH_BFX2 U15313 ( .A(n33786), .Z(n33788) );
  HS65_LH_BFX2 U15314 ( .A(n33791), .Z(n33789) );
  HS65_LH_BFX2 U15322 ( .A(n33788), .Z(n33790) );
  HS65_LH_BFX2 U15337 ( .A(n33793), .Z(n33791) );
  HS65_LH_BFX2 U15345 ( .A(n33790), .Z(n33792) );
  HS65_LH_BFX2 U15358 ( .A(n33795), .Z(n33793) );
  HS65_LH_BFX2 U15393 ( .A(n33792), .Z(n33794) );
  HS65_LH_BFX2 U15647 ( .A(n33797), .Z(n33795) );
  HS65_LH_BFX2 U15780 ( .A(n33798), .Z(n33796) );
  HS65_LH_BFX2 U15863 ( .A(n33799), .Z(n33797) );
  HS65_LH_BFX2 U15864 ( .A(n33800), .Z(n33798) );
  HS65_LH_BFX2 U15887 ( .A(n33801), .Z(n33799) );
  HS65_LH_BFX2 U15888 ( .A(n33802), .Z(n33800) );
  HS65_LH_BFX2 U16017 ( .A(n33803), .Z(n33801) );
  HS65_LH_BFX2 U16148 ( .A(n33804), .Z(n33802) );
  HS65_LH_BFX2 U16401 ( .A(n33805), .Z(n33803) );
  HS65_LH_BFX2 U16513 ( .A(n33806), .Z(n33804) );
  HS65_LH_BFX2 U16524 ( .A(n33807), .Z(n33805) );
  HS65_LH_BFX2 U16525 ( .A(n33808), .Z(n33806) );
  HS65_LH_BFX2 U16526 ( .A(n33809), .Z(n33807) );
  HS65_LH_BFX2 U16528 ( .A(n33810), .Z(n33808) );
  HS65_LH_BFX2 U16544 ( .A(n33811), .Z(n33809) );
  HS65_LH_BFX2 U16597 ( .A(n33812), .Z(n33810) );
  HS65_LH_BFX2 U16600 ( .A(n33813), .Z(n33811) );
  HS65_LH_BFX2 U16601 ( .A(n33814), .Z(n33812) );
  HS65_LH_BFX2 U16603 ( .A(n33815), .Z(n33813) );
  HS65_LH_BFX2 U16617 ( .A(n33816), .Z(n33814) );
  HS65_LH_BFX2 U16625 ( .A(n33817), .Z(n33815) );
  HS65_LH_BFX2 U16628 ( .A(n33818), .Z(n33816) );
  HS65_LH_BFX2 U16632 ( .A(n33819), .Z(n33817) );
  HS65_LH_BFX2 U16634 ( .A(n33794), .Z(n33818) );
  HS65_LH_BFX2 U16637 ( .A(n33820), .Z(n33819) );
  HS65_LH_BFX2 U16642 ( .A(n33821), .Z(n33820) );
  HS65_LH_BFX2 U16654 ( .A(n33822), .Z(n33821) );
  HS65_LH_BFX2 U16664 ( .A(n33823), .Z(n33822) );
  HS65_LH_BFX2 U16666 ( .A(n17970), .Z(n33823) );
  HS65_LH_BFX2 U16669 ( .A(n33825), .Z(n33824) );
  HS65_LH_BFX2 U16676 ( .A(n33826), .Z(n33825) );
  HS65_LH_BFX2 U16677 ( .A(n17870), .Z(n33826) );
  HS65_LH_BFX2 U16680 ( .A(n33828), .Z(n33827) );
  HS65_LH_BFX2 U16682 ( .A(n17946), .Z(n33828) );
  HS65_LH_BFX2 U16686 ( .A(n33831), .Z(n33829) );
  HS65_LH_BFX2 U16688 ( .A(n33832), .Z(n33830) );
  HS65_LH_BFX2 U16689 ( .A(n17792), .Z(n33831) );
  HS65_LH_BFX2 U16693 ( .A(n33833), .Z(n33832) );
  HS65_LH_BFX2 U16696 ( .A(n33834), .Z(n33833) );
  HS65_LH_BFX2 U16704 ( .A(n33835), .Z(n33834) );
  HS65_LH_BFX2 U16708 ( .A(n33836), .Z(n33835) );
  HS65_LH_BFX2 U16712 ( .A(n33837), .Z(n33836) );
  HS65_LH_BFX2 U16717 ( .A(n33838), .Z(n33837) );
  HS65_LH_BFX2 U16720 ( .A(n33839), .Z(n33838) );
  HS65_LH_BFX2 U16722 ( .A(n33840), .Z(n33839) );
  HS65_LH_BFX2 U16738 ( .A(n33841), .Z(n33840) );
  HS65_LH_BFX2 U16749 ( .A(n33842), .Z(n33841) );
  HS65_LH_BFX2 U16775 ( .A(n33843), .Z(n33842) );
  HS65_LH_BFX2 U16789 ( .A(n33844), .Z(n33843) );
  HS65_LH_BFX2 U16808 ( .A(n33845), .Z(n33844) );
  HS65_LH_BFX2 U16811 ( .A(n33846), .Z(n33845) );
  HS65_LH_BFX2 U16822 ( .A(n33847), .Z(n33846) );
  HS65_LH_BFX2 U16833 ( .A(n33848), .Z(n33847) );
  HS65_LH_BFX2 U16852 ( .A(n17585), .Z(n33848) );
  HS65_LH_BFX2 U16874 ( .A(n33858), .Z(n33849) );
  HS65_LH_BFX2 U16899 ( .A(n33852), .Z(n33850) );
  HS65_LH_IVX2 U16937 ( .A(n33855), .Z(n33851) );
  HS65_LH_IVX2 U16938 ( .A(n33851), .Z(n33852) );
  HS65_LH_BFX2 U16965 ( .A(n15538), .Z(n33853) );
  HS65_LH_BFX2 U16976 ( .A(n33853), .Z(n33854) );
  HS65_LH_BFX2 U16998 ( .A(n33857), .Z(n33855) );
  HS65_LH_BFX2 U17031 ( .A(n33854), .Z(n33856) );
  HS65_LH_BFX2 U17042 ( .A(n33859), .Z(n33857) );
  HS65_LH_BFX2 U17050 ( .A(n33860), .Z(n33858) );
  HS65_LH_BFX2 U17078 ( .A(n33861), .Z(n33859) );
  HS65_LH_BFX2 U17086 ( .A(n33862), .Z(n33860) );
  HS65_LH_BFX2 U17097 ( .A(n33863), .Z(n33861) );
  HS65_LH_BFX2 U17127 ( .A(n33864), .Z(n33862) );
  HS65_LH_BFX2 U17130 ( .A(n33865), .Z(n33863) );
  HS65_LH_BFX2 U17171 ( .A(n33866), .Z(n33864) );
  HS65_LH_BFX2 U17181 ( .A(n33867), .Z(n33865) );
  HS65_LH_BFX2 U17190 ( .A(n33868), .Z(n33866) );
  HS65_LH_BFX2 U17196 ( .A(n33869), .Z(n33867) );
  HS65_LH_BFX2 U17234 ( .A(n33870), .Z(n33868) );
  HS65_LH_BFX2 U17256 ( .A(n33871), .Z(n33869) );
  HS65_LH_BFX2 U17257 ( .A(n33872), .Z(n33870) );
  HS65_LH_BFX2 U17267 ( .A(n33873), .Z(n33871) );
  HS65_LH_BFX2 U17278 ( .A(n33874), .Z(n33872) );
  HS65_LH_BFX2 U17328 ( .A(n33875), .Z(n33873) );
  HS65_LH_BFX2 U17346 ( .A(n33876), .Z(n33874) );
  HS65_LH_BFX2 U17358 ( .A(n33877), .Z(n33875) );
  HS65_LH_BFX2 U17367 ( .A(n33878), .Z(n33876) );
  HS65_LH_BFX2 U17455 ( .A(n33879), .Z(n33877) );
  HS65_LH_BFX2 U17464 ( .A(n33856), .Z(n33878) );
  HS65_LH_BFX2 U17465 ( .A(n33881), .Z(n33879) );
  HS65_LH_BFX2 U17467 ( .A(n17592), .Z(n33880) );
  HS65_LH_BFX2 U17517 ( .A(n33883), .Z(n33881) );
  HS65_LH_BFX2 U17539 ( .A(n17315), .Z(n33882) );
  HS65_LH_BFX2 U17558 ( .A(n33884), .Z(n33883) );
  HS65_LH_BFX2 U17561 ( .A(n33885), .Z(n33884) );
  HS65_LH_BFX2 U17580 ( .A(n33886), .Z(n33885) );
  HS65_LH_BFX2 U17628 ( .A(n33887), .Z(n33886) );
  HS65_LH_BFX2 U17650 ( .A(n17876), .Z(n33887) );
  HS65_LH_BFX2 U17669 ( .A(n338), .Z(n33888) );
  HS65_LH_BFX2 U17735 ( .A(n33890), .Z(n33889) );
  HS65_LH_BFX2 U17760 ( .A(n33891), .Z(n33890) );
  HS65_LH_BFX2 U17779 ( .A(n33892), .Z(n33891) );
  HS65_LH_BFX2 U17782 ( .A(n17852), .Z(n33892) );
  HS65_LH_BFX2 U17787 ( .A(n33895), .Z(n33893) );
  HS65_LH_IVX2 U17801 ( .A(n326), .Z(n33894) );
  HS65_LH_IVX2 U17804 ( .A(n33894), .Z(n33895) );
  HS65_LH_BFX2 U17812 ( .A(n33897), .Z(n33896) );
  HS65_LH_BFX2 U17832 ( .A(n33898), .Z(n33897) );
  HS65_LH_BFX2 U17892 ( .A(n33899), .Z(n33898) );
  HS65_LH_BFX2 U17900 ( .A(n33900), .Z(n33899) );
  HS65_LH_BFX2 U17936 ( .A(n17929), .Z(n33900) );
  HS65_LH_BFX2 U17985 ( .A(n33903), .Z(n33901) );
  HS65_LH_IVX2 U17988 ( .A(n327), .Z(n33902) );
  HS65_LH_IVX2 U17999 ( .A(n33902), .Z(n33903) );
  HS65_LH_BFX2 U18010 ( .A(n33905), .Z(n33904) );
  HS65_LH_BFX2 U18043 ( .A(n33906), .Z(n33905) );
  HS65_LH_BFX2 U18052 ( .A(n33907), .Z(n33906) );
  HS65_LH_BFX2 U18068 ( .A(n33908), .Z(n33907) );
  HS65_LH_BFX2 U18076 ( .A(n17900), .Z(n33908) );
  HS65_LH_BFX2 U18079 ( .A(n33911), .Z(n33909) );
  HS65_LH_BFX2 U18098 ( .A(n33912), .Z(n33910) );
  HS65_LH_BFX2 U18109 ( .A(n330), .Z(n33911) );
  HS65_LH_BFX2 U18139 ( .A(n33913), .Z(n33912) );
  HS65_LH_BFX2 U18170 ( .A(n33914), .Z(n33913) );
  HS65_LH_BFX2 U18171 ( .A(n33915), .Z(n33914) );
  HS65_LH_BFX2 U18172 ( .A(n17759), .Z(n33915) );
  HS65_LH_BFX2 U18173 ( .A(n33919), .Z(n33916) );
  HS65_LH_BFX2 U18174 ( .A(n17268), .Z(n33917) );
  HS65_LH_BFX2 U18175 ( .A(n33921), .Z(n33918) );
  HS65_LH_BFX2 U18176 ( .A(n33922), .Z(n33919) );
  HS65_LH_BFX2 U18177 ( .A(n33917), .Z(n33920) );
  HS65_LH_BFX2 U18178 ( .A(n33926), .Z(n33921) );
  HS65_LH_BFX2 U18179 ( .A(n33925), .Z(n33922) );
  HS65_LH_BFX2 U18180 ( .A(n33920), .Z(n33923) );
  HS65_LH_IVX2 U18181 ( .A(n33931), .Z(n33924) );
  HS65_LH_IVX2 U18182 ( .A(n33924), .Z(n33925) );
  HS65_LH_BFX2 U18183 ( .A(n33932), .Z(n33926) );
  HS65_LH_BFX2 U18184 ( .A(n33923), .Z(n33927) );
  HS65_LH_IVX2 U18185 ( .A(n33927), .Z(n33928) );
  HS65_LH_IVX2 U18186 ( .A(n33928), .Z(n33929) );
  HS65_LH_IVX2 U18187 ( .A(n17848), .Z(n33930) );
  HS65_LH_IVX2 U18188 ( .A(n33930), .Z(n33931) );
  HS65_LH_BFX2 U18189 ( .A(n17303), .Z(n33932) );
  HS65_LH_IVX2 U18190 ( .A(n33937), .Z(n33933) );
  HS65_LH_IVX2 U18191 ( .A(n33933), .Z(n33934) );
  HS65_LH_BFX2 U18192 ( .A(n33936), .Z(n33935) );
  HS65_LH_BFX2 U18193 ( .A(n33938), .Z(n33936) );
  HS65_LH_BFX2 U18194 ( .A(n328), .Z(n33937) );
  HS65_LH_BFX2 U18195 ( .A(n33939), .Z(n33938) );
  HS65_LH_BFX2 U18196 ( .A(n33940), .Z(n33939) );
  HS65_LH_BFX2 U18197 ( .A(n33941), .Z(n33940) );
  HS65_LH_BFX2 U18198 ( .A(n17971), .Z(n33941) );
  HS65_LH_BFX2 U18199 ( .A(n33955), .Z(n33942) );
  HS65_LH_BFX2 U18200 ( .A(n33946), .Z(n33943) );
  HS65_LH_BFX2 U18201 ( .A(n17854), .Z(n33944) );
  HS65_LH_IVX2 U18202 ( .A(n17857), .Z(n33945) );
  HS65_LH_IVX2 U18203 ( .A(n33945), .Z(n33946) );
  HS65_LH_BFX2 U18204 ( .A(n33949), .Z(n33947) );
  HS65_LH_IVX2 U18205 ( .A(n17509), .Z(n33948) );
  HS65_LH_IVX2 U18206 ( .A(n33948), .Z(n33949) );
  HS65_LH_BFX2 U18207 ( .A(n33956), .Z(n33950) );
  HS65_LH_BFX2 U18208 ( .A(n17858), .Z(n33951) );
  HS65_LH_BFX2 U18209 ( .A(n33954), .Z(n33952) );
  HS65_LH_IVX2 U18210 ( .A(n329), .Z(n33953) );
  HS65_LH_IVX2 U18211 ( .A(n33953), .Z(n33954) );
  HS65_LH_BFX2 U18212 ( .A(n17568), .Z(n33955) );
  HS65_LH_BFX2 U18213 ( .A(n33957), .Z(n33956) );
  HS65_LH_BFX2 U18214 ( .A(n33958), .Z(n33957) );
  HS65_LH_BFX2 U18215 ( .A(n33959), .Z(n33958) );
  HS65_LH_BFX2 U18216 ( .A(n33960), .Z(n33959) );
  HS65_LH_BFX2 U18217 ( .A(n17878), .Z(n33960) );
  HS65_LH_BFX2 U18218 ( .A(n33963), .Z(n33961) );
  HS65_LH_IVX2 U18219 ( .A(n33967), .Z(n33962) );
  HS65_LH_IVX2 U18220 ( .A(n33962), .Z(n33963) );
  HS65_LH_BFX2 U18221 ( .A(n34023), .Z(n33964) );
  HS65_LH_BFX2 U18222 ( .A(n33966), .Z(n33965) );
  HS65_LH_BFX2 U18223 ( .A(n34022), .Z(n33966) );
  HS65_LH_BFX2 U18224 ( .A(n33968), .Z(n33967) );
  HS65_LH_BFX2 U18225 ( .A(n34024), .Z(n33968) );
  HS65_LH_BFX2 U18226 ( .A(n34267), .Z(n33969) );
  HS65_LH_IVX2 U18227 ( .A(n33975), .Z(n33970) );
  HS65_LH_IVX2 U18228 ( .A(n33970), .Z(n33971) );
  HS65_LH_IVX2 U18229 ( .A(n33977), .Z(n33972) );
  HS65_LH_IVX2 U18230 ( .A(n33972), .Z(n33973) );
  HS65_LH_IVX2 U18231 ( .A(n33979), .Z(n33974) );
  HS65_LH_IVX2 U18232 ( .A(n33974), .Z(n33975) );
  HS65_LH_IVX2 U18233 ( .A(n33981), .Z(n33976) );
  HS65_LH_IVX2 U18234 ( .A(n33976), .Z(n33977) );
  HS65_LH_IVX2 U18235 ( .A(n33983), .Z(n33978) );
  HS65_LH_IVX2 U18236 ( .A(n33978), .Z(n33979) );
  HS65_LH_IVX2 U18237 ( .A(n33985), .Z(n33980) );
  HS65_LH_IVX2 U18238 ( .A(n33980), .Z(n33981) );
  HS65_LH_IVX2 U18239 ( .A(n33987), .Z(n33982) );
  HS65_LH_IVX2 U18240 ( .A(n33982), .Z(n33983) );
  HS65_LH_IVX2 U18241 ( .A(n33989), .Z(n33984) );
  HS65_LH_IVX2 U18242 ( .A(n33984), .Z(n33985) );
  HS65_LH_IVX2 U18243 ( .A(n33992), .Z(n33986) );
  HS65_LH_IVX2 U18244 ( .A(n33986), .Z(n33987) );
  HS65_LH_IVX2 U18245 ( .A(n33991), .Z(n33988) );
  HS65_LH_IVX2 U18246 ( .A(n33988), .Z(n33989) );
  HS65_LH_IVX2 U18247 ( .A(n17775), .Z(n33990) );
  HS65_LH_IVX2 U18248 ( .A(n33990), .Z(n33991) );
  HS65_LH_BFX2 U18249 ( .A(n33994), .Z(n33992) );
  HS65_LH_IVX2 U18250 ( .A(n17577), .Z(n33993) );
  HS65_LH_IVX2 U18251 ( .A(n33993), .Z(n33994) );
  HS65_LH_BFX2 U18252 ( .A(n33998), .Z(n33995) );
  HS65_LH_BFX2 U18253 ( .A(n17445), .Z(n33996) );
  HS65_LH_IVX2 U18254 ( .A(n34007), .Z(n33997) );
  HS65_LH_IVX2 U18255 ( .A(n33997), .Z(n33998) );
  HS65_LH_BFX2 U18256 ( .A(n36976), .Z(n33999) );
  HS65_LH_BFX2 U18257 ( .A(n17642), .Z(n34000) );
  HS65_LH_IVX2 U18258 ( .A(n34000), .Z(n34001) );
  HS65_LH_IVX2 U18259 ( .A(n34001), .Z(n34002) );
  HS65_LH_BFX2 U18260 ( .A(n33996), .Z(n34003) );
  HS65_LH_IVX2 U18261 ( .A(n34010), .Z(n34004) );
  HS65_LH_IVX2 U18262 ( .A(n34004), .Z(n34005) );
  HS65_LH_IVX2 U18263 ( .A(n34009), .Z(n34006) );
  HS65_LH_IVX2 U18264 ( .A(n34006), .Z(n34007) );
  HS65_LH_IVX2 U18265 ( .A(n17643), .Z(n34008) );
  HS65_LH_IVX2 U18266 ( .A(n34008), .Z(n34009) );
  HS65_LH_BFX2 U18267 ( .A(n34011), .Z(n34010) );
  HS65_LH_BFX2 U18268 ( .A(n34003), .Z(n34011) );
  HS65_LH_BFX2 U18269 ( .A(n17826), .Z(n34012) );
  HS65_LH_BFX2 U18270 ( .A(n33096), .Z(n34013) );
  HS65_LH_BFX2 U18271 ( .A(n17743), .Z(n34014) );
  HS65_LH_BFX2 U18272 ( .A(n17744), .Z(n34015) );
  HS65_LH_BFX2 U18273 ( .A(n34018), .Z(n34016) );
  HS65_LH_BFX2 U18274 ( .A(n34019), .Z(n34017) );
  HS65_LH_BFX2 U18275 ( .A(n34020), .Z(n34018) );
  HS65_LH_BFX2 U18276 ( .A(n34021), .Z(n34019) );
  HS65_LH_BFX2 U18277 ( .A(n17440), .Z(n34020) );
  HS65_LH_BFX2 U18278 ( .A(n17446), .Z(n34021) );
  HS65_LH_BFX2 U18279 ( .A(n34025), .Z(n34022) );
  HS65_LH_BFX2 U18280 ( .A(n34026), .Z(n34023) );
  HS65_LH_BFX2 U18281 ( .A(n34027), .Z(n34024) );
  HS65_LH_BFX2 U18282 ( .A(n34030), .Z(n34025) );
  HS65_LH_BFX2 U18283 ( .A(n34029), .Z(n34026) );
  HS65_LH_BFX2 U18284 ( .A(n17786), .Z(n34027) );
  HS65_LH_IVX2 U18285 ( .A(n34031), .Z(n34028) );
  HS65_LH_IVX2 U18286 ( .A(n34028), .Z(n34029) );
  HS65_LH_BFX2 U18287 ( .A(n17777), .Z(n34030) );
  HS65_LH_BFX2 U18288 ( .A(n17776), .Z(n34031) );
  HS65_LH_BFX2 U18289 ( .A(n34369), .Z(n34032) );
  HS65_LH_BFX2 U18290 ( .A(n34035), .Z(n34033) );
  HS65_LH_BFX2 U18291 ( .A(n2669), .Z(n34034) );
  HS65_LH_BFX2 U18292 ( .A(n34037), .Z(n34035) );
  HS65_LH_BFX2 U18293 ( .A(n34034), .Z(n34036) );
  HS65_LH_BFX2 U18294 ( .A(n34039), .Z(n34037) );
  HS65_LH_BFX2 U18295 ( .A(n34036), .Z(n34038) );
  HS65_LH_BFX2 U18296 ( .A(n34041), .Z(n34039) );
  HS65_LH_BFX2 U18297 ( .A(n34038), .Z(n34040) );
  HS65_LH_BFX2 U18298 ( .A(n34044), .Z(n34041) );
  HS65_LH_BFX2 U18299 ( .A(n34040), .Z(n34042) );
  HS65_LH_IVX2 U18300 ( .A(n34049), .Z(n34043) );
  HS65_LH_IVX2 U18301 ( .A(n34043), .Z(n34044) );
  HS65_LH_BFX2 U18302 ( .A(n34042), .Z(n34045) );
  HS65_LH_IVX2 U18303 ( .A(n34045), .Z(n34046) );
  HS65_LH_IVX2 U18304 ( .A(n34046), .Z(n34047) );
  HS65_LH_IVX2 U18305 ( .A(n2670), .Z(n34048) );
  HS65_LH_IVX2 U18306 ( .A(n34048), .Z(n34049) );
  HS65_LH_IVX2 U18307 ( .A(n34073), .Z(n34050) );
  HS65_LH_IVX2 U18308 ( .A(n34050), .Z(n34051) );
  HS65_LH_BFX2 U18309 ( .A(n34149), .Z(n34052) );
  HS65_LH_BFX2 U18310 ( .A(n34057), .Z(n34053) );
  HS65_LH_BFX2 U18311 ( .A(n34059), .Z(n34054) );
  HS65_LH_IVX2 U18312 ( .A(n17762), .Z(n34251) );
  HS65_LH_BFX2 U18313 ( .A(n34062), .Z(n34055) );
  HS65_LH_IVX2 U18314 ( .A(n34076), .Z(n34056) );
  HS65_LH_IVX2 U18315 ( .A(n34056), .Z(n34057) );
  HS65_LH_IVX2 U18316 ( .A(n34078), .Z(n34058) );
  HS65_LH_IVX2 U18317 ( .A(n34058), .Z(n34059) );
  HS65_LH_BFX2 U18318 ( .A(n34065), .Z(n34060) );
  HS65_LH_IVX2 U18319 ( .A(n34080), .Z(n34061) );
  HS65_LH_IVX2 U18320 ( .A(n34061), .Z(n34062) );
  HS65_LH_BFX2 U18321 ( .A(n34067), .Z(n34063) );
  HS65_LH_IVX2 U18322 ( .A(n34082), .Z(n34064) );
  HS65_LH_IVX2 U18323 ( .A(n34064), .Z(n34065) );
  HS65_LH_IVX2 U18324 ( .A(n34085), .Z(n34066) );
  HS65_LH_IVX2 U18325 ( .A(n34066), .Z(n34067) );
  HS65_LH_BFX2 U18326 ( .A(n17856), .Z(n34068) );
  HS65_LH_BFX2 U18327 ( .A(n34071), .Z(n34069) );
  HS65_LH_IVX2 U18328 ( .A(n34087), .Z(n34070) );
  HS65_LH_IVX2 U18329 ( .A(n34070), .Z(n34071) );
  HS65_LH_IVX2 U18330 ( .A(n34089), .Z(n34072) );
  HS65_LH_IVX2 U18331 ( .A(n34072), .Z(n34073) );
  HS65_LH_BFX2 U18332 ( .A(n324), .Z(n34074) );
  HS65_LH_IVX2 U18333 ( .A(n34092), .Z(n34075) );
  HS65_LH_IVX2 U18334 ( .A(n34075), .Z(n34076) );
  HS65_LH_IVX2 U18335 ( .A(n34094), .Z(n34077) );
  HS65_LH_IVX2 U18336 ( .A(n34077), .Z(n34078) );
  HS65_LH_IVX2 U18337 ( .A(n34096), .Z(n34079) );
  HS65_LH_IVX2 U18338 ( .A(n34079), .Z(n34080) );
  HS65_LH_IVX2 U18339 ( .A(n34099), .Z(n34081) );
  HS65_LH_IVX2 U18340 ( .A(n34081), .Z(n34082) );
  HS65_LH_BFX2 U18341 ( .A(n34068), .Z(n34083) );
  HS65_LH_IVX2 U18342 ( .A(n34101), .Z(n34084) );
  HS65_LH_IVX2 U18343 ( .A(n34084), .Z(n34085) );
  HS65_LH_IVX2 U18344 ( .A(n34103), .Z(n34086) );
  HS65_LH_IVX2 U18345 ( .A(n34086), .Z(n34087) );
  HS65_LH_IVX2 U18346 ( .A(n34105), .Z(n34088) );
  HS65_LH_IVX2 U18347 ( .A(n34088), .Z(n34089) );
  HS65_LH_BFX2 U18348 ( .A(n34074), .Z(n34090) );
  HS65_LH_IVX2 U18349 ( .A(n34108), .Z(n34091) );
  HS65_LH_IVX2 U18350 ( .A(n34091), .Z(n34092) );
  HS65_LH_IVX2 U18351 ( .A(n34111), .Z(n34093) );
  HS65_LH_IVX2 U18352 ( .A(n34093), .Z(n34094) );
  HS65_LH_IVX2 U18353 ( .A(n34113), .Z(n34095) );
  HS65_LH_IVX2 U18354 ( .A(n34095), .Z(n34096) );
  HS65_LH_BFX2 U18355 ( .A(n34083), .Z(n34097) );
  HS65_LH_IVX2 U18356 ( .A(n34115), .Z(n34098) );
  HS65_LH_IVX2 U18357 ( .A(n34098), .Z(n34099) );
  HS65_LH_IVX2 U18358 ( .A(n34117), .Z(n34100) );
  HS65_LH_IVX2 U18359 ( .A(n34100), .Z(n34101) );
  HS65_LH_IVX2 U18360 ( .A(n34119), .Z(n34102) );
  HS65_LH_IVX2 U18361 ( .A(n34102), .Z(n34103) );
  HS65_LH_IVX2 U18362 ( .A(n34122), .Z(n34104) );
  HS65_LH_IVX2 U18363 ( .A(n34104), .Z(n34105) );
  HS65_LH_BFX2 U18364 ( .A(n34090), .Z(n34106) );
  HS65_LH_IVX2 U18365 ( .A(n34137), .Z(n34107) );
  HS65_LH_IVX2 U18366 ( .A(n34107), .Z(n34108) );
  HS65_LH_BFX2 U18367 ( .A(n34097), .Z(n34109) );
  HS65_LH_IVX2 U18368 ( .A(n34125), .Z(n34110) );
  HS65_LH_IVX2 U18369 ( .A(n34110), .Z(n34111) );
  HS65_LH_IVX2 U18370 ( .A(n34127), .Z(n34112) );
  HS65_LH_IVX2 U18371 ( .A(n34112), .Z(n34113) );
  HS65_LH_IVX2 U18372 ( .A(n34129), .Z(n34114) );
  HS65_LH_IVX2 U18373 ( .A(n34114), .Z(n34115) );
  HS65_LH_IVX2 U18374 ( .A(n34131), .Z(n34116) );
  HS65_LH_IVX2 U18375 ( .A(n34116), .Z(n34117) );
  HS65_LH_IVX2 U18376 ( .A(n34134), .Z(n34118) );
  HS65_LH_IVX2 U18377 ( .A(n34118), .Z(n34119) );
  HS65_LH_BFX2 U18378 ( .A(n34106), .Z(n34120) );
  HS65_LH_IVX2 U18379 ( .A(n34136), .Z(n34121) );
  HS65_LH_IVX2 U18380 ( .A(n34121), .Z(n34122) );
  HS65_LH_BFX2 U18381 ( .A(n34109), .Z(n34123) );
  HS65_LH_IVX2 U18382 ( .A(n34140), .Z(n34124) );
  HS65_LH_IVX2 U18383 ( .A(n34124), .Z(n34125) );
  HS65_LH_IVX2 U18384 ( .A(n34142), .Z(n34126) );
  HS65_LH_IVX2 U18385 ( .A(n34126), .Z(n34127) );
  HS65_LH_IVX2 U18386 ( .A(n34144), .Z(n34128) );
  HS65_LH_IVX2 U18387 ( .A(n34128), .Z(n34129) );
  HS65_LH_IVX2 U18388 ( .A(n34146), .Z(n34130) );
  HS65_LH_IVX2 U18389 ( .A(n34130), .Z(n34131) );
  HS65_LH_BFX2 U18390 ( .A(n34120), .Z(n34132) );
  HS65_LH_IVX2 U18391 ( .A(n34151), .Z(n34133) );
  HS65_LH_IVX2 U18392 ( .A(n34133), .Z(n34134) );
  HS65_LH_IVX2 U18393 ( .A(n34153), .Z(n34135) );
  HS65_LH_IVX2 U18394 ( .A(n34135), .Z(n34136) );
  HS65_LH_BFX2 U18395 ( .A(n34154), .Z(n34137) );
  HS65_LH_BFX2 U18396 ( .A(n34123), .Z(n34138) );
  HS65_LH_IVX2 U18397 ( .A(n34157), .Z(n34139) );
  HS65_LH_IVX2 U18398 ( .A(n34139), .Z(n34140) );
  HS65_LH_IVX2 U18399 ( .A(n34159), .Z(n34141) );
  HS65_LH_IVX2 U18400 ( .A(n34141), .Z(n34142) );
  HS65_LH_IVX2 U18401 ( .A(n34161), .Z(n34143) );
  HS65_LH_IVX2 U18402 ( .A(n34143), .Z(n34144) );
  HS65_LH_IVX2 U18403 ( .A(n34163), .Z(n34145) );
  HS65_LH_IVX2 U18404 ( .A(n34145), .Z(n34146) );
  HS65_LH_BFX2 U18405 ( .A(n34132), .Z(n34147) );
  HS65_LH_IVX2 U18406 ( .A(n34165), .Z(n34148) );
  HS65_LH_IVX2 U18407 ( .A(n34148), .Z(n34149) );
  HS65_LH_IVX2 U18408 ( .A(n34167), .Z(n34150) );
  HS65_LH_IVX2 U18409 ( .A(n34150), .Z(n34151) );
  HS65_LH_IVX2 U18410 ( .A(n34169), .Z(n34152) );
  HS65_LH_IVX2 U18411 ( .A(n34152), .Z(n34153) );
  HS65_LH_BFX2 U18412 ( .A(n34170), .Z(n34154) );
  HS65_LH_BFX2 U18413 ( .A(n34138), .Z(n34155) );
  HS65_LH_IVX2 U18414 ( .A(n34177), .Z(n34156) );
  HS65_LH_IVX2 U18415 ( .A(n34156), .Z(n34157) );
  HS65_LH_IVX2 U18416 ( .A(n34179), .Z(n34158) );
  HS65_LH_IVX2 U18417 ( .A(n34158), .Z(n34159) );
  HS65_LH_IVX2 U18418 ( .A(n34181), .Z(n34160) );
  HS65_LH_IVX2 U18419 ( .A(n34160), .Z(n34161) );
  HS65_LH_IVX2 U18420 ( .A(n34183), .Z(n34162) );
  HS65_LH_IVX2 U18421 ( .A(n34162), .Z(n34163) );
  HS65_LH_IVX2 U18422 ( .A(n34185), .Z(n34164) );
  HS65_LH_IVX2 U18423 ( .A(n34164), .Z(n34165) );
  HS65_LH_IVX2 U18424 ( .A(n34187), .Z(n34166) );
  HS65_LH_IVX2 U18425 ( .A(n34166), .Z(n34167) );
  HS65_LH_IVX2 U18426 ( .A(n34189), .Z(n34168) );
  HS65_LH_IVX2 U18427 ( .A(n34168), .Z(n34169) );
  HS65_LH_BFX2 U18428 ( .A(n34173), .Z(n34170) );
  HS65_LH_BFX2 U18429 ( .A(n34155), .Z(n34171) );
  HS65_LH_IVX2 U18430 ( .A(n34205), .Z(n34172) );
  HS65_LH_IVX2 U18431 ( .A(n34172), .Z(n34173) );
  HS65_LH_IVX2 U18432 ( .A(n34247), .Z(n34174) );
  HS65_LH_IVX2 U18433 ( .A(n34174), .Z(n34175) );
  HS65_LH_IVX2 U18434 ( .A(n34191), .Z(n34176) );
  HS65_LH_IVX2 U18435 ( .A(n34176), .Z(n34177) );
  HS65_LH_IVX2 U18436 ( .A(n34193), .Z(n34178) );
  HS65_LH_IVX2 U18437 ( .A(n34178), .Z(n34179) );
  HS65_LH_IVX2 U18438 ( .A(n34195), .Z(n34180) );
  HS65_LH_IVX2 U18439 ( .A(n34180), .Z(n34181) );
  HS65_LH_IVX2 U18440 ( .A(n34197), .Z(n34182) );
  HS65_LH_IVX2 U18441 ( .A(n34182), .Z(n34183) );
  HS65_LH_IVX2 U18442 ( .A(n34199), .Z(n34184) );
  HS65_LH_IVX2 U18443 ( .A(n34184), .Z(n34185) );
  HS65_LH_IVX2 U18444 ( .A(n34201), .Z(n34186) );
  HS65_LH_IVX2 U18445 ( .A(n34186), .Z(n34187) );
  HS65_LH_IVX2 U18446 ( .A(n34203), .Z(n34188) );
  HS65_LH_IVX2 U18447 ( .A(n34188), .Z(n34189) );
  HS65_LH_IVX2 U18448 ( .A(n34209), .Z(n34190) );
  HS65_LH_IVX2 U18449 ( .A(n34190), .Z(n34191) );
  HS65_LH_IVX2 U18450 ( .A(n34211), .Z(n34192) );
  HS65_LH_IVX2 U18451 ( .A(n34192), .Z(n34193) );
  HS65_LH_IVX2 U18452 ( .A(n34213), .Z(n34194) );
  HS65_LH_IVX2 U18453 ( .A(n34194), .Z(n34195) );
  HS65_LH_IVX2 U18454 ( .A(n34215), .Z(n34196) );
  HS65_LH_IVX2 U18455 ( .A(n34196), .Z(n34197) );
  HS65_LH_IVX2 U18456 ( .A(n34227), .Z(n34198) );
  HS65_LH_IVX2 U18457 ( .A(n34198), .Z(n34199) );
  HS65_LH_IVX2 U18458 ( .A(n34217), .Z(n34200) );
  HS65_LH_IVX2 U18459 ( .A(n34200), .Z(n34201) );
  HS65_LH_IVX2 U18460 ( .A(n34219), .Z(n34202) );
  HS65_LH_IVX2 U18461 ( .A(n34202), .Z(n34203) );
  HS65_LH_BFX2 U18462 ( .A(n34171), .Z(n34204) );
  HS65_LH_BFX2 U18463 ( .A(n34207), .Z(n34205) );
  HS65_LH_IVX2 U18464 ( .A(n34222), .Z(n34206) );
  HS65_LH_IVX2 U18465 ( .A(n34206), .Z(n34207) );
  HS65_LH_IVX2 U18466 ( .A(n34224), .Z(n34208) );
  HS65_LH_IVX2 U18467 ( .A(n34208), .Z(n34209) );
  HS65_LH_IVX2 U18468 ( .A(n34226), .Z(n34210) );
  HS65_LH_IVX2 U18469 ( .A(n34210), .Z(n34211) );
  HS65_LH_IVX2 U18470 ( .A(n34229), .Z(n34212) );
  HS65_LH_IVX2 U18471 ( .A(n34212), .Z(n34213) );
  HS65_LH_IVX2 U18472 ( .A(n34235), .Z(n34214) );
  HS65_LH_IVX2 U18473 ( .A(n34214), .Z(n34215) );
  HS65_LH_IVX2 U18474 ( .A(n34242), .Z(n34216) );
  HS65_LH_IVX2 U18475 ( .A(n34216), .Z(n34217) );
  HS65_LH_IVX2 U18476 ( .A(n34231), .Z(n34218) );
  HS65_LH_IVX2 U18477 ( .A(n34218), .Z(n34219) );
  HS65_LH_BFX2 U18478 ( .A(n34204), .Z(n34220) );
  HS65_LH_IVX2 U18479 ( .A(n34234), .Z(n34221) );
  HS65_LH_IVX2 U18480 ( .A(n34221), .Z(n34222) );
  HS65_LH_IVX2 U18481 ( .A(n34237), .Z(n34223) );
  HS65_LH_IVX2 U18482 ( .A(n34223), .Z(n34224) );
  HS65_LH_IVX2 U18483 ( .A(n34239), .Z(n34225) );
  HS65_LH_IVX2 U18484 ( .A(n34225), .Z(n34226) );
  HS65_LH_BFX2 U18485 ( .A(n34147), .Z(n34227) );
  HS65_LH_IVX2 U18486 ( .A(n34241), .Z(n34228) );
  HS65_LH_IVX2 U18487 ( .A(n34228), .Z(n34229) );
  HS65_LH_IVX2 U18488 ( .A(n34245), .Z(n34230) );
  HS65_LH_IVX2 U18489 ( .A(n34230), .Z(n34231) );
  HS65_LH_BFX2 U18490 ( .A(n34220), .Z(n34232) );
  HS65_LH_IVX2 U18491 ( .A(n17791), .Z(n34233) );
  HS65_LH_IVX2 U18492 ( .A(n34233), .Z(n34234) );
  HS65_LH_BFX2 U18493 ( .A(n34248), .Z(n34235) );
  HS65_LH_IVX2 U18494 ( .A(n34250), .Z(n34236) );
  HS65_LH_IVX2 U18495 ( .A(n34236), .Z(n34237) );
  HS65_LH_IVX2 U18496 ( .A(n34252), .Z(n34238) );
  HS65_LH_IVX2 U18497 ( .A(n34238), .Z(n34239) );
  HS65_LH_IVX2 U18498 ( .A(n34254), .Z(n34240) );
  HS65_LH_IVX2 U18499 ( .A(n34240), .Z(n34241) );
  HS65_LH_BFX2 U18500 ( .A(n34255), .Z(n34242) );
  HS65_LH_BFX2 U18501 ( .A(n34232), .Z(n34243) );
  HS65_LH_IVX2 U18502 ( .A(n17855), .Z(n34244) );
  HS65_LH_IVX2 U18503 ( .A(n34244), .Z(n34245) );
  HS65_LH_IVX2 U18504 ( .A(n34243), .Z(n34246) );
  HS65_LH_IVX2 U18505 ( .A(n34246), .Z(n34247) );
  HS65_LH_BFX2 U18506 ( .A(n34256), .Z(n34248) );
  HS65_LH_IVX2 U18507 ( .A(n17760), .Z(n34249) );
  HS65_LH_IVX2 U18508 ( .A(n34249), .Z(n34250) );
  HS65_LH_IVX2 U18509 ( .A(n34251), .Z(n34252) );
  HS65_LH_IVX2 U18510 ( .A(n17281), .Z(n34253) );
  HS65_LH_IVX2 U18511 ( .A(n34253), .Z(n34254) );
  HS65_LH_BFX2 U18512 ( .A(n34257), .Z(n34255) );
  HS65_LH_BFX2 U18513 ( .A(n34258), .Z(n34256) );
  HS65_LH_BFX2 U18514 ( .A(n34259), .Z(n34257) );
  HS65_LH_BFX2 U18515 ( .A(n34260), .Z(n34258) );
  HS65_LH_BFX2 U18516 ( .A(n17763), .Z(n34259) );
  HS65_LH_BFX2 U18517 ( .A(n34261), .Z(n34260) );
  HS65_LH_BFX2 U18518 ( .A(n15387), .Z(n34261) );
  HS65_LH_BFX2 U18519 ( .A(n34263), .Z(n34262) );
  HS65_LH_BFX2 U18520 ( .A(n34264), .Z(n34263) );
  HS65_LH_BFX2 U18521 ( .A(n34265), .Z(n34264) );
  HS65_LH_BFX2 U18522 ( .A(n34266), .Z(n34265) );
  HS65_LH_BFX2 U18523 ( .A(n17778), .Z(n34266) );
  HS65_LH_BFX2 U18524 ( .A(n34268), .Z(n34267) );
  HS65_LH_BFX2 U18525 ( .A(n34269), .Z(n34268) );
  HS65_LH_BFX2 U18526 ( .A(n34270), .Z(n34269) );
  HS65_LH_BFX2 U18527 ( .A(n34271), .Z(n34270) );
  HS65_LH_BFX2 U18528 ( .A(n17787), .Z(n34271) );
  HS65_LH_BFX2 U18529 ( .A(n34280), .Z(n34272) );
  HS65_LH_BFX2 U18530 ( .A(n34276), .Z(n34273) );
  HS65_LH_BFX2 U18531 ( .A(n34278), .Z(n34274) );
  HS65_LH_IVX2 U18532 ( .A(n34282), .Z(n34275) );
  HS65_LH_IVX2 U18533 ( .A(n34275), .Z(n34276) );
  HS65_LH_IVX2 U18534 ( .A(n34284), .Z(n34277) );
  HS65_LH_IVX2 U18535 ( .A(n34277), .Z(n34278) );
  HS65_LH_BFX2 U18536 ( .A(n17299), .Z(n34279) );
  HS65_LH_BFX2 U18537 ( .A(n34286), .Z(n34280) );
  HS65_LH_IVX2 U18538 ( .A(n34288), .Z(n34281) );
  HS65_LH_IVX2 U18539 ( .A(n34281), .Z(n34282) );
  HS65_LH_IVX2 U18540 ( .A(n34290), .Z(n34283) );
  HS65_LH_IVX2 U18541 ( .A(n34283), .Z(n34284) );
  HS65_LH_BFX2 U18542 ( .A(n34279), .Z(n34285) );
  HS65_LH_BFX2 U18543 ( .A(n34292), .Z(n34286) );
  HS65_LH_IVX2 U18544 ( .A(n34295), .Z(n34287) );
  HS65_LH_IVX2 U18545 ( .A(n34287), .Z(n34288) );
  HS65_LH_IVX2 U18546 ( .A(n34297), .Z(n34289) );
  HS65_LH_IVX2 U18547 ( .A(n34289), .Z(n34290) );
  HS65_LH_BFX2 U18548 ( .A(n34285), .Z(n34291) );
  HS65_LH_BFX2 U18549 ( .A(n34298), .Z(n34292) );
  HS65_LH_BFX2 U18550 ( .A(n34291), .Z(n34293) );
  HS65_LH_IVX2 U18551 ( .A(n34301), .Z(n34294) );
  HS65_LH_IVX2 U18552 ( .A(n34294), .Z(n34295) );
  HS65_LH_IVX2 U18553 ( .A(n34303), .Z(n34296) );
  HS65_LH_IVX2 U18554 ( .A(n34296), .Z(n34297) );
  HS65_LH_BFX2 U18555 ( .A(n34304), .Z(n34298) );
  HS65_LH_BFX2 U18556 ( .A(n34293), .Z(n34299) );
  HS65_LH_IVX2 U18557 ( .A(n34307), .Z(n34300) );
  HS65_LH_IVX2 U18558 ( .A(n34300), .Z(n34301) );
  HS65_LH_IVX2 U18559 ( .A(n34309), .Z(n34302) );
  HS65_LH_IVX2 U18560 ( .A(n34302), .Z(n34303) );
  HS65_LH_BFX2 U18561 ( .A(n34310), .Z(n34304) );
  HS65_LH_BFX2 U18562 ( .A(n34299), .Z(n34305) );
  HS65_LH_IVX2 U18563 ( .A(n34313), .Z(n34306) );
  HS65_LH_IVX2 U18564 ( .A(n34306), .Z(n34307) );
  HS65_LH_IVX2 U18565 ( .A(n34315), .Z(n34308) );
  HS65_LH_IVX2 U18566 ( .A(n34308), .Z(n34309) );
  HS65_LH_BFX2 U18567 ( .A(n34316), .Z(n34310) );
  HS65_LH_BFX2 U18568 ( .A(n34305), .Z(n34311) );
  HS65_LH_IVX2 U18569 ( .A(n34319), .Z(n34312) );
  HS65_LH_IVX2 U18570 ( .A(n34312), .Z(n34313) );
  HS65_LH_IVX2 U18571 ( .A(n34321), .Z(n34314) );
  HS65_LH_IVX2 U18572 ( .A(n34314), .Z(n34315) );
  HS65_LH_BFX2 U18573 ( .A(n34322), .Z(n34316) );
  HS65_LH_BFX2 U18574 ( .A(n34311), .Z(n34317) );
  HS65_LH_IVX2 U18575 ( .A(n34325), .Z(n34318) );
  HS65_LH_IVX2 U18576 ( .A(n34318), .Z(n34319) );
  HS65_LH_IVX2 U18577 ( .A(n34327), .Z(n34320) );
  HS65_LH_IVX2 U18578 ( .A(n34320), .Z(n34321) );
  HS65_LH_BFX2 U18579 ( .A(n34328), .Z(n34322) );
  HS65_LH_BFX2 U18580 ( .A(n34317), .Z(n34323) );
  HS65_LH_IVX2 U18581 ( .A(n34331), .Z(n34324) );
  HS65_LH_IVX2 U18582 ( .A(n34324), .Z(n34325) );
  HS65_LH_IVX2 U18583 ( .A(n34333), .Z(n34326) );
  HS65_LH_IVX2 U18584 ( .A(n34326), .Z(n34327) );
  HS65_LH_BFX2 U18585 ( .A(n34334), .Z(n34328) );
  HS65_LH_BFX2 U18586 ( .A(n34323), .Z(n34329) );
  HS65_LH_IVX2 U18587 ( .A(n34337), .Z(n34330) );
  HS65_LH_IVX2 U18588 ( .A(n34330), .Z(n34331) );
  HS65_LH_IVX2 U18589 ( .A(n34339), .Z(n34332) );
  HS65_LH_IVX2 U18590 ( .A(n34332), .Z(n34333) );
  HS65_LH_BFX2 U18591 ( .A(n34340), .Z(n34334) );
  HS65_LH_BFX2 U18592 ( .A(n34329), .Z(n34335) );
  HS65_LH_IVX2 U18593 ( .A(n34346), .Z(n34336) );
  HS65_LH_IVX2 U18594 ( .A(n34336), .Z(n34337) );
  HS65_LH_IVX2 U18595 ( .A(n34344), .Z(n34338) );
  HS65_LH_IVX2 U18596 ( .A(n34338), .Z(n34339) );
  HS65_LH_BFX2 U18597 ( .A(n34342), .Z(n34340) );
  HS65_LH_BFX2 U18598 ( .A(n34335), .Z(n34341) );
  HS65_LH_BFX2 U18599 ( .A(n34347), .Z(n34342) );
  HS65_LH_IVX2 U18600 ( .A(n34349), .Z(n34343) );
  HS65_LH_IVX2 U18601 ( .A(n34343), .Z(n34344) );
  HS65_LH_BFX2 U18602 ( .A(n34341), .Z(n34345) );
  HS65_LH_BFX2 U18603 ( .A(n34352), .Z(n34346) );
  HS65_LH_BFX2 U18604 ( .A(n34351), .Z(n34347) );
  HS65_LH_IVX2 U18605 ( .A(n34358), .Z(n34348) );
  HS65_LH_IVX2 U18606 ( .A(n34348), .Z(n34349) );
  HS65_LH_BFX2 U18607 ( .A(n34345), .Z(n34350) );
  HS65_LH_BFX2 U18608 ( .A(n34356), .Z(n34351) );
  HS65_LH_BFX2 U18609 ( .A(n34354), .Z(n34352) );
  HS65_LH_IVX2 U18610 ( .A(n34363), .Z(n34353) );
  HS65_LH_IVX2 U18611 ( .A(n34353), .Z(n34354) );
  HS65_LH_IVX2 U18612 ( .A(n17692), .Z(n34355) );
  HS65_LH_IVX2 U18613 ( .A(n34355), .Z(n34356) );
  HS65_LH_IVX2 U18614 ( .A(n34361), .Z(n34357) );
  HS65_LH_IVX2 U18615 ( .A(n34357), .Z(n34358) );
  HS65_LH_BFX2 U18616 ( .A(n34350), .Z(n34359) );
  HS65_LH_IVX2 U18617 ( .A(n34366), .Z(n34360) );
  HS65_LH_IVX2 U18618 ( .A(n34360), .Z(n34361) );
  HS65_LH_BFX2 U18619 ( .A(n34359), .Z(n34362) );
  HS65_LH_BFX2 U18620 ( .A(n34365), .Z(n34363) );
  HS65_LH_BFX2 U18621 ( .A(n34362), .Z(n34364) );
  HS65_LH_BFX2 U18622 ( .A(n34370), .Z(n34365) );
  HS65_LH_BFX2 U18623 ( .A(n34371), .Z(n34366) );
  HS65_LH_BFX2 U18624 ( .A(n34364), .Z(n34367) );
  HS65_LH_IVX2 U18625 ( .A(n34367), .Z(n34368) );
  HS65_LH_IVX2 U18626 ( .A(n34368), .Z(n34369) );
  HS65_LH_BFX2 U18627 ( .A(n17294), .Z(n34370) );
  HS65_LH_BFX2 U18628 ( .A(n17435), .Z(n34371) );
  HS65_LH_BFX2 U18629 ( .A(n34373), .Z(n34372) );
  HS65_LH_BFX2 U18630 ( .A(n34374), .Z(n34373) );
  HS65_LH_BFX2 U18631 ( .A(n34375), .Z(n34374) );
  HS65_LH_BFX2 U18632 ( .A(n34376), .Z(n34375) );
  HS65_LH_BFX2 U18633 ( .A(n17772), .Z(n34376) );
  HS65_LH_BFX2 U18634 ( .A(n34379), .Z(n34377) );
  HS65_LH_BFX2 U18635 ( .A(n34380), .Z(n34378) );
  HS65_LH_BFX2 U18636 ( .A(n34381), .Z(n34379) );
  HS65_LH_BFX2 U18637 ( .A(n34382), .Z(n34380) );
  HS65_LH_BFX2 U18638 ( .A(n34383), .Z(n34381) );
  HS65_LH_BFX2 U18639 ( .A(n34384), .Z(n34382) );
  HS65_LH_BFX2 U18640 ( .A(n34385), .Z(n34383) );
  HS65_LH_BFX2 U18641 ( .A(n34386), .Z(n34384) );
  HS65_LH_BFX2 U18642 ( .A(n17768), .Z(n34385) );
  HS65_LH_BFX2 U18643 ( .A(n17769), .Z(n34386) );
  HS65_LH_BFX2 U18644 ( .A(n34388), .Z(n34387) );
  HS65_LH_BFX2 U18645 ( .A(n34389), .Z(n34388) );
  HS65_LH_BFX2 U18646 ( .A(n34390), .Z(n34389) );
  HS65_LH_BFX2 U18647 ( .A(n34391), .Z(n34390) );
  HS65_LH_BFX2 U18648 ( .A(n17582), .Z(n34391) );
  HS65_LH_BFX2 U18649 ( .A(n34394), .Z(n34392) );
  HS65_LH_IVX2 U18650 ( .A(n34398), .Z(n34393) );
  HS65_LH_IVX2 U18651 ( .A(n34393), .Z(n34394) );
  HS65_LH_BFX2 U18652 ( .A(n34396), .Z(n34395) );
  HS65_LH_BFX2 U18653 ( .A(n34399), .Z(n34396) );
  HS65_LH_BFX2 U18654 ( .A(n34400), .Z(n34397) );
  HS65_LH_BFX2 U18655 ( .A(n34401), .Z(n34398) );
  HS65_LH_BFX2 U18656 ( .A(n34402), .Z(n34399) );
  HS65_LH_BFX2 U18657 ( .A(n34403), .Z(n34400) );
  HS65_LH_BFX2 U18658 ( .A(n34404), .Z(n34401) );
  HS65_LH_BFX2 U18659 ( .A(n34405), .Z(n34402) );
  HS65_LH_BFX2 U18660 ( .A(n34406), .Z(n34403) );
  HS65_LH_BFX2 U18661 ( .A(n34407), .Z(n34404) );
  HS65_LH_BFX2 U18662 ( .A(n34408), .Z(n34405) );
  HS65_LH_BFX2 U18663 ( .A(n34409), .Z(n34406) );
  HS65_LH_BFX2 U18664 ( .A(n34410), .Z(n34407) );
  HS65_LH_BFX2 U18665 ( .A(n34411), .Z(n34408) );
  HS65_LH_BFX2 U18666 ( .A(n34412), .Z(n34409) );
  HS65_LH_BFX2 U18667 ( .A(n34413), .Z(n34410) );
  HS65_LH_BFX2 U18668 ( .A(n34414), .Z(n34411) );
  HS65_LH_BFX2 U18669 ( .A(n34415), .Z(n34412) );
  HS65_LH_BFX2 U18670 ( .A(n34416), .Z(n34413) );
  HS65_LH_BFX2 U18671 ( .A(n34417), .Z(n34414) );
  HS65_LH_BFX2 U18672 ( .A(n34418), .Z(n34415) );
  HS65_LH_BFX2 U18673 ( .A(n34419), .Z(n34416) );
  HS65_LH_BFX2 U18674 ( .A(n34420), .Z(n34417) );
  HS65_LH_BFX2 U18675 ( .A(n34421), .Z(n34418) );
  HS65_LH_BFX2 U18676 ( .A(n1896), .Z(n34419) );
  HS65_LH_BFX2 U18677 ( .A(n1897), .Z(n34420) );
  HS65_LH_BFX2 U18678 ( .A(n34422), .Z(n34421) );
  HS65_LH_BFX2 U18679 ( .A(n34423), .Z(n34422) );
  HS65_LH_BFX2 U18680 ( .A(n34424), .Z(n34423) );
  HS65_LH_BFX2 U18681 ( .A(n17861), .Z(n34424) );
  HS65_LH_BFX2 U18682 ( .A(n34426), .Z(n34425) );
  HS65_LH_BFX2 U18683 ( .A(n34427), .Z(n34426) );
  HS65_LH_BFX2 U18684 ( .A(n34428), .Z(n34427) );
  HS65_LH_BFX2 U18685 ( .A(n34429), .Z(n34428) );
  HS65_LH_BFX2 U18686 ( .A(n34430), .Z(n34429) );
  HS65_LH_BFX2 U18687 ( .A(n17789), .Z(n34430) );
  HS65_LH_BFX2 U18688 ( .A(n34434), .Z(n34431) );
  HS65_LH_BFX2 U18689 ( .A(n34438), .Z(n34432) );
  HS65_LH_IVX2 U18690 ( .A(n34447), .Z(n34433) );
  HS65_LH_IVX2 U18691 ( .A(n34433), .Z(n34434) );
  HS65_LH_BFX2 U18692 ( .A(n34440), .Z(n34435) );
  HS65_LH_BFX2 U18693 ( .A(n34443), .Z(n34436) );
  HS65_LH_IVX2 U18694 ( .A(n34449), .Z(n34437) );
  HS65_LH_IVX2 U18695 ( .A(n34437), .Z(n34438) );
  HS65_LH_IVX2 U18696 ( .A(n34451), .Z(n34439) );
  HS65_LH_IVX2 U18697 ( .A(n34439), .Z(n34440) );
  HS65_LH_BFX2 U18698 ( .A(n34445), .Z(n34441) );
  HS65_LH_IVX2 U18699 ( .A(n34453), .Z(n34442) );
  HS65_LH_IVX2 U18700 ( .A(n34442), .Z(n34443) );
  HS65_LH_IVX2 U18701 ( .A(n34455), .Z(n34444) );
  HS65_LH_IVX2 U18702 ( .A(n34444), .Z(n34445) );
  HS65_LH_IVX2 U18703 ( .A(n34457), .Z(n34446) );
  HS65_LH_IVX2 U18704 ( .A(n34446), .Z(n34447) );
  HS65_LH_IVX2 U18705 ( .A(n34459), .Z(n34448) );
  HS65_LH_IVX2 U18706 ( .A(n34448), .Z(n34449) );
  HS65_LH_IVX2 U18707 ( .A(n34461), .Z(n34450) );
  HS65_LH_IVX2 U18708 ( .A(n34450), .Z(n34451) );
  HS65_LH_IVX2 U18709 ( .A(n34463), .Z(n34452) );
  HS65_LH_IVX2 U18710 ( .A(n34452), .Z(n34453) );
  HS65_LH_IVX2 U18711 ( .A(n34465), .Z(n34454) );
  HS65_LH_IVX2 U18712 ( .A(n34454), .Z(n34455) );
  HS65_LH_IVX2 U18713 ( .A(n34474), .Z(n34456) );
  HS65_LH_IVX2 U18714 ( .A(n34456), .Z(n34457) );
  HS65_LH_IVX2 U18715 ( .A(n34467), .Z(n34458) );
  HS65_LH_IVX2 U18716 ( .A(n34458), .Z(n34459) );
  HS65_LH_IVX2 U18717 ( .A(n34469), .Z(n34460) );
  HS65_LH_IVX2 U18718 ( .A(n34460), .Z(n34461) );
  HS65_LH_IVX2 U18719 ( .A(n34471), .Z(n34462) );
  HS65_LH_IVX2 U18720 ( .A(n34462), .Z(n34463) );
  HS65_LH_IVX2 U18721 ( .A(n34473), .Z(n34464) );
  HS65_LH_IVX2 U18722 ( .A(n34464), .Z(n34465) );
  HS65_LH_IVX2 U18723 ( .A(n34476), .Z(n34466) );
  HS65_LH_IVX2 U18724 ( .A(n34466), .Z(n34467) );
  HS65_LH_IVX2 U18725 ( .A(n34478), .Z(n34468) );
  HS65_LH_IVX2 U18726 ( .A(n34468), .Z(n34469) );
  HS65_LH_IVX2 U18727 ( .A(n34480), .Z(n34470) );
  HS65_LH_IVX2 U18728 ( .A(n34470), .Z(n34471) );
  HS65_LH_IVX2 U18729 ( .A(n34482), .Z(n34472) );
  HS65_LH_IVX2 U18730 ( .A(n34472), .Z(n34473) );
  HS65_LH_BFX2 U18731 ( .A(n34483), .Z(n34474) );
  HS65_LH_IVX2 U18732 ( .A(n34485), .Z(n34475) );
  HS65_LH_IVX2 U18733 ( .A(n34475), .Z(n34476) );
  HS65_LH_IVX2 U18734 ( .A(n34487), .Z(n34477) );
  HS65_LH_IVX2 U18735 ( .A(n34477), .Z(n34478) );
  HS65_LH_IVX2 U18736 ( .A(n34489), .Z(n34479) );
  HS65_LH_IVX2 U18737 ( .A(n34479), .Z(n34480) );
  HS65_LH_IVX2 U18738 ( .A(n34491), .Z(n34481) );
  HS65_LH_IVX2 U18739 ( .A(n34481), .Z(n34482) );
  HS65_LH_BFX2 U18740 ( .A(n34492), .Z(n34483) );
  HS65_LH_IVX2 U18741 ( .A(n34494), .Z(n34484) );
  HS65_LH_IVX2 U18742 ( .A(n34484), .Z(n34485) );
  HS65_LH_IVX2 U18743 ( .A(n34496), .Z(n34486) );
  HS65_LH_IVX2 U18744 ( .A(n34486), .Z(n34487) );
  HS65_LH_IVX2 U18745 ( .A(n34498), .Z(n34488) );
  HS65_LH_IVX2 U18746 ( .A(n34488), .Z(n34489) );
  HS65_LH_IVX2 U18747 ( .A(n34500), .Z(n34490) );
  HS65_LH_IVX2 U18748 ( .A(n34490), .Z(n34491) );
  HS65_LH_BFX2 U18749 ( .A(n34501), .Z(n34492) );
  HS65_LH_IVX2 U18750 ( .A(n34503), .Z(n34493) );
  HS65_LH_IVX2 U18751 ( .A(n34493), .Z(n34494) );
  HS65_LH_IVX2 U18752 ( .A(n34505), .Z(n34495) );
  HS65_LH_IVX2 U18753 ( .A(n34495), .Z(n34496) );
  HS65_LH_IVX2 U18754 ( .A(n34507), .Z(n34497) );
  HS65_LH_IVX2 U18755 ( .A(n34497), .Z(n34498) );
  HS65_LH_IVX2 U18756 ( .A(n34509), .Z(n34499) );
  HS65_LH_IVX2 U18757 ( .A(n34499), .Z(n34500) );
  HS65_LH_BFX2 U18758 ( .A(n34510), .Z(n34501) );
  HS65_LH_IVX2 U18759 ( .A(n34512), .Z(n34502) );
  HS65_LH_IVX2 U18760 ( .A(n34502), .Z(n34503) );
  HS65_LH_IVX2 U18761 ( .A(n34514), .Z(n34504) );
  HS65_LH_IVX2 U18762 ( .A(n34504), .Z(n34505) );
  HS65_LH_IVX2 U18763 ( .A(n34516), .Z(n34506) );
  HS65_LH_IVX2 U18764 ( .A(n34506), .Z(n34507) );
  HS65_LH_IVX2 U18765 ( .A(n34518), .Z(n34508) );
  HS65_LH_IVX2 U18766 ( .A(n34508), .Z(n34509) );
  HS65_LH_BFX2 U18767 ( .A(n34519), .Z(n34510) );
  HS65_LH_IVX2 U18768 ( .A(n34521), .Z(n34511) );
  HS65_LH_IVX2 U18769 ( .A(n34511), .Z(n34512) );
  HS65_LH_IVX2 U18770 ( .A(n34523), .Z(n34513) );
  HS65_LH_IVX2 U18771 ( .A(n34513), .Z(n34514) );
  HS65_LH_IVX2 U18772 ( .A(n34525), .Z(n34515) );
  HS65_LH_IVX2 U18773 ( .A(n34515), .Z(n34516) );
  HS65_LH_IVX2 U18774 ( .A(n34527), .Z(n34517) );
  HS65_LH_IVX2 U18775 ( .A(n34517), .Z(n34518) );
  HS65_LH_BFX2 U18776 ( .A(n35564), .Z(n34519) );
  HS65_LH_IVX2 U18777 ( .A(n34529), .Z(n34520) );
  HS65_LH_IVX2 U18778 ( .A(n34520), .Z(n34521) );
  HS65_LH_IVX2 U18779 ( .A(n34531), .Z(n34522) );
  HS65_LH_IVX2 U18780 ( .A(n34522), .Z(n34523) );
  HS65_LH_IVX2 U18781 ( .A(n34533), .Z(n34524) );
  HS65_LH_IVX2 U18782 ( .A(n34524), .Z(n34525) );
  HS65_LH_IVX2 U18783 ( .A(n34535), .Z(n34526) );
  HS65_LH_IVX2 U18784 ( .A(n34526), .Z(n34527) );
  HS65_LH_IVX2 U18785 ( .A(n34537), .Z(n34528) );
  HS65_LH_IVX2 U18786 ( .A(n34528), .Z(n34529) );
  HS65_LH_IVX2 U18787 ( .A(n34539), .Z(n34530) );
  HS65_LH_IVX2 U18788 ( .A(n34530), .Z(n34531) );
  HS65_LH_IVX2 U18789 ( .A(n34541), .Z(n34532) );
  HS65_LH_IVX2 U18790 ( .A(n34532), .Z(n34533) );
  HS65_LH_IVX2 U18791 ( .A(n34543), .Z(n34534) );
  HS65_LH_IVX2 U18792 ( .A(n34534), .Z(n34535) );
  HS65_LH_IVX2 U18793 ( .A(n34545), .Z(n34536) );
  HS65_LH_IVX2 U18794 ( .A(n34536), .Z(n34537) );
  HS65_LH_IVX2 U18795 ( .A(n34547), .Z(n34538) );
  HS65_LH_IVX2 U18796 ( .A(n34538), .Z(n34539) );
  HS65_LH_IVX2 U18797 ( .A(n34549), .Z(n34540) );
  HS65_LH_IVX2 U18798 ( .A(n34540), .Z(n34541) );
  HS65_LH_IVX2 U18799 ( .A(n34551), .Z(n34542) );
  HS65_LH_IVX2 U18800 ( .A(n34542), .Z(n34543) );
  HS65_LH_IVX2 U18801 ( .A(n34553), .Z(n34544) );
  HS65_LH_IVX2 U18802 ( .A(n34544), .Z(n34545) );
  HS65_LH_IVX2 U18803 ( .A(n34555), .Z(n34546) );
  HS65_LH_IVX2 U18804 ( .A(n34546), .Z(n34547) );
  HS65_LH_IVX2 U18805 ( .A(n34557), .Z(n34548) );
  HS65_LH_IVX2 U18806 ( .A(n34548), .Z(n34549) );
  HS65_LH_IVX2 U18807 ( .A(n34559), .Z(n34550) );
  HS65_LH_IVX2 U18808 ( .A(n34550), .Z(n34551) );
  HS65_LH_IVX2 U18809 ( .A(n34561), .Z(n34552) );
  HS65_LH_IVX2 U18810 ( .A(n34552), .Z(n34553) );
  HS65_LH_IVX2 U18811 ( .A(n34563), .Z(n34554) );
  HS65_LH_IVX2 U18812 ( .A(n34554), .Z(n34555) );
  HS65_LH_IVX2 U18813 ( .A(n34565), .Z(n34556) );
  HS65_LH_IVX2 U18814 ( .A(n34556), .Z(n34557) );
  HS65_LH_IVX2 U18815 ( .A(n34567), .Z(n34558) );
  HS65_LH_IVX2 U18816 ( .A(n34558), .Z(n34559) );
  HS65_LH_IVX2 U18817 ( .A(n34569), .Z(n34560) );
  HS65_LH_IVX2 U18818 ( .A(n34560), .Z(n34561) );
  HS65_LH_IVX2 U18819 ( .A(n34571), .Z(n34562) );
  HS65_LH_IVX2 U18820 ( .A(n34562), .Z(n34563) );
  HS65_LH_IVX2 U18821 ( .A(n34573), .Z(n34564) );
  HS65_LH_IVX2 U18822 ( .A(n34564), .Z(n34565) );
  HS65_LH_IVX2 U18823 ( .A(n34575), .Z(n34566) );
  HS65_LH_IVX2 U18824 ( .A(n34566), .Z(n34567) );
  HS65_LH_IVX2 U18825 ( .A(n34578), .Z(n34568) );
  HS65_LH_IVX2 U18826 ( .A(n34568), .Z(n34569) );
  HS65_LH_IVX2 U18827 ( .A(n17298), .Z(n34570) );
  HS65_LH_IVX2 U18828 ( .A(n34570), .Z(n34571) );
  HS65_LH_IVX2 U18829 ( .A(n34577), .Z(n34572) );
  HS65_LH_IVX2 U18830 ( .A(n34572), .Z(n34573) );
  HS65_LH_IVX2 U18831 ( .A(n17570), .Z(n34574) );
  HS65_LH_IVX2 U18832 ( .A(n34574), .Z(n34575) );
  HS65_LH_IVX2 U18833 ( .A(n17438), .Z(n34576) );
  HS65_LH_IVX2 U18834 ( .A(n34576), .Z(n34577) );
  HS65_LH_BFX2 U18835 ( .A(n17439), .Z(n34578) );
  HS65_LH_BFX2 U18836 ( .A(n34585), .Z(n34579) );
  HS65_LH_BFX2 U18837 ( .A(n34583), .Z(n34580) );
  HS65_LH_BFX2 U18838 ( .A(n17295), .Z(n34581) );
  HS65_LH_IVX2 U18839 ( .A(n34588), .Z(n34582) );
  HS65_LH_IVX2 U18840 ( .A(n34582), .Z(n34583) );
  HS65_LH_BFX2 U18841 ( .A(n17513), .Z(n34584) );
  HS65_LH_BFX2 U18842 ( .A(n34590), .Z(n34585) );
  HS65_LH_BFX2 U18843 ( .A(n34581), .Z(n34586) );
  HS65_LH_IVX2 U18844 ( .A(n34594), .Z(n34587) );
  HS65_LH_IVX2 U18845 ( .A(n34587), .Z(n34588) );
  HS65_LH_BFX2 U18846 ( .A(n34584), .Z(n34589) );
  HS65_LH_BFX2 U18847 ( .A(n34597), .Z(n34590) );
  HS65_LH_BFX2 U18848 ( .A(n34586), .Z(n34591) );
  HS65_LH_BFX2 U18849 ( .A(n34589), .Z(n34592) );
  HS65_LH_IVX2 U18850 ( .A(n34600), .Z(n34593) );
  HS65_LH_IVX2 U18851 ( .A(n34593), .Z(n34594) );
  HS65_LH_IVX2 U18852 ( .A(n34602), .Z(n34595) );
  HS65_LH_IVX2 U18853 ( .A(n34595), .Z(n34596) );
  HS65_LH_BFX2 U18854 ( .A(n34603), .Z(n34597) );
  HS65_LH_BFX2 U18855 ( .A(n34591), .Z(n34598) );
  HS65_LH_IVX2 U18856 ( .A(n34606), .Z(n34599) );
  HS65_LH_IVX2 U18857 ( .A(n34599), .Z(n34600) );
  HS65_LH_IVX2 U18858 ( .A(n34608), .Z(n34601) );
  HS65_LH_IVX2 U18859 ( .A(n34601), .Z(n34602) );
  HS65_LH_BFX2 U18860 ( .A(n34609), .Z(n34603) );
  HS65_LH_BFX2 U18861 ( .A(n34598), .Z(n34604) );
  HS65_LH_IVX2 U18862 ( .A(n34612), .Z(n34605) );
  HS65_LH_IVX2 U18863 ( .A(n34605), .Z(n34606) );
  HS65_LH_IVX2 U18864 ( .A(n34614), .Z(n34607) );
  HS65_LH_IVX2 U18865 ( .A(n34607), .Z(n34608) );
  HS65_LH_BFX2 U18866 ( .A(n34615), .Z(n34609) );
  HS65_LH_BFX2 U18867 ( .A(n34604), .Z(n34610) );
  HS65_LH_IVX2 U18868 ( .A(n34618), .Z(n34611) );
  HS65_LH_IVX2 U18869 ( .A(n34611), .Z(n34612) );
  HS65_LH_IVX2 U18870 ( .A(n34620), .Z(n34613) );
  HS65_LH_IVX2 U18871 ( .A(n34613), .Z(n34614) );
  HS65_LH_BFX2 U18872 ( .A(n34621), .Z(n34615) );
  HS65_LH_BFX2 U18873 ( .A(n34610), .Z(n34616) );
  HS65_LH_IVX2 U18874 ( .A(n34624), .Z(n34617) );
  HS65_LH_IVX2 U18875 ( .A(n34617), .Z(n34618) );
  HS65_LH_IVX2 U18876 ( .A(n34626), .Z(n34619) );
  HS65_LH_IVX2 U18877 ( .A(n34619), .Z(n34620) );
  HS65_LH_BFX2 U18878 ( .A(n34627), .Z(n34621) );
  HS65_LH_BFX2 U18879 ( .A(n34616), .Z(n34622) );
  HS65_LH_IVX2 U18880 ( .A(n34630), .Z(n34623) );
  HS65_LH_IVX2 U18881 ( .A(n34623), .Z(n34624) );
  HS65_LH_IVX2 U18882 ( .A(n34632), .Z(n34625) );
  HS65_LH_IVX2 U18883 ( .A(n34625), .Z(n34626) );
  HS65_LH_BFX2 U18884 ( .A(n34633), .Z(n34627) );
  HS65_LH_BFX2 U18885 ( .A(n34622), .Z(n34628) );
  HS65_LH_IVX2 U18886 ( .A(n34636), .Z(n34629) );
  HS65_LH_IVX2 U18887 ( .A(n34629), .Z(n34630) );
  HS65_LH_IVX2 U18888 ( .A(n34638), .Z(n34631) );
  HS65_LH_IVX2 U18889 ( .A(n34631), .Z(n34632) );
  HS65_LH_BFX2 U18890 ( .A(n34639), .Z(n34633) );
  HS65_LH_BFX2 U18891 ( .A(n34628), .Z(n34634) );
  HS65_LH_IVX2 U18892 ( .A(n34645), .Z(n34635) );
  HS65_LH_IVX2 U18893 ( .A(n34635), .Z(n34636) );
  HS65_LH_IVX2 U18894 ( .A(n34643), .Z(n34637) );
  HS65_LH_IVX2 U18895 ( .A(n34637), .Z(n34638) );
  HS65_LH_BFX2 U18896 ( .A(n34641), .Z(n34639) );
  HS65_LH_BFX2 U18897 ( .A(n34634), .Z(n34640) );
  HS65_LH_BFX2 U18898 ( .A(n34646), .Z(n34641) );
  HS65_LH_IVX2 U18899 ( .A(n34664), .Z(n34642) );
  HS65_LH_IVX2 U18900 ( .A(n34642), .Z(n34643) );
  HS65_LH_BFX2 U18901 ( .A(n34640), .Z(n34644) );
  HS65_LH_BFX2 U18902 ( .A(n34648), .Z(n34645) );
  HS65_LH_BFX2 U18903 ( .A(n34650), .Z(n34646) );
  HS65_LH_IVX2 U18904 ( .A(n34653), .Z(n34647) );
  HS65_LH_IVX2 U18905 ( .A(n34647), .Z(n34648) );
  HS65_LH_BFX2 U18906 ( .A(n34644), .Z(n34649) );
  HS65_LH_BFX2 U18907 ( .A(n34655), .Z(n34650) );
  HS65_LH_BFX2 U18908 ( .A(n34592), .Z(n34651) );
  HS65_LH_IVX2 U18909 ( .A(n34659), .Z(n34652) );
  HS65_LH_IVX2 U18910 ( .A(n34652), .Z(n34653) );
  HS65_LH_BFX2 U18911 ( .A(n34649), .Z(n34654) );
  HS65_LH_BFX2 U18912 ( .A(n34660), .Z(n34655) );
  HS65_LH_BFX2 U18913 ( .A(n34651), .Z(n34656) );
  HS65_LH_BFX2 U18914 ( .A(n34654), .Z(n34657) );
  HS65_LH_IVX2 U18915 ( .A(n34666), .Z(n34658) );
  HS65_LH_IVX2 U18916 ( .A(n34658), .Z(n34659) );
  HS65_LH_BFX2 U18917 ( .A(n34667), .Z(n34660) );
  HS65_LH_BFX2 U18918 ( .A(n34656), .Z(n34661) );
  HS65_LH_BFX2 U18919 ( .A(n34657), .Z(n34662) );
  HS65_LH_IVX2 U18920 ( .A(n34672), .Z(n34663) );
  HS65_LH_IVX2 U18921 ( .A(n34663), .Z(n34664) );
  HS65_LH_IVX2 U18922 ( .A(n34674), .Z(n34665) );
  HS65_LH_IVX2 U18923 ( .A(n34665), .Z(n34666) );
  HS65_LH_BFX2 U18924 ( .A(n34675), .Z(n34667) );
  HS65_LH_BFX2 U18925 ( .A(n34662), .Z(n34668) );
  HS65_LH_IVX2 U18926 ( .A(n34680), .Z(n34669) );
  HS65_LH_IVX2 U18927 ( .A(n34669), .Z(n34670) );
  HS65_LH_IVX2 U18928 ( .A(n34677), .Z(n34671) );
  HS65_LH_IVX2 U18929 ( .A(n34671), .Z(n34672) );
  HS65_LH_IVX2 U18930 ( .A(n34679), .Z(n34673) );
  HS65_LH_IVX2 U18931 ( .A(n34673), .Z(n34674) );
  HS65_LH_BFX2 U18932 ( .A(n34681), .Z(n34675) );
  HS65_LH_IVX2 U18933 ( .A(n34661), .Z(n34676) );
  HS65_LH_IVX2 U18934 ( .A(n34676), .Z(n34677) );
  HS65_LH_IVX2 U18935 ( .A(n29540), .Z(n34678) );
  HS65_LH_IVX2 U18936 ( .A(n34678), .Z(n34679) );
  HS65_LH_BFX2 U18937 ( .A(n34682), .Z(n34680) );
  HS65_LH_BFX2 U18938 ( .A(n29766), .Z(n34681) );
  HS65_LH_BFX2 U18939 ( .A(n34683), .Z(n34682) );
  HS65_LH_BFX2 U18940 ( .A(n34668), .Z(n34683) );
  HS65_LH_BFX2 U18941 ( .A(n34715), .Z(n34684) );
  HS65_LH_OAI112X1 U18942 ( .A(n34687), .B(n34693), .C(n34702), .D(n34713), 
        .Z(n213) );
  HS65_LH_BFX2 U18943 ( .A(n17640), .Z(n34685) );
  HS65_LH_BFX2 U18944 ( .A(n34692), .Z(n34686) );
  HS65_LH_BFX2 U18945 ( .A(n34695), .Z(n34687) );
  HS65_LH_BFX2 U18946 ( .A(n34697), .Z(n34688) );
  HS65_LH_IVX2 U18947 ( .A(n34719), .Z(n34689) );
  HS65_LH_IVX2 U18948 ( .A(n34689), .Z(n34690) );
  HS65_LH_IVX2 U18949 ( .A(n34721), .Z(n34691) );
  HS65_LH_IVX2 U18950 ( .A(n34691), .Z(n34692) );
  HS65_LH_BFX2 U18951 ( .A(n34699), .Z(n34693) );
  HS65_LH_IVX2 U18952 ( .A(n34723), .Z(n34694) );
  HS65_LH_IVX2 U18953 ( .A(n34694), .Z(n34695) );
  HS65_LH_IVX2 U18954 ( .A(n34725), .Z(n34696) );
  HS65_LH_IVX2 U18955 ( .A(n34696), .Z(n34697) );
  HS65_LH_IVX2 U18956 ( .A(n34727), .Z(n34698) );
  HS65_LH_IVX2 U18957 ( .A(n34698), .Z(n34699) );
  HS65_LH_BFX2 U18958 ( .A(n34705), .Z(n34700) );
  HS65_LH_BFX2 U18959 ( .A(n34707), .Z(n34701) );
  HS65_LH_BFX2 U18960 ( .A(n34709), .Z(n34702) );
  HS65_LH_BFX2 U18961 ( .A(n34711), .Z(n34703) );
  HS65_LH_IVX2 U18962 ( .A(n34729), .Z(n34704) );
  HS65_LH_IVX2 U18963 ( .A(n34704), .Z(n34705) );
  HS65_LH_IVX2 U18964 ( .A(n34731), .Z(n34706) );
  HS65_LH_IVX2 U18965 ( .A(n34706), .Z(n34707) );
  HS65_LH_IVX2 U18966 ( .A(n34733), .Z(n34708) );
  HS65_LH_IVX2 U18967 ( .A(n34708), .Z(n34709) );
  HS65_LH_IVX2 U18968 ( .A(n34735), .Z(n34710) );
  HS65_LH_IVX2 U18969 ( .A(n34710), .Z(n34711) );
  HS65_LH_BFX2 U18970 ( .A(n17437), .Z(n34712) );
  HS65_LH_BFX2 U18971 ( .A(n34717), .Z(n34713) );
  HS65_LH_IVX2 U18972 ( .A(n34737), .Z(n34714) );
  HS65_LH_IVX2 U18973 ( .A(n34714), .Z(n34715) );
  HS65_LH_IVX2 U18974 ( .A(n34739), .Z(n34716) );
  HS65_LH_IVX2 U18975 ( .A(n34716), .Z(n34717) );
  HS65_LH_IVX2 U18976 ( .A(n34741), .Z(n34718) );
  HS65_LH_IVX2 U18977 ( .A(n34718), .Z(n34719) );
  HS65_LH_IVX2 U18978 ( .A(n34743), .Z(n34720) );
  HS65_LH_IVX2 U18979 ( .A(n34720), .Z(n34721) );
  HS65_LH_IVX2 U18980 ( .A(n34745), .Z(n34722) );
  HS65_LH_IVX2 U18981 ( .A(n34722), .Z(n34723) );
  HS65_LH_IVX2 U18982 ( .A(n34747), .Z(n34724) );
  HS65_LH_IVX2 U18983 ( .A(n34724), .Z(n34725) );
  HS65_LH_IVX2 U18984 ( .A(n34749), .Z(n34726) );
  HS65_LH_IVX2 U18985 ( .A(n34726), .Z(n34727) );
  HS65_LH_IVX2 U18986 ( .A(n34751), .Z(n34728) );
  HS65_LH_IVX2 U18987 ( .A(n34728), .Z(n34729) );
  HS65_LH_IVX2 U18988 ( .A(n34753), .Z(n34730) );
  HS65_LH_IVX2 U18989 ( .A(n34730), .Z(n34731) );
  HS65_LH_IVX2 U18990 ( .A(n34755), .Z(n34732) );
  HS65_LH_IVX2 U18991 ( .A(n34732), .Z(n34733) );
  HS65_LH_IVX2 U18992 ( .A(n34757), .Z(n34734) );
  HS65_LH_IVX2 U18993 ( .A(n34734), .Z(n34735) );
  HS65_LH_IVX2 U18994 ( .A(n34759), .Z(n34736) );
  HS65_LH_IVX2 U18995 ( .A(n34736), .Z(n34737) );
  HS65_LH_IVX2 U18996 ( .A(n34761), .Z(n34738) );
  HS65_LH_IVX2 U18997 ( .A(n34738), .Z(n34739) );
  HS65_LH_IVX2 U18998 ( .A(n34763), .Z(n34740) );
  HS65_LH_IVX2 U18999 ( .A(n34740), .Z(n34741) );
  HS65_LH_IVX2 U19000 ( .A(n34765), .Z(n34742) );
  HS65_LH_IVX2 U19001 ( .A(n34742), .Z(n34743) );
  HS65_LH_IVX2 U19002 ( .A(n34767), .Z(n34744) );
  HS65_LH_IVX2 U19003 ( .A(n34744), .Z(n34745) );
  HS65_LH_IVX2 U19004 ( .A(n34769), .Z(n34746) );
  HS65_LH_IVX2 U19005 ( .A(n34746), .Z(n34747) );
  HS65_LH_IVX2 U19006 ( .A(n34771), .Z(n34748) );
  HS65_LH_IVX2 U19007 ( .A(n34748), .Z(n34749) );
  HS65_LH_IVX2 U19008 ( .A(n34773), .Z(n34750) );
  HS65_LH_IVX2 U19009 ( .A(n34750), .Z(n34751) );
  HS65_LH_IVX2 U19010 ( .A(n34775), .Z(n34752) );
  HS65_LH_IVX2 U19011 ( .A(n34752), .Z(n34753) );
  HS65_LH_IVX2 U19012 ( .A(n34777), .Z(n34754) );
  HS65_LH_IVX2 U19013 ( .A(n34754), .Z(n34755) );
  HS65_LH_IVX2 U19014 ( .A(n34779), .Z(n34756) );
  HS65_LH_IVX2 U19015 ( .A(n34756), .Z(n34757) );
  HS65_LH_IVX2 U19016 ( .A(n34781), .Z(n34758) );
  HS65_LH_IVX2 U19017 ( .A(n34758), .Z(n34759) );
  HS65_LH_IVX2 U19018 ( .A(n34783), .Z(n34760) );
  HS65_LH_IVX2 U19019 ( .A(n34760), .Z(n34761) );
  HS65_LH_IVX2 U19020 ( .A(n34785), .Z(n34762) );
  HS65_LH_IVX2 U19021 ( .A(n34762), .Z(n34763) );
  HS65_LH_IVX2 U19022 ( .A(n34787), .Z(n34764) );
  HS65_LH_IVX2 U19023 ( .A(n34764), .Z(n34765) );
  HS65_LH_IVX2 U19024 ( .A(n34789), .Z(n34766) );
  HS65_LH_IVX2 U19025 ( .A(n34766), .Z(n34767) );
  HS65_LH_IVX2 U19026 ( .A(n34791), .Z(n34768) );
  HS65_LH_IVX2 U19027 ( .A(n34768), .Z(n34769) );
  HS65_LH_IVX2 U19028 ( .A(n34793), .Z(n34770) );
  HS65_LH_IVX2 U19029 ( .A(n34770), .Z(n34771) );
  HS65_LH_IVX2 U19030 ( .A(n34795), .Z(n34772) );
  HS65_LH_IVX2 U19031 ( .A(n34772), .Z(n34773) );
  HS65_LH_IVX2 U19032 ( .A(n34797), .Z(n34774) );
  HS65_LH_IVX2 U19033 ( .A(n34774), .Z(n34775) );
  HS65_LH_IVX2 U19034 ( .A(n34799), .Z(n34776) );
  HS65_LH_IVX2 U19035 ( .A(n34776), .Z(n34777) );
  HS65_LH_IVX2 U19036 ( .A(n34801), .Z(n34778) );
  HS65_LH_IVX2 U19037 ( .A(n34778), .Z(n34779) );
  HS65_LH_IVX2 U19038 ( .A(n34803), .Z(n34780) );
  HS65_LH_IVX2 U19039 ( .A(n34780), .Z(n34781) );
  HS65_LH_IVX2 U19040 ( .A(n34805), .Z(n34782) );
  HS65_LH_IVX2 U19041 ( .A(n34782), .Z(n34783) );
  HS65_LH_IVX2 U19042 ( .A(n34807), .Z(n34784) );
  HS65_LH_IVX2 U19043 ( .A(n34784), .Z(n34785) );
  HS65_LH_IVX2 U19044 ( .A(n34809), .Z(n34786) );
  HS65_LH_IVX2 U19045 ( .A(n34786), .Z(n34787) );
  HS65_LH_IVX2 U19046 ( .A(n34811), .Z(n34788) );
  HS65_LH_IVX2 U19047 ( .A(n34788), .Z(n34789) );
  HS65_LH_IVX2 U19048 ( .A(n34813), .Z(n34790) );
  HS65_LH_IVX2 U19049 ( .A(n34790), .Z(n34791) );
  HS65_LH_IVX2 U19050 ( .A(n34815), .Z(n34792) );
  HS65_LH_IVX2 U19051 ( .A(n34792), .Z(n34793) );
  HS65_LH_IVX2 U19052 ( .A(n34817), .Z(n34794) );
  HS65_LH_IVX2 U19053 ( .A(n34794), .Z(n34795) );
  HS65_LH_IVX2 U19054 ( .A(n34819), .Z(n34796) );
  HS65_LH_IVX2 U19055 ( .A(n34796), .Z(n34797) );
  HS65_LH_IVX2 U19056 ( .A(n34821), .Z(n34798) );
  HS65_LH_IVX2 U19057 ( .A(n34798), .Z(n34799) );
  HS65_LH_IVX2 U19058 ( .A(n34823), .Z(n34800) );
  HS65_LH_IVX2 U19059 ( .A(n34800), .Z(n34801) );
  HS65_LH_IVX2 U19060 ( .A(n34825), .Z(n34802) );
  HS65_LH_IVX2 U19061 ( .A(n34802), .Z(n34803) );
  HS65_LH_IVX2 U19062 ( .A(n34827), .Z(n34804) );
  HS65_LH_IVX2 U19063 ( .A(n34804), .Z(n34805) );
  HS65_LH_IVX2 U19064 ( .A(n34829), .Z(n34806) );
  HS65_LH_IVX2 U19065 ( .A(n34806), .Z(n34807) );
  HS65_LH_IVX2 U19066 ( .A(n34831), .Z(n34808) );
  HS65_LH_IVX2 U19067 ( .A(n34808), .Z(n34809) );
  HS65_LH_IVX2 U19068 ( .A(n34833), .Z(n34810) );
  HS65_LH_IVX2 U19069 ( .A(n34810), .Z(n34811) );
  HS65_LH_IVX2 U19070 ( .A(n34835), .Z(n34812) );
  HS65_LH_IVX2 U19071 ( .A(n34812), .Z(n34813) );
  HS65_LH_IVX2 U19072 ( .A(n34837), .Z(n34814) );
  HS65_LH_IVX2 U19073 ( .A(n34814), .Z(n34815) );
  HS65_LH_IVX2 U19074 ( .A(n34839), .Z(n34816) );
  HS65_LH_IVX2 U19075 ( .A(n34816), .Z(n34817) );
  HS65_LH_IVX2 U19076 ( .A(n34841), .Z(n34818) );
  HS65_LH_IVX2 U19077 ( .A(n34818), .Z(n34819) );
  HS65_LH_IVX2 U19078 ( .A(n34843), .Z(n34820) );
  HS65_LH_IVX2 U19079 ( .A(n34820), .Z(n34821) );
  HS65_LH_IVX2 U19080 ( .A(n34845), .Z(n34822) );
  HS65_LH_IVX2 U19081 ( .A(n34822), .Z(n34823) );
  HS65_LH_IVX2 U19082 ( .A(n34847), .Z(n34824) );
  HS65_LH_IVX2 U19083 ( .A(n34824), .Z(n34825) );
  HS65_LH_IVX2 U19084 ( .A(n34849), .Z(n34826) );
  HS65_LH_IVX2 U19085 ( .A(n34826), .Z(n34827) );
  HS65_LH_IVX2 U19086 ( .A(n34851), .Z(n34828) );
  HS65_LH_IVX2 U19087 ( .A(n34828), .Z(n34829) );
  HS65_LH_IVX2 U19088 ( .A(n34853), .Z(n34830) );
  HS65_LH_IVX2 U19089 ( .A(n34830), .Z(n34831) );
  HS65_LH_IVX2 U19090 ( .A(n34855), .Z(n34832) );
  HS65_LH_IVX2 U19091 ( .A(n34832), .Z(n34833) );
  HS65_LH_IVX2 U19092 ( .A(n34857), .Z(n34834) );
  HS65_LH_IVX2 U19093 ( .A(n34834), .Z(n34835) );
  HS65_LH_IVX2 U19094 ( .A(n34859), .Z(n34836) );
  HS65_LH_IVX2 U19095 ( .A(n34836), .Z(n34837) );
  HS65_LH_IVX2 U19096 ( .A(n34861), .Z(n34838) );
  HS65_LH_IVX2 U19097 ( .A(n34838), .Z(n34839) );
  HS65_LH_IVX2 U19098 ( .A(n34863), .Z(n34840) );
  HS65_LH_IVX2 U19099 ( .A(n34840), .Z(n34841) );
  HS65_LH_IVX2 U19100 ( .A(n34865), .Z(n34842) );
  HS65_LH_IVX2 U19101 ( .A(n34842), .Z(n34843) );
  HS65_LH_IVX2 U19102 ( .A(n34867), .Z(n34844) );
  HS65_LH_IVX2 U19103 ( .A(n34844), .Z(n34845) );
  HS65_LH_IVX2 U19104 ( .A(n34869), .Z(n34846) );
  HS65_LH_IVX2 U19105 ( .A(n34846), .Z(n34847) );
  HS65_LH_IVX2 U19106 ( .A(n34871), .Z(n34848) );
  HS65_LH_IVX2 U19107 ( .A(n34848), .Z(n34849) );
  HS65_LH_IVX2 U19108 ( .A(n34873), .Z(n34850) );
  HS65_LH_IVX2 U19109 ( .A(n34850), .Z(n34851) );
  HS65_LH_IVX2 U19110 ( .A(n34875), .Z(n34852) );
  HS65_LH_IVX2 U19111 ( .A(n34852), .Z(n34853) );
  HS65_LH_IVX2 U19112 ( .A(n34877), .Z(n34854) );
  HS65_LH_IVX2 U19113 ( .A(n34854), .Z(n34855) );
  HS65_LH_IVX2 U19114 ( .A(n34879), .Z(n34856) );
  HS65_LH_IVX2 U19115 ( .A(n34856), .Z(n34857) );
  HS65_LH_IVX2 U19116 ( .A(n34881), .Z(n34858) );
  HS65_LH_IVX2 U19117 ( .A(n34858), .Z(n34859) );
  HS65_LH_IVX2 U19118 ( .A(n34883), .Z(n34860) );
  HS65_LH_IVX2 U19119 ( .A(n34860), .Z(n34861) );
  HS65_LH_IVX2 U19120 ( .A(n34885), .Z(n34862) );
  HS65_LH_IVX2 U19121 ( .A(n34862), .Z(n34863) );
  HS65_LH_IVX2 U19122 ( .A(n34887), .Z(n34864) );
  HS65_LH_IVX2 U19123 ( .A(n34864), .Z(n34865) );
  HS65_LH_IVX2 U19124 ( .A(n34889), .Z(n34866) );
  HS65_LH_IVX2 U19125 ( .A(n34866), .Z(n34867) );
  HS65_LH_IVX2 U19126 ( .A(n34891), .Z(n34868) );
  HS65_LH_IVX2 U19127 ( .A(n34868), .Z(n34869) );
  HS65_LH_IVX2 U19128 ( .A(n34893), .Z(n34870) );
  HS65_LH_IVX2 U19129 ( .A(n34870), .Z(n34871) );
  HS65_LH_IVX2 U19130 ( .A(n34895), .Z(n34872) );
  HS65_LH_IVX2 U19131 ( .A(n34872), .Z(n34873) );
  HS65_LH_IVX2 U19132 ( .A(n34897), .Z(n34874) );
  HS65_LH_IVX2 U19133 ( .A(n34874), .Z(n34875) );
  HS65_LH_IVX2 U19134 ( .A(n34899), .Z(n34876) );
  HS65_LH_IVX2 U19135 ( .A(n34876), .Z(n34877) );
  HS65_LH_IVX2 U19136 ( .A(n34901), .Z(n34878) );
  HS65_LH_IVX2 U19137 ( .A(n34878), .Z(n34879) );
  HS65_LH_IVX2 U19138 ( .A(n34903), .Z(n34880) );
  HS65_LH_IVX2 U19139 ( .A(n34880), .Z(n34881) );
  HS65_LH_IVX2 U19140 ( .A(n34905), .Z(n34882) );
  HS65_LH_IVX2 U19141 ( .A(n34882), .Z(n34883) );
  HS65_LH_IVX2 U19142 ( .A(n34907), .Z(n34884) );
  HS65_LH_IVX2 U19143 ( .A(n34884), .Z(n34885) );
  HS65_LH_IVX2 U19144 ( .A(n34909), .Z(n34886) );
  HS65_LH_IVX2 U19145 ( .A(n34886), .Z(n34887) );
  HS65_LH_IVX2 U19146 ( .A(n34911), .Z(n34888) );
  HS65_LH_IVX2 U19147 ( .A(n34888), .Z(n34889) );
  HS65_LH_IVX2 U19148 ( .A(n34913), .Z(n34890) );
  HS65_LH_IVX2 U19149 ( .A(n34890), .Z(n34891) );
  HS65_LH_IVX2 U19150 ( .A(n34915), .Z(n34892) );
  HS65_LH_IVX2 U19151 ( .A(n34892), .Z(n34893) );
  HS65_LH_IVX2 U19152 ( .A(n34917), .Z(n34894) );
  HS65_LH_IVX2 U19153 ( .A(n34894), .Z(n34895) );
  HS65_LH_IVX2 U19154 ( .A(n34919), .Z(n34896) );
  HS65_LH_IVX2 U19155 ( .A(n34896), .Z(n34897) );
  HS65_LH_IVX2 U19156 ( .A(n34921), .Z(n34898) );
  HS65_LH_IVX2 U19157 ( .A(n34898), .Z(n34899) );
  HS65_LH_IVX2 U19158 ( .A(n34923), .Z(n34900) );
  HS65_LH_IVX2 U19159 ( .A(n34900), .Z(n34901) );
  HS65_LH_IVX2 U19160 ( .A(n34925), .Z(n34902) );
  HS65_LH_IVX2 U19161 ( .A(n34902), .Z(n34903) );
  HS65_LH_IVX2 U19162 ( .A(n34927), .Z(n34904) );
  HS65_LH_IVX2 U19163 ( .A(n34904), .Z(n34905) );
  HS65_LH_IVX2 U19164 ( .A(n34929), .Z(n34906) );
  HS65_LH_IVX2 U19165 ( .A(n34906), .Z(n34907) );
  HS65_LH_IVX2 U19166 ( .A(n34931), .Z(n34908) );
  HS65_LH_IVX2 U19167 ( .A(n34908), .Z(n34909) );
  HS65_LH_IVX2 U19168 ( .A(n34933), .Z(n34910) );
  HS65_LH_IVX2 U19169 ( .A(n34910), .Z(n34911) );
  HS65_LH_IVX2 U19170 ( .A(n34935), .Z(n34912) );
  HS65_LH_IVX2 U19171 ( .A(n34912), .Z(n34913) );
  HS65_LH_IVX2 U19172 ( .A(n34937), .Z(n34914) );
  HS65_LH_IVX2 U19173 ( .A(n34914), .Z(n34915) );
  HS65_LH_IVX2 U19174 ( .A(n34939), .Z(n34916) );
  HS65_LH_IVX2 U19175 ( .A(n34916), .Z(n34917) );
  HS65_LH_IVX2 U19176 ( .A(n34941), .Z(n34918) );
  HS65_LH_IVX2 U19177 ( .A(n34918), .Z(n34919) );
  HS65_LH_IVX2 U19178 ( .A(n34943), .Z(n34920) );
  HS65_LH_IVX2 U19179 ( .A(n34920), .Z(n34921) );
  HS65_LH_IVX2 U19180 ( .A(n34945), .Z(n34922) );
  HS65_LH_IVX2 U19181 ( .A(n34922), .Z(n34923) );
  HS65_LH_IVX2 U19182 ( .A(n34947), .Z(n34924) );
  HS65_LH_IVX2 U19183 ( .A(n34924), .Z(n34925) );
  HS65_LH_IVX2 U19184 ( .A(n34949), .Z(n34926) );
  HS65_LH_IVX2 U19185 ( .A(n34926), .Z(n34927) );
  HS65_LH_IVX2 U19186 ( .A(n34951), .Z(n34928) );
  HS65_LH_IVX2 U19187 ( .A(n34928), .Z(n34929) );
  HS65_LH_IVX2 U19188 ( .A(n34953), .Z(n34930) );
  HS65_LH_IVX2 U19189 ( .A(n34930), .Z(n34931) );
  HS65_LH_IVX2 U19190 ( .A(n34955), .Z(n34932) );
  HS65_LH_IVX2 U19191 ( .A(n34932), .Z(n34933) );
  HS65_LH_IVX2 U19192 ( .A(n34957), .Z(n34934) );
  HS65_LH_IVX2 U19193 ( .A(n34934), .Z(n34935) );
  HS65_LH_IVX2 U19194 ( .A(n34959), .Z(n34936) );
  HS65_LH_IVX2 U19195 ( .A(n34936), .Z(n34937) );
  HS65_LH_IVX2 U19196 ( .A(n34961), .Z(n34938) );
  HS65_LH_IVX2 U19197 ( .A(n34938), .Z(n34939) );
  HS65_LH_IVX2 U19198 ( .A(n34963), .Z(n34940) );
  HS65_LH_IVX2 U19199 ( .A(n34940), .Z(n34941) );
  HS65_LH_IVX2 U19200 ( .A(n34965), .Z(n34942) );
  HS65_LH_IVX2 U19201 ( .A(n34942), .Z(n34943) );
  HS65_LH_IVX2 U19202 ( .A(n34967), .Z(n34944) );
  HS65_LH_IVX2 U19203 ( .A(n34944), .Z(n34945) );
  HS65_LH_IVX2 U19204 ( .A(n34969), .Z(n34946) );
  HS65_LH_IVX2 U19205 ( .A(n34946), .Z(n34947) );
  HS65_LH_IVX2 U19206 ( .A(n34971), .Z(n34948) );
  HS65_LH_IVX2 U19207 ( .A(n34948), .Z(n34949) );
  HS65_LH_IVX2 U19208 ( .A(n34973), .Z(n34950) );
  HS65_LH_IVX2 U19209 ( .A(n34950), .Z(n34951) );
  HS65_LH_IVX2 U19210 ( .A(n34975), .Z(n34952) );
  HS65_LH_IVX2 U19211 ( .A(n34952), .Z(n34953) );
  HS65_LH_IVX2 U19212 ( .A(n34977), .Z(n34954) );
  HS65_LH_IVX2 U19213 ( .A(n34954), .Z(n34955) );
  HS65_LH_IVX2 U19214 ( .A(n34979), .Z(n34956) );
  HS65_LH_IVX2 U19215 ( .A(n34956), .Z(n34957) );
  HS65_LH_IVX2 U19216 ( .A(n34981), .Z(n34958) );
  HS65_LH_IVX2 U19217 ( .A(n34958), .Z(n34959) );
  HS65_LH_IVX2 U19218 ( .A(n34983), .Z(n34960) );
  HS65_LH_IVX2 U19219 ( .A(n34960), .Z(n34961) );
  HS65_LH_IVX2 U19220 ( .A(n34985), .Z(n34962) );
  HS65_LH_IVX2 U19221 ( .A(n34962), .Z(n34963) );
  HS65_LH_IVX2 U19222 ( .A(n34987), .Z(n34964) );
  HS65_LH_IVX2 U19223 ( .A(n34964), .Z(n34965) );
  HS65_LH_IVX2 U19224 ( .A(n34989), .Z(n34966) );
  HS65_LH_IVX2 U19225 ( .A(n34966), .Z(n34967) );
  HS65_LH_IVX2 U19226 ( .A(n34991), .Z(n34968) );
  HS65_LH_IVX2 U19227 ( .A(n34968), .Z(n34969) );
  HS65_LH_IVX2 U19228 ( .A(n34993), .Z(n34970) );
  HS65_LH_IVX2 U19229 ( .A(n34970), .Z(n34971) );
  HS65_LH_IVX2 U19230 ( .A(n34995), .Z(n34972) );
  HS65_LH_IVX2 U19231 ( .A(n34972), .Z(n34973) );
  HS65_LH_IVX2 U19232 ( .A(n34997), .Z(n34974) );
  HS65_LH_IVX2 U19233 ( .A(n34974), .Z(n34975) );
  HS65_LH_IVX2 U19234 ( .A(n34999), .Z(n34976) );
  HS65_LH_IVX2 U19235 ( .A(n34976), .Z(n34977) );
  HS65_LH_IVX2 U19236 ( .A(n35001), .Z(n34978) );
  HS65_LH_IVX2 U19237 ( .A(n34978), .Z(n34979) );
  HS65_LH_IVX2 U19238 ( .A(n35003), .Z(n34980) );
  HS65_LH_IVX2 U19239 ( .A(n34980), .Z(n34981) );
  HS65_LH_IVX2 U19240 ( .A(n35005), .Z(n34982) );
  HS65_LH_IVX2 U19241 ( .A(n34982), .Z(n34983) );
  HS65_LH_IVX2 U19242 ( .A(n35007), .Z(n34984) );
  HS65_LH_IVX2 U19243 ( .A(n34984), .Z(n34985) );
  HS65_LH_IVX2 U19244 ( .A(n35009), .Z(n34986) );
  HS65_LH_IVX2 U19245 ( .A(n34986), .Z(n34987) );
  HS65_LH_IVX2 U19246 ( .A(n35011), .Z(n34988) );
  HS65_LH_IVX2 U19247 ( .A(n34988), .Z(n34989) );
  HS65_LH_IVX2 U19248 ( .A(n35013), .Z(n34990) );
  HS65_LH_IVX2 U19249 ( .A(n34990), .Z(n34991) );
  HS65_LH_IVX2 U19250 ( .A(n35015), .Z(n34992) );
  HS65_LH_IVX2 U19251 ( .A(n34992), .Z(n34993) );
  HS65_LH_IVX2 U19252 ( .A(n35017), .Z(n34994) );
  HS65_LH_IVX2 U19253 ( .A(n34994), .Z(n34995) );
  HS65_LH_IVX2 U19254 ( .A(n35019), .Z(n34996) );
  HS65_LH_IVX2 U19255 ( .A(n34996), .Z(n34997) );
  HS65_LH_IVX2 U19256 ( .A(n35021), .Z(n34998) );
  HS65_LH_IVX2 U19257 ( .A(n34998), .Z(n34999) );
  HS65_LH_IVX2 U19259 ( .A(n35023), .Z(n35000) );
  HS65_LH_IVX2 U19260 ( .A(n35000), .Z(n35001) );
  HS65_LH_IVX2 U19261 ( .A(n35025), .Z(n35002) );
  HS65_LH_IVX2 U19262 ( .A(n35002), .Z(n35003) );
  HS65_LH_IVX2 U19263 ( .A(n35058), .Z(n35004) );
  HS65_LH_IVX2 U19264 ( .A(n35004), .Z(n35005) );
  HS65_LH_IVX2 U19265 ( .A(n35027), .Z(n35006) );
  HS65_LH_IVX2 U19266 ( .A(n35006), .Z(n35007) );
  HS65_LH_IVX2 U19267 ( .A(n35044), .Z(n35008) );
  HS65_LH_IVX2 U19268 ( .A(n35008), .Z(n35009) );
  HS65_LH_IVX2 U19269 ( .A(n35031), .Z(n35010) );
  HS65_LH_IVX2 U19270 ( .A(n35010), .Z(n35011) );
  HS65_LH_IVX2 U19271 ( .A(n35046), .Z(n35012) );
  HS65_LH_IVX2 U19272 ( .A(n35012), .Z(n35013) );
  HS65_LH_IVX2 U19273 ( .A(n35033), .Z(n35014) );
  HS65_LH_IVX2 U19274 ( .A(n35014), .Z(n35015) );
  HS65_LH_IVX2 U19275 ( .A(n35035), .Z(n35016) );
  HS65_LH_IVX2 U19276 ( .A(n35016), .Z(n35017) );
  HS65_LH_IVX2 U19277 ( .A(n35054), .Z(n35018) );
  HS65_LH_IVX2 U19278 ( .A(n35018), .Z(n35019) );
  HS65_LH_IVX2 U19279 ( .A(n35037), .Z(n35020) );
  HS65_LH_IVX2 U19280 ( .A(n35020), .Z(n35021) );
  HS65_LH_IVX2 U19281 ( .A(n35055), .Z(n35022) );
  HS65_LH_IVX2 U19282 ( .A(n35022), .Z(n35023) );
  HS65_LH_IVX2 U19283 ( .A(n15730), .Z(n35024) );
  HS65_LH_IVX2 U19284 ( .A(n35024), .Z(n35025) );
  HS65_LH_IVX2 U19285 ( .A(n35040), .Z(n35026) );
  HS65_LH_IVX2 U19286 ( .A(n35026), .Z(n35027) );
  HS65_LH_IVX2 U19287 ( .A(n213), .Z(n35028) );
  HS65_LH_IVX2 U19288 ( .A(n35028), .Z(n35029) );
  HS65_LH_IVX2 U19289 ( .A(n35042), .Z(n35030) );
  HS65_LH_IVX2 U19290 ( .A(n35030), .Z(n35031) );
  HS65_LH_IVX2 U19291 ( .A(n35048), .Z(n35032) );
  HS65_LH_IVX2 U19292 ( .A(n35032), .Z(n35033) );
  HS65_LH_IVX2 U19293 ( .A(n35050), .Z(n35034) );
  HS65_LH_IVX2 U19294 ( .A(n35034), .Z(n35035) );
  HS65_LH_IVX2 U19295 ( .A(n35052), .Z(n35036) );
  HS65_LH_IVX2 U19296 ( .A(n35036), .Z(n35037) );
  HS65_LH_BFX2 U19297 ( .A(n34685), .Z(n35038) );
  HS65_LH_IVX2 U19298 ( .A(n17847), .Z(n35039) );
  HS65_LH_IVX2 U19299 ( .A(n35039), .Z(n35040) );
  HS65_LH_IVX2 U19300 ( .A(n35060), .Z(n35041) );
  HS65_LH_IVX2 U19301 ( .A(n35041), .Z(n35042) );
  HS65_LH_IVX2 U19302 ( .A(n17443), .Z(n35043) );
  HS65_LH_IVX2 U19303 ( .A(n35043), .Z(n35044) );
  HS65_LH_IVX2 U19304 ( .A(n17442), .Z(n35045) );
  HS65_LH_IVX2 U19305 ( .A(n35045), .Z(n35046) );
  HS65_LH_IVX2 U19306 ( .A(n17641), .Z(n35047) );
  HS65_LH_IVX2 U19307 ( .A(n35047), .Z(n35048) );
  HS65_LH_IVX2 U19308 ( .A(n35062), .Z(n35049) );
  HS65_LH_IVX2 U19309 ( .A(n35049), .Z(n35050) );
  HS65_LH_IVX2 U19310 ( .A(n35064), .Z(n35051) );
  HS65_LH_IVX2 U19311 ( .A(n35051), .Z(n35052) );
  HS65_LH_IVX2 U19312 ( .A(n17441), .Z(n35053) );
  HS65_LH_IVX2 U19313 ( .A(n35053), .Z(n35054) );
  HS65_LH_BFX2 U19314 ( .A(n34712), .Z(n35055) );
  HS65_LH_BFX2 U19315 ( .A(n35038), .Z(n35056) );
  HS65_LH_IVX2 U19316 ( .A(n35056), .Z(n35057) );
  HS65_LH_IVX2 U19317 ( .A(n35057), .Z(n35058) );
  HS65_LH_IVX2 U19318 ( .A(n17725), .Z(n35059) );
  HS65_LH_IVX2 U19319 ( .A(n35059), .Z(n35060) );
  HS65_LH_IVX2 U19320 ( .A(n17374), .Z(n35061) );
  HS65_LH_IVX2 U19321 ( .A(n35061), .Z(n35062) );
  HS65_LH_IVX2 U19322 ( .A(n17269), .Z(n35063) );
  HS65_LH_IVX2 U19323 ( .A(n35063), .Z(n35064) );
  HS65_LH_BFX2 U19324 ( .A(n35067), .Z(n35065) );
  HS65_LH_BFX2 U19325 ( .A(n17849), .Z(n35066) );
  HS65_LH_BFX2 U19326 ( .A(n35069), .Z(n35067) );
  HS65_LH_BFX2 U19327 ( .A(n35066), .Z(n35068) );
  HS65_LH_BFX2 U19328 ( .A(n35071), .Z(n35069) );
  HS65_LH_BFX2 U19329 ( .A(n35068), .Z(n35070) );
  HS65_LH_BFX2 U19330 ( .A(n35073), .Z(n35071) );
  HS65_LH_BFX2 U19331 ( .A(n35070), .Z(n35072) );
  HS65_LH_BFX2 U19332 ( .A(n35075), .Z(n35073) );
  HS65_LH_BFX2 U19333 ( .A(n35072), .Z(n35074) );
  HS65_LH_BFX2 U19334 ( .A(n35077), .Z(n35075) );
  HS65_LH_BFX2 U19335 ( .A(n35074), .Z(n35076) );
  HS65_LH_BFX2 U19336 ( .A(n35079), .Z(n35077) );
  HS65_LH_BFX2 U19337 ( .A(n35076), .Z(n35078) );
  HS65_LH_BFX2 U19338 ( .A(n35081), .Z(n35079) );
  HS65_LH_BFX2 U19339 ( .A(n35078), .Z(n35080) );
  HS65_LH_BFX2 U19340 ( .A(n35083), .Z(n35081) );
  HS65_LH_BFX2 U19341 ( .A(n35080), .Z(n35082) );
  HS65_LH_BFX2 U19342 ( .A(n35085), .Z(n35083) );
  HS65_LH_BFX2 U19343 ( .A(n35082), .Z(n35084) );
  HS65_LH_BFX2 U19344 ( .A(n35087), .Z(n35085) );
  HS65_LH_BFX2 U19345 ( .A(n35084), .Z(n35086) );
  HS65_LH_BFX2 U19346 ( .A(n35089), .Z(n35087) );
  HS65_LH_BFX2 U19347 ( .A(n35086), .Z(n35088) );
  HS65_LH_BFX2 U19348 ( .A(n35091), .Z(n35089) );
  HS65_LH_BFX2 U19349 ( .A(n35088), .Z(n35090) );
  HS65_LH_BFX2 U19350 ( .A(n35093), .Z(n35091) );
  HS65_LH_BFX2 U19351 ( .A(n35090), .Z(n35092) );
  HS65_LH_BFX2 U19352 ( .A(n35095), .Z(n35093) );
  HS65_LH_BFX2 U19353 ( .A(n35092), .Z(n35094) );
  HS65_LH_BFX2 U19354 ( .A(n35097), .Z(n35095) );
  HS65_LH_BFX2 U19355 ( .A(n35094), .Z(n35096) );
  HS65_LH_BFX2 U19356 ( .A(n35099), .Z(n35097) );
  HS65_LH_BFX2 U19357 ( .A(n35096), .Z(n35098) );
  HS65_LH_BFX2 U19358 ( .A(n35102), .Z(n35099) );
  HS65_LH_BFX2 U19359 ( .A(n35098), .Z(n35100) );
  HS65_LH_IVX2 U19360 ( .A(n15389), .Z(n35101) );
  HS65_LH_IVX2 U19361 ( .A(n35101), .Z(n35102) );
  HS65_LH_BFX2 U19362 ( .A(n35100), .Z(n35103) );
  HS65_LH_BFX2 U19363 ( .A(n35103), .Z(n35104) );
  HS65_LH_IVX2 U19364 ( .A(n35107), .Z(n35105) );
  HS65_LH_IVX2 U19365 ( .A(n35105), .Z(n35106) );
  HS65_LH_BFX2 U19366 ( .A(n35104), .Z(n35107) );
  HS65_LH_BFX2 U19367 ( .A(n35110), .Z(n35108) );
  HS65_LH_IVX2 U19368 ( .A(n35113), .Z(n35109) );
  HS65_LH_IVX2 U19369 ( .A(n35109), .Z(n35110) );
  HS65_LH_BFX2 U19370 ( .A(n35112), .Z(n35111) );
  HS65_LH_BFX2 U19371 ( .A(n35114), .Z(n35112) );
  HS65_LH_BFX2 U19372 ( .A(n35115), .Z(n35113) );
  HS65_LH_BFX2 U19373 ( .A(n35116), .Z(n35114) );
  HS65_LH_BFX2 U19374 ( .A(n35117), .Z(n35115) );
  HS65_LH_BFX2 U19375 ( .A(n35118), .Z(n35116) );
  HS65_LH_BFX2 U19376 ( .A(n35119), .Z(n35117) );
  HS65_LH_BFX2 U19377 ( .A(n35120), .Z(n35118) );
  HS65_LH_BFX2 U19378 ( .A(n35121), .Z(n35119) );
  HS65_LH_BFX2 U19379 ( .A(n35122), .Z(n35120) );
  HS65_LH_BFX2 U19380 ( .A(n35123), .Z(n35121) );
  HS65_LH_BFX2 U19381 ( .A(n35124), .Z(n35122) );
  HS65_LH_BFX2 U19382 ( .A(n35125), .Z(n35123) );
  HS65_LH_BFX2 U19383 ( .A(n35126), .Z(n35124) );
  HS65_LH_BFX2 U19384 ( .A(n35127), .Z(n35125) );
  HS65_LH_BFX2 U19385 ( .A(n35128), .Z(n35126) );
  HS65_LH_BFX2 U19386 ( .A(n35129), .Z(n35127) );
  HS65_LH_BFX2 U19387 ( .A(n35130), .Z(n35128) );
  HS65_LH_BFX2 U19388 ( .A(n35131), .Z(n35129) );
  HS65_LH_BFX2 U19389 ( .A(n35132), .Z(n35130) );
  HS65_LH_BFX2 U19391 ( .A(n35133), .Z(n35131) );
  HS65_LH_BFX2 U19392 ( .A(n35134), .Z(n35132) );
  HS65_LH_BFX2 U19393 ( .A(n35135), .Z(n35133) );
  HS65_LH_BFX2 U19394 ( .A(n35136), .Z(n35134) );
  HS65_LH_BFX2 U19395 ( .A(n35137), .Z(n35135) );
  HS65_LH_BFX2 U19396 ( .A(n35138), .Z(n35136) );
  HS65_LH_BFX2 U19397 ( .A(n35139), .Z(n35137) );
  HS65_LH_BFX2 U19398 ( .A(n35140), .Z(n35138) );
  HS65_LH_BFX2 U19399 ( .A(n35141), .Z(n35139) );
  HS65_LH_BFX2 U19400 ( .A(n35142), .Z(n35140) );
  HS65_LH_BFX2 U19401 ( .A(n35143), .Z(n35141) );
  HS65_LH_BFX2 U19402 ( .A(n35144), .Z(n35142) );
  HS65_LH_BFX2 U19403 ( .A(n35145), .Z(n35143) );
  HS65_LH_BFX2 U19404 ( .A(n35146), .Z(n35144) );
  HS65_LH_BFX2 U19405 ( .A(n35147), .Z(n35145) );
  HS65_LH_BFX2 U19406 ( .A(n35148), .Z(n35146) );
  HS65_LH_BFX2 U19407 ( .A(n35149), .Z(n35147) );
  HS65_LH_BFX2 U19408 ( .A(n35150), .Z(n35148) );
  HS65_LH_BFX2 U19409 ( .A(n14750), .Z(n35149) );
  HS65_LH_BFX2 U19410 ( .A(n35151), .Z(n35150) );
  HS65_LH_BFX2 U19411 ( .A(n17925), .Z(n35151) );
  HS65_LH_BFX2 U19412 ( .A(n35154), .Z(n35152) );
  HS65_LH_IVX2 U19413 ( .A(n35157), .Z(n35153) );
  HS65_LH_IVX2 U19414 ( .A(n35153), .Z(n35154) );
  HS65_LH_BFX2 U19415 ( .A(n35156), .Z(n35155) );
  HS65_LH_BFX2 U19416 ( .A(n35158), .Z(n35156) );
  HS65_LH_BFX2 U19417 ( .A(n35159), .Z(n35157) );
  HS65_LH_BFX2 U19418 ( .A(n35160), .Z(n35158) );
  HS65_LH_BFX2 U19419 ( .A(n35161), .Z(n35159) );
  HS65_LH_BFX2 U19420 ( .A(n35162), .Z(n35160) );
  HS65_LH_BFX2 U19421 ( .A(n35163), .Z(n35161) );
  HS65_LH_BFX2 U19422 ( .A(n35164), .Z(n35162) );
  HS65_LH_BFX2 U19423 ( .A(n35165), .Z(n35163) );
  HS65_LH_BFX2 U19424 ( .A(n35166), .Z(n35164) );
  HS65_LH_BFX2 U19425 ( .A(n35167), .Z(n35165) );
  HS65_LH_BFX2 U19426 ( .A(n35168), .Z(n35166) );
  HS65_LH_BFX2 U19427 ( .A(n35169), .Z(n35167) );
  HS65_LH_BFX2 U19428 ( .A(n35170), .Z(n35168) );
  HS65_LH_BFX2 U19429 ( .A(n35171), .Z(n35169) );
  HS65_LH_BFX2 U19430 ( .A(n35172), .Z(n35170) );
  HS65_LH_BFX2 U19431 ( .A(n35173), .Z(n35171) );
  HS65_LH_BFX2 U19432 ( .A(n35174), .Z(n35172) );
  HS65_LH_BFX2 U19433 ( .A(n35175), .Z(n35173) );
  HS65_LH_BFX2 U19434 ( .A(n35176), .Z(n35174) );
  HS65_LH_BFX2 U19435 ( .A(n35177), .Z(n35175) );
  HS65_LH_BFX2 U19436 ( .A(n35178), .Z(n35176) );
  HS65_LH_BFX2 U19437 ( .A(n35179), .Z(n35177) );
  HS65_LH_BFX2 U19438 ( .A(n35180), .Z(n35178) );
  HS65_LH_BFX2 U19439 ( .A(n35181), .Z(n35179) );
  HS65_LH_BFX2 U19440 ( .A(n35182), .Z(n35180) );
  HS65_LH_BFX2 U19441 ( .A(n35183), .Z(n35181) );
  HS65_LH_BFX2 U19442 ( .A(n35184), .Z(n35182) );
  HS65_LH_BFX2 U19443 ( .A(n35185), .Z(n35183) );
  HS65_LH_BFX2 U19444 ( .A(n35186), .Z(n35184) );
  HS65_LH_BFX2 U19445 ( .A(n35187), .Z(n35185) );
  HS65_LH_BFX2 U19446 ( .A(n35188), .Z(n35186) );
  HS65_LH_BFX2 U19447 ( .A(n35189), .Z(n35187) );
  HS65_LH_BFX2 U19448 ( .A(n35190), .Z(n35188) );
  HS65_LH_BFX2 U19449 ( .A(n35191), .Z(n35189) );
  HS65_LH_BFX2 U19450 ( .A(n35192), .Z(n35190) );
  HS65_LH_BFX2 U19451 ( .A(n14840), .Z(n35191) );
  HS65_LH_BFX2 U19452 ( .A(n35193), .Z(n35192) );
  HS65_LH_BFX2 U19453 ( .A(n35194), .Z(n35193) );
  HS65_LH_BFX2 U19454 ( .A(n17917), .Z(n35194) );
  HS65_LH_BFX2 U19455 ( .A(n35196), .Z(n35195) );
  HS65_LH_BFX2 U19456 ( .A(n35197), .Z(n35196) );
  HS65_LH_BFX2 U19457 ( .A(n35198), .Z(n35197) );
  HS65_LH_BFX2 U19458 ( .A(n35199), .Z(n35198) );
  HS65_LH_BFX2 U19459 ( .A(n35200), .Z(n35199) );
  HS65_LH_BFX2 U19460 ( .A(n35201), .Z(n35200) );
  HS65_LH_BFX2 U19461 ( .A(n35202), .Z(n35201) );
  HS65_LH_BFX2 U19462 ( .A(n35203), .Z(n35202) );
  HS65_LH_BFX2 U19463 ( .A(n35204), .Z(n35203) );
  HS65_LH_BFX2 U19464 ( .A(n35205), .Z(n35204) );
  HS65_LH_BFX2 U19465 ( .A(n35206), .Z(n35205) );
  HS65_LH_BFX2 U19466 ( .A(n35207), .Z(n35206) );
  HS65_LH_BFX2 U19467 ( .A(n35208), .Z(n35207) );
  HS65_LH_BFX2 U19468 ( .A(n35209), .Z(n35208) );
  HS65_LH_BFX2 U19469 ( .A(n35210), .Z(n35209) );
  HS65_LH_BFX2 U19470 ( .A(n35211), .Z(n35210) );
  HS65_LH_BFX2 U19471 ( .A(n35212), .Z(n35211) );
  HS65_LH_BFX2 U19472 ( .A(n15423), .Z(n35212) );
  HS65_LH_BFX2 U19473 ( .A(n32636), .Z(n35213) );
  HS65_LH_IVX2 U19474 ( .A(n37036), .Z(n35214) );
  HS65_LH_IVX2 U19475 ( .A(n35214), .Z(n35215) );
  HS65_LH_BFX2 U19476 ( .A(n35222), .Z(n35216) );
  HS65_LH_IVX2 U19477 ( .A(n35247), .Z(n35217) );
  HS65_LH_IVX2 U19478 ( .A(n35217), .Z(n35218) );
  HS65_LH_BFX2 U19479 ( .A(n35226), .Z(n35219) );
  HS65_LH_BFX2 U19480 ( .A(n35228), .Z(n35220) );
  HS65_LH_IVX2 U19481 ( .A(n35249), .Z(n35221) );
  HS65_LH_IVX2 U19482 ( .A(n35221), .Z(n35222) );
  HS65_LH_IVX2 U19483 ( .A(n35251), .Z(n35223) );
  HS65_LH_IVX2 U19484 ( .A(n35223), .Z(n35224) );
  HS65_LH_IVX2 U19485 ( .A(n35253), .Z(n35225) );
  HS65_LH_IVX2 U19486 ( .A(n35225), .Z(n35226) );
  HS65_LH_IVX2 U19487 ( .A(n35255), .Z(n35227) );
  HS65_LH_IVX2 U19488 ( .A(n35227), .Z(n35228) );
  HS65_LH_BFX2 U19489 ( .A(n35256), .Z(n35229) );
  HS65_LH_BFX2 U19490 ( .A(n17569), .Z(n35230) );
  HS65_LH_BFX2 U19491 ( .A(n35419), .Z(n35231) );
  HS65_LH_BFX2 U19492 ( .A(n17574), .Z(n35232) );
  HS65_LH_IVX2 U19493 ( .A(n35521), .Z(n35522) );
  HS65_LH_BFX2 U19494 ( .A(n35245), .Z(n35233) );
  HS65_LH_BFX2 U19495 ( .A(n197), .Z(n35234) );
  HS65_LH_BFX2 U19496 ( .A(n31206), .Z(n35235) );
  HS65_LH_IVX2 U19497 ( .A(n35269), .Z(n35236) );
  HS65_LH_IVX2 U19498 ( .A(n35236), .Z(n35237) );
  HS65_LH_IVX2 U19499 ( .A(n35271), .Z(n35238) );
  HS65_LH_IVX2 U19500 ( .A(n35238), .Z(n35239) );
  HS65_LH_IVX2 U19501 ( .A(n35273), .Z(n35240) );
  HS65_LH_IVX2 U19502 ( .A(n35240), .Z(n35241) );
  HS65_LH_IVX2 U19503 ( .A(n37047), .Z(n35242) );
  HS65_LH_IVX2 U19504 ( .A(n35242), .Z(n35243) );
  HS65_LH_IVX2 U19505 ( .A(n35298), .Z(n35244) );
  HS65_LH_IVX2 U19506 ( .A(n35244), .Z(n35245) );
  HS65_LH_IVX2 U19507 ( .A(n35275), .Z(n35246) );
  HS65_LH_IVX2 U19508 ( .A(n35246), .Z(n35247) );
  HS65_LH_IVX2 U19509 ( .A(n35277), .Z(n35248) );
  HS65_LH_IVX2 U19510 ( .A(n35248), .Z(n35249) );
  HS65_LH_IVX2 U19511 ( .A(n35279), .Z(n35250) );
  HS65_LH_IVX2 U19512 ( .A(n35250), .Z(n35251) );
  HS65_LH_IVX2 U19513 ( .A(n35281), .Z(n35252) );
  HS65_LH_IVX2 U19514 ( .A(n35252), .Z(n35253) );
  HS65_LH_IVX2 U19515 ( .A(n35283), .Z(n35254) );
  HS65_LH_IVX2 U19516 ( .A(n35254), .Z(n35255) );
  HS65_LH_IVX2 U19517 ( .A(n40985), .Z(n35520) );
  HS65_LH_BFX2 U19518 ( .A(n35259), .Z(n35256) );
  HS65_LH_BFX2 U19519 ( .A(n35230), .Z(n35257) );
  HS65_LH_IVX2 U19520 ( .A(n35287), .Z(n35258) );
  HS65_LH_IVX2 U19521 ( .A(n35258), .Z(n35259) );
  HS65_LH_BFX2 U19522 ( .A(n17297), .Z(n35260) );
  HS65_LH_BFX2 U19523 ( .A(n35232), .Z(n35261) );
  HS65_LH_IVX2 U19524 ( .A(n35290), .Z(n35262) );
  HS65_LH_IVX2 U19525 ( .A(n35262), .Z(n35263) );
  HS65_LH_BFX2 U19526 ( .A(n35234), .Z(n35264) );
  HS65_LH_BFX2 U19527 ( .A(n35235), .Z(n35265) );
  HS65_LH_IVX2 U19528 ( .A(n35370), .Z(n35266) );
  HS65_LH_IVX2 U19529 ( .A(n35266), .Z(n35267) );
  HS65_LH_IVX2 U19530 ( .A(n35292), .Z(n35268) );
  HS65_LH_IVX2 U19531 ( .A(n35268), .Z(n35269) );
  HS65_LH_IVX2 U19532 ( .A(n35294), .Z(n35270) );
  HS65_LH_IVX2 U19533 ( .A(n35270), .Z(n35271) );
  HS65_LH_IVX2 U19534 ( .A(n35296), .Z(n35272) );
  HS65_LH_IVX2 U19535 ( .A(n35272), .Z(n35273) );
  HS65_LH_IVX2 U19536 ( .A(n35300), .Z(n35274) );
  HS65_LH_IVX2 U19537 ( .A(n35274), .Z(n35275) );
  HS65_LH_IVX2 U19538 ( .A(n35302), .Z(n35276) );
  HS65_LH_IVX2 U19539 ( .A(n35276), .Z(n35277) );
  HS65_LH_IVX2 U19540 ( .A(n35306), .Z(n35278) );
  HS65_LH_IVX2 U19541 ( .A(n35278), .Z(n35279) );
  HS65_LH_IVX2 U19542 ( .A(n35308), .Z(n35280) );
  HS65_LH_IVX2 U19543 ( .A(n35280), .Z(n35281) );
  HS65_LH_IVX2 U19544 ( .A(n35310), .Z(n35282) );
  HS65_LH_IVX2 U19545 ( .A(n35282), .Z(n35283) );
  HS65_LH_BFX2 U19546 ( .A(n35257), .Z(n35284) );
  HS65_LH_BFX2 U19547 ( .A(n35260), .Z(n35285) );
  HS65_LH_IVX2 U19548 ( .A(n35314), .Z(n35286) );
  HS65_LH_IVX2 U19549 ( .A(n35286), .Z(n35287) );
  HS65_LH_BFX2 U19550 ( .A(n35265), .Z(n35288) );
  HS65_LH_IVX2 U19551 ( .A(n35318), .Z(n35289) );
  HS65_LH_IVX2 U19552 ( .A(n35289), .Z(n35290) );
  HS65_LH_IVX2 U19553 ( .A(n35320), .Z(n35291) );
  HS65_LH_IVX2 U19554 ( .A(n35291), .Z(n35292) );
  HS65_LH_IVX2 U19555 ( .A(n35322), .Z(n35293) );
  HS65_LH_IVX2 U19556 ( .A(n35293), .Z(n35294) );
  HS65_LH_IVX2 U19557 ( .A(n35324), .Z(n35295) );
  HS65_LH_IVX2 U19558 ( .A(n35295), .Z(n35296) );
  HS65_LH_IVX2 U19559 ( .A(n35304), .Z(n35297) );
  HS65_LH_IVX2 U19560 ( .A(n35297), .Z(n35298) );
  HS65_LH_IVX2 U19561 ( .A(n35326), .Z(n35299) );
  HS65_LH_IVX2 U19562 ( .A(n35299), .Z(n35300) );
  HS65_LH_IVX2 U19563 ( .A(n35328), .Z(n35301) );
  HS65_LH_IVX2 U19564 ( .A(n35301), .Z(n35302) );
  HS65_LH_IVX2 U19565 ( .A(n35330), .Z(n35303) );
  HS65_LH_IVX2 U19566 ( .A(n35303), .Z(n35304) );
  HS65_LH_IVX2 U19567 ( .A(n35332), .Z(n35305) );
  HS65_LH_IVX2 U19568 ( .A(n35305), .Z(n35306) );
  HS65_LH_IVX2 U19569 ( .A(n35334), .Z(n35307) );
  HS65_LH_IVX2 U19570 ( .A(n35307), .Z(n35308) );
  HS65_LH_IVX2 U19571 ( .A(n35336), .Z(n35309) );
  HS65_LH_IVX2 U19572 ( .A(n35309), .Z(n35310) );
  HS65_LH_BFX2 U19573 ( .A(n35284), .Z(n35311) );
  HS65_LH_BFX2 U19574 ( .A(n35285), .Z(n35312) );
  HS65_LH_IVX2 U19575 ( .A(n35341), .Z(n35313) );
  HS65_LH_IVX2 U19576 ( .A(n35313), .Z(n35314) );
  HS65_LH_BFX2 U19577 ( .A(n35288), .Z(n35315) );
  HS65_LH_BFX2 U19578 ( .A(n35264), .Z(n35316) );
  HS65_LH_IVX2 U19579 ( .A(n35344), .Z(n35317) );
  HS65_LH_IVX2 U19580 ( .A(n35317), .Z(n35318) );
  HS65_LH_IVX2 U19581 ( .A(n35346), .Z(n35319) );
  HS65_LH_IVX2 U19582 ( .A(n35319), .Z(n35320) );
  HS65_LH_IVX2 U19583 ( .A(n35348), .Z(n35321) );
  HS65_LH_IVX2 U19584 ( .A(n35321), .Z(n35322) );
  HS65_LH_IVX2 U19585 ( .A(n35350), .Z(n35323) );
  HS65_LH_IVX2 U19586 ( .A(n35323), .Z(n35324) );
  HS65_LH_IVX2 U19587 ( .A(n35352), .Z(n35325) );
  HS65_LH_IVX2 U19588 ( .A(n35325), .Z(n35326) );
  HS65_LH_IVX2 U19589 ( .A(n35354), .Z(n35327) );
  HS65_LH_IVX2 U19590 ( .A(n35327), .Z(n35328) );
  HS65_LH_IVX2 U19591 ( .A(n35356), .Z(n35329) );
  HS65_LH_IVX2 U19592 ( .A(n35329), .Z(n35330) );
  HS65_LH_IVX2 U19593 ( .A(n35358), .Z(n35331) );
  HS65_LH_IVX2 U19594 ( .A(n35331), .Z(n35332) );
  HS65_LH_IVX2 U19595 ( .A(n35360), .Z(n35333) );
  HS65_LH_IVX2 U19596 ( .A(n35333), .Z(n35334) );
  HS65_LH_IVX2 U19597 ( .A(n35362), .Z(n35335) );
  HS65_LH_IVX2 U19598 ( .A(n35335), .Z(n35336) );
  HS65_LH_BFX2 U19599 ( .A(n35311), .Z(n35337) );
  HS65_LH_BFX2 U19600 ( .A(n35312), .Z(n35338) );
  HS65_LH_BFX2 U19601 ( .A(n35315), .Z(n35339) );
  HS65_LH_IVX2 U19602 ( .A(n35368), .Z(n35340) );
  HS65_LH_IVX2 U19603 ( .A(n35340), .Z(n35341) );
  HS65_LH_BFX2 U19604 ( .A(n35316), .Z(n35342) );
  HS65_LH_IVX2 U19605 ( .A(n35372), .Z(n35343) );
  HS65_LH_IVX2 U19606 ( .A(n35343), .Z(n35344) );
  HS65_LH_IVX2 U19607 ( .A(n35374), .Z(n35345) );
  HS65_LH_IVX2 U19608 ( .A(n35345), .Z(n35346) );
  HS65_LH_IVX2 U19609 ( .A(n35376), .Z(n35347) );
  HS65_LH_IVX2 U19610 ( .A(n35347), .Z(n35348) );
  HS65_LH_IVX2 U19611 ( .A(n35378), .Z(n35349) );
  HS65_LH_IVX2 U19612 ( .A(n35349), .Z(n35350) );
  HS65_LH_IVX2 U19613 ( .A(n35380), .Z(n35351) );
  HS65_LH_IVX2 U19614 ( .A(n35351), .Z(n35352) );
  HS65_LH_IVX2 U19615 ( .A(n35382), .Z(n35353) );
  HS65_LH_IVX2 U19616 ( .A(n35353), .Z(n35354) );
  HS65_LH_IVX2 U19617 ( .A(n35384), .Z(n35355) );
  HS65_LH_IVX2 U19618 ( .A(n35355), .Z(n35356) );
  HS65_LH_IVX2 U19619 ( .A(n35386), .Z(n35357) );
  HS65_LH_IVX2 U19620 ( .A(n35357), .Z(n35358) );
  HS65_LH_IVX2 U19621 ( .A(n35388), .Z(n35359) );
  HS65_LH_IVX2 U19622 ( .A(n35359), .Z(n35360) );
  HS65_LH_IVX2 U19623 ( .A(n35390), .Z(n35361) );
  HS65_LH_IVX2 U19624 ( .A(n35361), .Z(n35362) );
  HS65_LH_BFX2 U19625 ( .A(n35337), .Z(n35363) );
  HS65_LH_BFX2 U19626 ( .A(n35338), .Z(n35364) );
  HS65_LH_BFX2 U19627 ( .A(n35339), .Z(n35365) );
  HS65_LH_BFX2 U19628 ( .A(n35342), .Z(n35366) );
  HS65_LH_IVX2 U19629 ( .A(n35395), .Z(n35367) );
  HS65_LH_IVX2 U19630 ( .A(n35367), .Z(n35368) );
  HS65_LH_IVX2 U19631 ( .A(n35427), .Z(n35369) );
  HS65_LH_IVX2 U19632 ( .A(n35369), .Z(n35370) );
  HS65_LH_IVX2 U19633 ( .A(n35397), .Z(n35371) );
  HS65_LH_IVX2 U19634 ( .A(n35371), .Z(n35372) );
  HS65_LH_IVX2 U19635 ( .A(n35399), .Z(n35373) );
  HS65_LH_IVX2 U19636 ( .A(n35373), .Z(n35374) );
  HS65_LH_IVX2 U19637 ( .A(n35401), .Z(n35375) );
  HS65_LH_IVX2 U19638 ( .A(n35375), .Z(n35376) );
  HS65_LH_IVX2 U19639 ( .A(n35403), .Z(n35377) );
  HS65_LH_IVX2 U19640 ( .A(n35377), .Z(n35378) );
  HS65_LH_IVX2 U19641 ( .A(n35405), .Z(n35379) );
  HS65_LH_IVX2 U19642 ( .A(n35379), .Z(n35380) );
  HS65_LH_IVX2 U19643 ( .A(n35407), .Z(n35381) );
  HS65_LH_IVX2 U19644 ( .A(n35381), .Z(n35382) );
  HS65_LH_IVX2 U19645 ( .A(n35409), .Z(n35383) );
  HS65_LH_IVX2 U19646 ( .A(n35383), .Z(n35384) );
  HS65_LH_IVX2 U19647 ( .A(n35412), .Z(n35385) );
  HS65_LH_IVX2 U19648 ( .A(n35385), .Z(n35386) );
  HS65_LH_IVX2 U19649 ( .A(n35414), .Z(n35387) );
  HS65_LH_IVX2 U19650 ( .A(n35387), .Z(n35388) );
  HS65_LH_IVX2 U19651 ( .A(n35416), .Z(n35389) );
  HS65_LH_IVX2 U19652 ( .A(n35389), .Z(n35390) );
  HS65_LH_BFX2 U19653 ( .A(n35363), .Z(n35391) );
  HS65_LH_BFX2 U19654 ( .A(n35364), .Z(n35392) );
  HS65_LH_BFX2 U19655 ( .A(n35365), .Z(n35393) );
  HS65_LH_IVX2 U19656 ( .A(n35575), .Z(n35394) );
  HS65_LH_IVX2 U19657 ( .A(n35394), .Z(n35395) );
  HS65_LH_IVX2 U19658 ( .A(n35572), .Z(n35396) );
  HS65_LH_IVX2 U19659 ( .A(n35396), .Z(n35397) );
  HS65_LH_IVX2 U19660 ( .A(n35566), .Z(n35398) );
  HS65_LH_IVX2 U19661 ( .A(n35398), .Z(n35399) );
  HS65_LH_IVX2 U19662 ( .A(n35568), .Z(n35400) );
  HS65_LH_IVX2 U19663 ( .A(n35400), .Z(n35401) );
  HS65_LH_IVX2 U19664 ( .A(n35570), .Z(n35402) );
  HS65_LH_IVX2 U19665 ( .A(n35402), .Z(n35403) );
  HS65_LH_IVX2 U19666 ( .A(n35429), .Z(n35404) );
  HS65_LH_IVX2 U19667 ( .A(n35404), .Z(n35405) );
  HS65_LH_IVX2 U19668 ( .A(n35431), .Z(n35406) );
  HS65_LH_IVX2 U19669 ( .A(n35406), .Z(n35407) );
  HS65_LH_IVX2 U19670 ( .A(n35433), .Z(n35408) );
  HS65_LH_IVX2 U19671 ( .A(n35408), .Z(n35409) );
  HS65_LH_BFX2 U19672 ( .A(n35391), .Z(n35410) );
  HS65_LH_IVX2 U19673 ( .A(n35576), .Z(n35411) );
  HS65_LH_IVX2 U19674 ( .A(n35411), .Z(n35412) );
  HS65_LH_IVX2 U19675 ( .A(n35435), .Z(n35413) );
  HS65_LH_IVX2 U19676 ( .A(n35413), .Z(n35414) );
  HS65_LH_IVX2 U19677 ( .A(n35437), .Z(n35415) );
  HS65_LH_IVX2 U19678 ( .A(n35415), .Z(n35416) );
  HS65_LH_BFX2 U19679 ( .A(n35392), .Z(n35417) );
  HS65_LH_IVX2 U19680 ( .A(n35439), .Z(n35418) );
  HS65_LH_IVX2 U19681 ( .A(n35418), .Z(n35419) );
  HS65_LH_BFX2 U19682 ( .A(n35422), .Z(n35420) );
  HS65_LH_IVX2 U19683 ( .A(n35589), .Z(n35421) );
  HS65_LH_IVX2 U19684 ( .A(n35421), .Z(n35422) );
  HS65_LH_BFX2 U19685 ( .A(n35366), .Z(n35423) );
  HS65_LH_IVX2 U19686 ( .A(n35393), .Z(n35424) );
  HS65_LH_IVX2 U19687 ( .A(n35424), .Z(n35425) );
  HS65_LH_IVX2 U19688 ( .A(n35452), .Z(n35426) );
  HS65_LH_IVX2 U19689 ( .A(n35426), .Z(n35427) );
  HS65_LH_IVX2 U19690 ( .A(n35441), .Z(n35428) );
  HS65_LH_IVX2 U19691 ( .A(n35428), .Z(n35429) );
  HS65_LH_IVX2 U19692 ( .A(n35443), .Z(n35430) );
  HS65_LH_IVX2 U19693 ( .A(n35430), .Z(n35431) );
  HS65_LH_IVX2 U19694 ( .A(n35445), .Z(n35432) );
  HS65_LH_IVX2 U19695 ( .A(n35432), .Z(n35433) );
  HS65_LH_IVX2 U19696 ( .A(n35447), .Z(n35434) );
  HS65_LH_IVX2 U19697 ( .A(n35434), .Z(n35435) );
  HS65_LH_IVX2 U19698 ( .A(n35449), .Z(n35436) );
  HS65_LH_IVX2 U19699 ( .A(n35436), .Z(n35437) );
  HS65_LH_IVX2 U19700 ( .A(n35451), .Z(n35438) );
  HS65_LH_IVX2 U19701 ( .A(n35438), .Z(n35439) );
  HS65_LH_IVX2 U19702 ( .A(n35454), .Z(n35440) );
  HS65_LH_IVX2 U19703 ( .A(n35440), .Z(n35441) );
  HS65_LH_IVX2 U19704 ( .A(n35456), .Z(n35442) );
  HS65_LH_IVX2 U19705 ( .A(n35442), .Z(n35443) );
  HS65_LH_IVX2 U19706 ( .A(n35458), .Z(n35444) );
  HS65_LH_IVX2 U19707 ( .A(n35444), .Z(n35445) );
  HS65_LH_IVX2 U19708 ( .A(n35460), .Z(n35446) );
  HS65_LH_IVX2 U19709 ( .A(n35446), .Z(n35447) );
  HS65_LH_IVX2 U19710 ( .A(n35462), .Z(n35448) );
  HS65_LH_IVX2 U19711 ( .A(n35448), .Z(n35449) );
  HS65_LH_IVX2 U19712 ( .A(n35464), .Z(n35450) );
  HS65_LH_IVX2 U19713 ( .A(n35450), .Z(n35451) );
  HS65_LH_BFX2 U19714 ( .A(n35515), .Z(n35452) );
  HS65_LH_IVX2 U19715 ( .A(n35477), .Z(n35453) );
  HS65_LH_IVX2 U19716 ( .A(n35453), .Z(n35454) );
  HS65_LH_IVX2 U19717 ( .A(n35467), .Z(n35455) );
  HS65_LH_IVX2 U19718 ( .A(n35455), .Z(n35456) );
  HS65_LH_IVX2 U19719 ( .A(n35469), .Z(n35457) );
  HS65_LH_IVX2 U19720 ( .A(n35457), .Z(n35458) );
  HS65_LH_IVX2 U19721 ( .A(n35471), .Z(n35459) );
  HS65_LH_IVX2 U19722 ( .A(n35459), .Z(n35460) );
  HS65_LH_IVX2 U19723 ( .A(n35473), .Z(n35461) );
  HS65_LH_IVX2 U19724 ( .A(n35461), .Z(n35462) );
  HS65_LH_IVX2 U19725 ( .A(n35476), .Z(n35463) );
  HS65_LH_IVX2 U19726 ( .A(n35463), .Z(n35464) );
  HS65_LH_BFX2 U19727 ( .A(n35423), .Z(n35465) );
  HS65_LH_IVX2 U19728 ( .A(n35479), .Z(n35466) );
  HS65_LH_IVX2 U19729 ( .A(n35466), .Z(n35467) );
  HS65_LH_IVX2 U19730 ( .A(n35481), .Z(n35468) );
  HS65_LH_IVX2 U19731 ( .A(n35468), .Z(n35469) );
  HS65_LH_IVX2 U19732 ( .A(n35483), .Z(n35470) );
  HS65_LH_IVX2 U19733 ( .A(n35470), .Z(n35471) );
  HS65_LH_IVX2 U19734 ( .A(n35486), .Z(n35472) );
  HS65_LH_IVX2 U19735 ( .A(n35472), .Z(n35473) );
  HS65_LH_BFX2 U19736 ( .A(n35465), .Z(n35474) );
  HS65_LH_IVX2 U19737 ( .A(n35488), .Z(n35475) );
  HS65_LH_IVX2 U19738 ( .A(n35475), .Z(n35476) );
  HS65_LH_BFX2 U19739 ( .A(n35489), .Z(n35477) );
  HS65_LH_IVX2 U19740 ( .A(n35498), .Z(n35478) );
  HS65_LH_IVX2 U19741 ( .A(n35478), .Z(n35479) );
  HS65_LH_IVX2 U19742 ( .A(n35499), .Z(n35480) );
  HS65_LH_IVX2 U19743 ( .A(n35480), .Z(n35481) );
  HS65_LH_IVX2 U19744 ( .A(n35492), .Z(n35482) );
  HS65_LH_IVX2 U19745 ( .A(n35482), .Z(n35483) );
  HS65_LH_BFX2 U19746 ( .A(n35474), .Z(n35484) );
  HS65_LH_IVX2 U19747 ( .A(n35494), .Z(n35485) );
  HS65_LH_IVX2 U19748 ( .A(n35485), .Z(n35486) );
  HS65_LH_IVX2 U19749 ( .A(n35496), .Z(n35487) );
  HS65_LH_IVX2 U19750 ( .A(n35487), .Z(n35488) );
  HS65_LH_BFX2 U19751 ( .A(n35497), .Z(n35489) );
  HS65_LH_BFX2 U19752 ( .A(n35484), .Z(n35490) );
  HS65_LH_IVX2 U19753 ( .A(n35504), .Z(n35491) );
  HS65_LH_IVX2 U19754 ( .A(n35491), .Z(n35492) );
  HS65_LH_IVX2 U19755 ( .A(n35506), .Z(n35493) );
  HS65_LH_IVX2 U19756 ( .A(n35493), .Z(n35494) );
  HS65_LH_IVX2 U19757 ( .A(n35508), .Z(n35495) );
  HS65_LH_IVX2 U19758 ( .A(n35495), .Z(n35496) );
  HS65_LH_BFX2 U19759 ( .A(n35509), .Z(n35497) );
  HS65_LH_BFX2 U19760 ( .A(n35510), .Z(n35498) );
  HS65_LH_BFX2 U19761 ( .A(n35502), .Z(n35499) );
  HS65_LH_BFX2 U19762 ( .A(n35490), .Z(n35500) );
  HS65_LH_IVX2 U19763 ( .A(n35523), .Z(n35501) );
  HS65_LH_IVX2 U19764 ( .A(n35501), .Z(n35502) );
  HS65_LH_IVX2 U19765 ( .A(n35517), .Z(n35503) );
  HS65_LH_IVX2 U19766 ( .A(n35503), .Z(n35504) );
  HS65_LH_IVX2 U19767 ( .A(n35519), .Z(n35505) );
  HS65_LH_IVX2 U19768 ( .A(n35505), .Z(n35506) );
  HS65_LH_IVX2 U19769 ( .A(n35538), .Z(n35507) );
  HS65_LH_IVX2 U19770 ( .A(n35507), .Z(n35508) );
  HS65_LH_BFX2 U19771 ( .A(n35524), .Z(n35509) );
  HS65_LH_BFX2 U19772 ( .A(n35513), .Z(n35510) );
  HS65_LH_BFX2 U19773 ( .A(n35500), .Z(n35511) );
  HS65_LH_IVX2 U19774 ( .A(n35526), .Z(n35512) );
  HS65_LH_IVX2 U19775 ( .A(n35512), .Z(n35513) );
  HS65_LH_IVX2 U19776 ( .A(n35533), .Z(n35514) );
  HS65_LH_IVX2 U19777 ( .A(n35514), .Z(n35515) );
  HS65_LH_IVX2 U19778 ( .A(n35529), .Z(n35516) );
  HS65_LH_IVX2 U19779 ( .A(n35516), .Z(n35517) );
  HS65_LH_IVX2 U19780 ( .A(n35531), .Z(n35518) );
  HS65_LH_IVX2 U19781 ( .A(n35518), .Z(n35519) );
  HS65_LH_IVX2 U19782 ( .A(n35520), .Z(n35521) );
  HS65_LH_IVX2 U19783 ( .A(n35522), .Z(n35523) );
  HS65_LH_BFX2 U19784 ( .A(n35532), .Z(n35524) );
  HS65_LH_IVX2 U19785 ( .A(n17511), .Z(n35525) );
  HS65_LH_IVX2 U19786 ( .A(n35525), .Z(n35526) );
  HS65_LH_BFX2 U19787 ( .A(n35417), .Z(n35527) );
  HS65_LH_IVX2 U19788 ( .A(n35536), .Z(n35528) );
  HS65_LH_IVX2 U19789 ( .A(n35528), .Z(n35529) );
  HS65_LH_IVX2 U19790 ( .A(n195), .Z(n35530) );
  HS65_LH_IVX2 U19791 ( .A(n35530), .Z(n35531) );
  HS65_LH_BFX2 U19792 ( .A(n35539), .Z(n35532) );
  HS65_LH_BFX2 U19793 ( .A(n35540), .Z(n35533) );
  HS65_LH_BFX2 U19794 ( .A(n35527), .Z(n35534) );
  HS65_LH_IVX2 U19795 ( .A(n35542), .Z(n35535) );
  HS65_LH_IVX2 U19796 ( .A(n35535), .Z(n35536) );
  HS65_LH_IVX2 U19797 ( .A(n35534), .Z(n35537) );
  HS65_LH_IVX2 U19798 ( .A(n35537), .Z(n35538) );
  HS65_LH_BFX2 U19799 ( .A(n35541), .Z(n35539) );
  HS65_LH_BFX2 U19800 ( .A(n35511), .Z(n35540) );
  HS65_LH_BFX2 U19801 ( .A(n35543), .Z(n35541) );
  HS65_LH_BFX2 U19802 ( .A(n17300), .Z(n35542) );
  HS65_LH_BFX2 U19803 ( .A(n17512), .Z(n35543) );
  HS65_LH_BFX2 U19804 ( .A(n35545), .Z(n35544) );
  HS65_LH_BFX2 U19805 ( .A(n35546), .Z(n35545) );
  HS65_LH_BFX2 U19806 ( .A(n35547), .Z(n35546) );
  HS65_LH_BFX2 U19807 ( .A(n35548), .Z(n35547) );
  HS65_LH_BFX2 U19808 ( .A(n35549), .Z(n35548) );
  HS65_LH_BFX2 U19809 ( .A(n35550), .Z(n35549) );
  HS65_LH_BFX2 U19810 ( .A(n35551), .Z(n35550) );
  HS65_LH_BFX2 U19811 ( .A(n35552), .Z(n35551) );
  HS65_LH_BFX2 U19812 ( .A(n35553), .Z(n35552) );
  HS65_LH_BFX2 U19813 ( .A(n35554), .Z(n35553) );
  HS65_LH_BFX2 U19814 ( .A(n35555), .Z(n35554) );
  HS65_LH_BFX2 U19815 ( .A(n35556), .Z(n35555) );
  HS65_LH_BFX2 U19816 ( .A(n35557), .Z(n35556) );
  HS65_LH_BFX2 U19817 ( .A(n35558), .Z(n35557) );
  HS65_LH_BFX2 U19818 ( .A(n35559), .Z(n35558) );
  HS65_LH_BFX2 U19819 ( .A(n35560), .Z(n35559) );
  HS65_LH_BFX2 U19820 ( .A(n35561), .Z(n35560) );
  HS65_LH_BFX2 U19821 ( .A(n14538), .Z(n35561) );
  HS65_LH_BFX2 U19822 ( .A(n17604), .Z(n35562) );
  HS65_LH_IVX2 U19823 ( .A(n35590), .Z(n35563) );
  HS65_LH_IVX2 U19824 ( .A(n35563), .Z(n35564) );
  HS65_LH_IVX2 U19825 ( .A(n35579), .Z(n35565) );
  HS65_LH_IVX2 U19826 ( .A(n35565), .Z(n35566) );
  HS65_LH_IVX2 U19827 ( .A(n35583), .Z(n35567) );
  HS65_LH_IVX2 U19828 ( .A(n35567), .Z(n35568) );
  HS65_LH_IVX2 U19829 ( .A(n35581), .Z(n35569) );
  HS65_LH_IVX2 U19830 ( .A(n35569), .Z(n35570) );
  HS65_LH_IVX2 U19831 ( .A(n35585), .Z(n35571) );
  HS65_LH_IVX2 U19832 ( .A(n35571), .Z(n35572) );
  HS65_LH_BFX2 U19833 ( .A(n35410), .Z(n35573) );
  HS65_LH_BFX2 U19834 ( .A(n35586), .Z(n35574) );
  HS65_LH_BFX2 U19835 ( .A(n35587), .Z(n35575) );
  HS65_LH_BFX2 U19836 ( .A(n35591), .Z(n35576) );
  HS65_LH_BFX2 U19837 ( .A(n35573), .Z(n35577) );
  HS65_LH_IVX2 U19838 ( .A(n35594), .Z(n35578) );
  HS65_LH_IVX2 U19839 ( .A(n35578), .Z(n35579) );
  HS65_LH_IVX2 U19840 ( .A(n35596), .Z(n35580) );
  HS65_LH_IVX2 U19841 ( .A(n35580), .Z(n35581) );
  HS65_LH_IVX2 U19842 ( .A(n35598), .Z(n35582) );
  HS65_LH_IVX2 U19843 ( .A(n35582), .Z(n35583) );
  HS65_LH_IVX2 U19844 ( .A(n35600), .Z(n35584) );
  HS65_LH_IVX2 U19845 ( .A(n35584), .Z(n35585) );
  HS65_LH_BFX2 U19846 ( .A(n35601), .Z(n35586) );
  HS65_LH_BFX2 U19847 ( .A(n35602), .Z(n35587) );
  HS65_LH_IVX2 U19848 ( .A(n35604), .Z(n35588) );
  HS65_LH_IVX2 U19849 ( .A(n35588), .Z(n35589) );
  HS65_LH_BFX2 U19850 ( .A(n35605), .Z(n35590) );
  HS65_LH_BFX2 U19851 ( .A(n35606), .Z(n35591) );
  HS65_LH_BFX2 U19852 ( .A(n35577), .Z(n35592) );
  HS65_LH_IVX2 U19853 ( .A(n35611), .Z(n35593) );
  HS65_LH_IVX2 U19854 ( .A(n35593), .Z(n35594) );
  HS65_LH_IVX2 U19855 ( .A(n35613), .Z(n35595) );
  HS65_LH_IVX2 U19856 ( .A(n35595), .Z(n35596) );
  HS65_LH_IVX2 U19857 ( .A(n35615), .Z(n35597) );
  HS65_LH_IVX2 U19858 ( .A(n35597), .Z(n35598) );
  HS65_LH_IVX2 U19859 ( .A(n35617), .Z(n35599) );
  HS65_LH_IVX2 U19860 ( .A(n35599), .Z(n35600) );
  HS65_LH_BFX2 U19861 ( .A(n35618), .Z(n35601) );
  HS65_LH_BFX2 U19862 ( .A(n35619), .Z(n35602) );
  HS65_LH_IVX2 U19863 ( .A(n35650), .Z(n35603) );
  HS65_LH_IVX2 U19864 ( .A(n35603), .Z(n35604) );
  HS65_LH_BFX2 U19865 ( .A(n35608), .Z(n35605) );
  HS65_LH_BFX2 U19866 ( .A(n35620), .Z(n35606) );
  HS65_LH_IVX2 U19867 ( .A(n35623), .Z(n35607) );
  HS65_LH_IVX2 U19868 ( .A(n35607), .Z(n35608) );
  HS65_LH_BFX2 U19869 ( .A(n35592), .Z(n35609) );
  HS65_LH_IVX2 U19870 ( .A(n35625), .Z(n35610) );
  HS65_LH_IVX2 U19871 ( .A(n35610), .Z(n35611) );
  HS65_LH_IVX2 U19872 ( .A(n35627), .Z(n35612) );
  HS65_LH_IVX2 U19873 ( .A(n35612), .Z(n35613) );
  HS65_LH_IVX2 U19874 ( .A(n35629), .Z(n35614) );
  HS65_LH_IVX2 U19875 ( .A(n35614), .Z(n35615) );
  HS65_LH_IVX2 U19876 ( .A(n35631), .Z(n35616) );
  HS65_LH_IVX2 U19877 ( .A(n35616), .Z(n35617) );
  HS65_LH_BFX2 U19878 ( .A(n35632), .Z(n35618) );
  HS65_LH_BFX2 U19879 ( .A(n35633), .Z(n35619) );
  HS65_LH_BFX2 U19880 ( .A(n35637), .Z(n35620) );
  HS65_LH_BFX2 U19881 ( .A(n35609), .Z(n35621) );
  HS65_LH_IVX2 U19882 ( .A(n35640), .Z(n35622) );
  HS65_LH_IVX2 U19883 ( .A(n35622), .Z(n35623) );
  HS65_LH_IVX2 U19884 ( .A(n35642), .Z(n35624) );
  HS65_LH_IVX2 U19885 ( .A(n35624), .Z(n35625) );
  HS65_LH_IVX2 U19886 ( .A(n17316), .Z(n35626) );
  HS65_LH_IVX2 U19887 ( .A(n35626), .Z(n35627) );
  HS65_LH_IVX2 U19888 ( .A(n35657), .Z(n35628) );
  HS65_LH_IVX2 U19889 ( .A(n35628), .Z(n35629) );
  HS65_LH_IVX2 U19890 ( .A(n35644), .Z(n35630) );
  HS65_LH_IVX2 U19891 ( .A(n35630), .Z(n35631) );
  HS65_LH_BFX2 U19892 ( .A(n35635), .Z(n35632) );
  HS65_LH_BFX2 U19893 ( .A(n35645), .Z(n35633) );
  HS65_LH_IVX2 U19894 ( .A(n35647), .Z(n35634) );
  HS65_LH_IVX2 U19895 ( .A(n35634), .Z(n35635) );
  HS65_LH_BFX2 U19896 ( .A(n17632), .Z(n35636) );
  HS65_LH_BFX2 U19897 ( .A(n35651), .Z(n35637) );
  HS65_LH_BFX2 U19898 ( .A(n35621), .Z(n35638) );
  HS65_LH_IVX2 U19899 ( .A(n35656), .Z(n35639) );
  HS65_LH_IVX2 U19900 ( .A(n35639), .Z(n35640) );
  HS65_LH_IVX2 U19901 ( .A(n17785), .Z(n35641) );
  HS65_LH_IVX2 U19902 ( .A(n35641), .Z(n35642) );
  HS65_LH_IVX2 U19903 ( .A(n35660), .Z(n35643) );
  HS65_LH_IVX2 U19904 ( .A(n35643), .Z(n35644) );
  HS65_LH_BFX2 U19905 ( .A(n35658), .Z(n35645) );
  HS65_LH_IVX2 U19906 ( .A(n35662), .Z(n35646) );
  HS65_LH_IVX2 U19907 ( .A(n35646), .Z(n35647) );
  HS65_LH_BFX2 U19908 ( .A(n35636), .Z(n35648) );
  HS65_LH_IVX2 U19909 ( .A(n35648), .Z(n35649) );
  HS65_LH_IVX2 U19910 ( .A(n35649), .Z(n35650) );
  HS65_LH_BFX2 U19911 ( .A(n35663), .Z(n35651) );
  HS65_LH_BFX2 U19912 ( .A(n35638), .Z(n35652) );
  HS65_LH_IVX2 U19913 ( .A(n35652), .Z(n35653) );
  HS65_LH_IVX2 U19914 ( .A(n35653), .Z(n35654) );
  HS65_LH_IVX2 U19915 ( .A(n35666), .Z(n35655) );
  HS65_LH_IVX2 U19916 ( .A(n35655), .Z(n35656) );
  HS65_LH_BFX2 U19917 ( .A(n35664), .Z(n35657) );
  HS65_LH_BFX2 U19918 ( .A(n35667), .Z(n35658) );
  HS65_LH_IVX2 U19919 ( .A(n35261), .Z(n35659) );
  HS65_LH_IVX2 U19920 ( .A(n35659), .Z(n35660) );
  HS65_LH_IVX2 U19921 ( .A(n35668), .Z(n35661) );
  HS65_LH_IVX2 U19922 ( .A(n35661), .Z(n35662) );
  HS65_LH_BFX2 U19923 ( .A(n31197), .Z(n35663) );
  HS65_LH_BFX2 U19924 ( .A(n17788), .Z(n35664) );
  HS65_LH_IVX2 U19925 ( .A(n40991), .Z(n35665) );
  HS65_LH_IVX2 U19926 ( .A(n35665), .Z(n35666) );
  HS65_LH_BFX2 U19927 ( .A(n17436), .Z(n35667) );
  HS65_LH_BFX2 U19928 ( .A(n270), .Z(n35668) );
  HS65_LH_IVX2 U19929 ( .A(n35696), .Z(n35669) );
  HS65_LH_IVX2 U19930 ( .A(n35669), .Z(n35670) );
  HS65_LH_NAND2X2 U19931 ( .A(n15817), .B(n15816), .Z(n15825) );
  HS65_LH_BFX2 U19932 ( .A(n15825), .Z(n35671) );
  HS65_LH_BFX2 U19933 ( .A(n35674), .Z(n35672) );
  HS65_LH_BFX2 U19934 ( .A(n2645), .Z(n35673) );
  HS65_LH_BFX2 U19935 ( .A(n35676), .Z(n35674) );
  HS65_LH_BFX2 U19936 ( .A(n35673), .Z(n35675) );
  HS65_LH_BFX2 U19937 ( .A(n35678), .Z(n35676) );
  HS65_LH_BFX2 U19938 ( .A(n35675), .Z(n35677) );
  HS65_LH_BFX2 U19939 ( .A(n35680), .Z(n35678) );
  HS65_LH_BFX2 U19940 ( .A(n35677), .Z(n35679) );
  HS65_LH_BFX2 U19941 ( .A(n35682), .Z(n35680) );
  HS65_LH_BFX2 U19942 ( .A(n35679), .Z(n35681) );
  HS65_LH_BFX2 U19943 ( .A(n35684), .Z(n35682) );
  HS65_LH_BFX2 U19944 ( .A(n35681), .Z(n35683) );
  HS65_LH_BFX2 U19945 ( .A(n35686), .Z(n35684) );
  HS65_LH_BFX2 U19946 ( .A(n35683), .Z(n35685) );
  HS65_LH_BFX2 U19947 ( .A(n35688), .Z(n35686) );
  HS65_LH_BFX2 U19948 ( .A(n35685), .Z(n35687) );
  HS65_LH_BFX2 U19949 ( .A(n35690), .Z(n35688) );
  HS65_LH_BFX2 U19950 ( .A(n35687), .Z(n35689) );
  HS65_LH_BFX2 U19951 ( .A(n35692), .Z(n35690) );
  HS65_LH_BFX2 U19952 ( .A(n35689), .Z(n35691) );
  HS65_LH_BFX2 U19953 ( .A(n35694), .Z(n35692) );
  HS65_LH_BFX2 U19954 ( .A(n35691), .Z(n35693) );
  HS65_LH_BFX2 U19955 ( .A(n35697), .Z(n35694) );
  HS65_LH_IVX2 U19956 ( .A(n15824), .Z(n35695) );
  HS65_LH_IVX2 U19957 ( .A(n35695), .Z(n35696) );
  HS65_LH_BFX2 U19958 ( .A(n35700), .Z(n35697) );
  HS65_LH_BFX2 U19959 ( .A(n36045), .Z(n35698) );
  HS65_LH_IVX2 U19960 ( .A(n2646), .Z(n35699) );
  HS65_LH_IVX2 U19961 ( .A(n35699), .Z(n35700) );
  HS65_LH_IVX2 U19962 ( .A(n35693), .Z(n35701) );
  HS65_LH_IVX2 U19963 ( .A(n35701), .Z(n35702) );
  HS65_LH_BFX2 U19964 ( .A(n35734), .Z(n35703) );
  HS65_LH_BFX2 U19965 ( .A(n37854), .Z(n35704) );
  HS65_LH_BFX2 U19966 ( .A(n35707), .Z(n35705) );
  HS65_LH_BFX2 U19967 ( .A(n2045), .Z(n35706) );
  HS65_LH_BFX2 U19968 ( .A(n35709), .Z(n35707) );
  HS65_LH_BFX2 U19969 ( .A(n35706), .Z(n35708) );
  HS65_LH_BFX2 U19970 ( .A(n35711), .Z(n35709) );
  HS65_LH_BFX2 U19971 ( .A(n35708), .Z(n35710) );
  HS65_LH_BFX2 U19972 ( .A(n35713), .Z(n35711) );
  HS65_LH_BFX2 U19973 ( .A(n35710), .Z(n35712) );
  HS65_LH_BFX2 U19974 ( .A(n35715), .Z(n35713) );
  HS65_LH_BFX2 U19975 ( .A(n35712), .Z(n35714) );
  HS65_LH_BFX2 U19976 ( .A(n35717), .Z(n35715) );
  HS65_LH_BFX2 U19977 ( .A(n35714), .Z(n35716) );
  HS65_LH_BFX2 U19978 ( .A(n35719), .Z(n35717) );
  HS65_LH_BFX2 U19979 ( .A(n35716), .Z(n35718) );
  HS65_LH_BFX2 U19980 ( .A(n35721), .Z(n35719) );
  HS65_LH_BFX2 U19981 ( .A(n35718), .Z(n35720) );
  HS65_LH_BFX2 U19982 ( .A(n35723), .Z(n35721) );
  HS65_LH_BFX2 U19983 ( .A(n35720), .Z(n35722) );
  HS65_LH_BFX2 U19984 ( .A(n35725), .Z(n35723) );
  HS65_LH_BFX2 U19985 ( .A(n35722), .Z(n35724) );
  HS65_LH_BFX2 U19986 ( .A(n35727), .Z(n35725) );
  HS65_LH_BFX2 U19987 ( .A(n35724), .Z(n35726) );
  HS65_LH_BFX2 U19988 ( .A(n35729), .Z(n35727) );
  HS65_LH_BFX2 U19989 ( .A(n35726), .Z(n35728) );
  HS65_LH_BFX2 U19990 ( .A(n35731), .Z(n35729) );
  HS65_LH_BFX2 U19991 ( .A(n35728), .Z(n35730) );
  HS65_LH_BFX2 U19992 ( .A(n35735), .Z(n35731) );
  HS65_LH_BFX2 U19993 ( .A(n16326), .Z(n35732) );
  HS65_LH_IVX2 U19994 ( .A(n35730), .Z(n35733) );
  HS65_LH_IVX2 U19995 ( .A(n35733), .Z(n35734) );
  HS65_LH_BFX2 U19996 ( .A(n2046), .Z(n35735) );
  HS65_LH_BFX2 U19997 ( .A(n35739), .Z(n35736) );
  HS65_LH_BFX2 U19998 ( .A(n35741), .Z(n35737) );
  HS65_LH_IVX2 U19999 ( .A(n35745), .Z(n35738) );
  HS65_LH_IVX2 U20000 ( .A(n35738), .Z(n35739) );
  HS65_LH_IVX2 U20001 ( .A(n35747), .Z(n35740) );
  HS65_LH_IVX2 U20002 ( .A(n35740), .Z(n35741) );
  HS65_LH_BFX2 U20003 ( .A(n35749), .Z(n35742) );
  HS65_LH_BFX2 U20004 ( .A(n2550), .Z(n35743) );
  HS65_LH_IVX2 U20005 ( .A(n35751), .Z(n35744) );
  HS65_LH_IVX2 U20006 ( .A(n35744), .Z(n35745) );
  HS65_LH_IVX2 U20007 ( .A(n35753), .Z(n35746) );
  HS65_LH_IVX2 U20008 ( .A(n35746), .Z(n35747) );
  HS65_LH_IVX2 U20009 ( .A(n35755), .Z(n35748) );
  HS65_LH_IVX2 U20010 ( .A(n35748), .Z(n35749) );
  HS65_LH_IVX2 U20011 ( .A(n35757), .Z(n35750) );
  HS65_LH_IVX2 U20012 ( .A(n35750), .Z(n35751) );
  HS65_LH_IVX2 U20013 ( .A(n35759), .Z(n35752) );
  HS65_LH_IVX2 U20014 ( .A(n35752), .Z(n35753) );
  HS65_LH_IVX2 U20015 ( .A(n35761), .Z(n35754) );
  HS65_LH_IVX2 U20016 ( .A(n35754), .Z(n35755) );
  HS65_LH_IVX2 U20017 ( .A(n35766), .Z(n35756) );
  HS65_LH_IVX2 U20018 ( .A(n35756), .Z(n35757) );
  HS65_LH_IVX2 U20019 ( .A(n35763), .Z(n35758) );
  HS65_LH_IVX2 U20020 ( .A(n35758), .Z(n35759) );
  HS65_LH_IVX2 U20021 ( .A(n35765), .Z(n35760) );
  HS65_LH_IVX2 U20022 ( .A(n35760), .Z(n35761) );
  HS65_LH_IVX2 U20023 ( .A(n35768), .Z(n35762) );
  HS65_LH_IVX2 U20024 ( .A(n35762), .Z(n35763) );
  HS65_LH_IVX2 U20025 ( .A(n35770), .Z(n35764) );
  HS65_LH_IVX2 U20026 ( .A(n35764), .Z(n35765) );
  HS65_LH_BFX2 U20027 ( .A(n35771), .Z(n35766) );
  HS65_LH_IVX2 U20028 ( .A(n35773), .Z(n35767) );
  HS65_LH_IVX2 U20029 ( .A(n35767), .Z(n35768) );
  HS65_LH_IVX2 U20030 ( .A(n35775), .Z(n35769) );
  HS65_LH_IVX2 U20031 ( .A(n35769), .Z(n35770) );
  HS65_LH_BFX2 U20032 ( .A(n35776), .Z(n35771) );
  HS65_LH_IVX2 U20033 ( .A(n35778), .Z(n35772) );
  HS65_LH_IVX2 U20034 ( .A(n35772), .Z(n35773) );
  HS65_LH_IVX2 U20035 ( .A(n35780), .Z(n35774) );
  HS65_LH_IVX2 U20036 ( .A(n35774), .Z(n35775) );
  HS65_LH_BFX2 U20037 ( .A(n35781), .Z(n35776) );
  HS65_LH_IVX2 U20038 ( .A(n35785), .Z(n35777) );
  HS65_LH_IVX2 U20039 ( .A(n35777), .Z(n35778) );
  HS65_LH_IVX2 U20040 ( .A(n35783), .Z(n35779) );
  HS65_LH_IVX2 U20041 ( .A(n35779), .Z(n35780) );
  HS65_LH_BFX2 U20042 ( .A(n35784), .Z(n35781) );
  HS65_LH_IVX2 U20043 ( .A(n35788), .Z(n35782) );
  HS65_LH_IVX2 U20044 ( .A(n35782), .Z(n35783) );
  HS65_LH_BFX2 U20045 ( .A(n35790), .Z(n35784) );
  HS65_LH_BFX2 U20046 ( .A(n35792), .Z(n35785) );
  HS65_LH_IVX2 U20047 ( .A(n35798), .Z(n35787) );
  HS65_LH_IVX2 U20048 ( .A(n35787), .Z(n35788) );
  HS65_LH_BFX2 U20049 ( .A(n35795), .Z(n35789) );
  HS65_LH_BFX2 U20050 ( .A(n35794), .Z(n35790) );
  HS65_LH_IVX2 U20051 ( .A(n2549), .Z(n35791) );
  HS65_LH_IVX2 U20052 ( .A(n35791), .Z(n35792) );
  HS65_LH_IVX2 U20053 ( .A(n35797), .Z(n35793) );
  HS65_LH_IVX2 U20054 ( .A(n35793), .Z(n35794) );
  HS65_LH_BFX2 U20055 ( .A(n15905), .Z(n35795) );
  HS65_LH_IVX2 U20056 ( .A(n35800), .Z(n35796) );
  HS65_LH_IVX2 U20057 ( .A(n35796), .Z(n35797) );
  HS65_LH_BFX2 U20058 ( .A(n35801), .Z(n35798) );
  HS65_LH_IVX2 U20059 ( .A(n35803), .Z(n35799) );
  HS65_LH_IVX2 U20060 ( .A(n35799), .Z(n35800) );
  HS65_LH_BFX2 U20061 ( .A(n35743), .Z(n35801) );
  HS65_LH_BFX2 U20062 ( .A(n15907), .Z(n35802) );
  HS65_LH_BFX2 U20063 ( .A(n35804), .Z(n35803) );
  HS65_LH_BFX2 U20064 ( .A(n35805), .Z(n35804) );
  HS65_LH_BFX2 U20065 ( .A(n35806), .Z(n35805) );
  HS65_LH_BFX2 U20066 ( .A(n35807), .Z(n35806) );
  HS65_LH_BFX2 U20067 ( .A(n35808), .Z(n35807) );
  HS65_LH_BFX2 U20068 ( .A(n17868), .Z(n35808) );
  HS65_LH_IVX2 U20069 ( .A(n37261), .Z(n35809) );
  HS65_LH_IVX2 U20070 ( .A(n35809), .Z(n35810) );
  HS65_LH_BFX2 U20071 ( .A(n2310), .Z(n35811) );
  HS65_LH_IVX2 U20072 ( .A(n35816), .Z(n35812) );
  HS65_LH_IVX2 U20073 ( .A(n35812), .Z(n35813) );
  HS65_LH_BFX2 U20074 ( .A(n35815), .Z(n35814) );
  HS65_LH_BFX2 U20075 ( .A(n35817), .Z(n35815) );
  HS65_LH_BFX2 U20076 ( .A(n35818), .Z(n35816) );
  HS65_LH_BFX2 U20077 ( .A(n35819), .Z(n35817) );
  HS65_LH_BFX2 U20078 ( .A(n35820), .Z(n35818) );
  HS65_LH_BFX2 U20079 ( .A(n35821), .Z(n35819) );
  HS65_LH_BFX2 U20080 ( .A(n35822), .Z(n35820) );
  HS65_LH_BFX2 U20081 ( .A(n35823), .Z(n35821) );
  HS65_LH_BFX2 U20082 ( .A(n35824), .Z(n35822) );
  HS65_LH_BFX2 U20083 ( .A(n35825), .Z(n35823) );
  HS65_LH_BFX2 U20084 ( .A(n35826), .Z(n35824) );
  HS65_LH_BFX2 U20085 ( .A(n35827), .Z(n35825) );
  HS65_LH_BFX2 U20086 ( .A(n35828), .Z(n35826) );
  HS65_LH_BFX2 U20087 ( .A(n35829), .Z(n35827) );
  HS65_LH_BFX2 U20088 ( .A(n35830), .Z(n35828) );
  HS65_LH_BFX2 U20089 ( .A(n35831), .Z(n35829) );
  HS65_LH_BFX2 U20090 ( .A(n35832), .Z(n35830) );
  HS65_LH_BFX2 U20091 ( .A(n35833), .Z(n35831) );
  HS65_LH_BFX2 U20092 ( .A(n35834), .Z(n35832) );
  HS65_LH_BFX2 U20093 ( .A(n35835), .Z(n35833) );
  HS65_LH_BFX2 U20094 ( .A(n35836), .Z(n35834) );
  HS65_LH_BFX2 U20095 ( .A(n35837), .Z(n35835) );
  HS65_LH_BFX2 U20096 ( .A(n35838), .Z(n35836) );
  HS65_LH_BFX2 U20097 ( .A(n35841), .Z(n35837) );
  HS65_LH_BFX2 U20098 ( .A(n35840), .Z(n35838) );
  HS65_LH_BFX2 U20099 ( .A(n16105), .Z(n35839) );
  HS65_LH_BFX2 U20100 ( .A(n35842), .Z(n35840) );
  HS65_LH_BFX2 U20101 ( .A(n2309), .Z(n35841) );
  HS65_LH_BFX2 U20102 ( .A(n35811), .Z(n35842) );
  HS65_LH_BFX2 U20103 ( .A(n35848), .Z(n35843) );
  HS65_LH_BFX2 U20104 ( .A(n37804), .Z(n35844) );
  HS65_LH_BFX2 U20105 ( .A(n35847), .Z(n35845) );
  HS65_LH_IVX2 U20106 ( .A(n35850), .Z(n35846) );
  HS65_LH_IVX2 U20107 ( .A(n35846), .Z(n35847) );
  HS65_LH_BFX2 U20108 ( .A(n35849), .Z(n35848) );
  HS65_LH_BFX2 U20109 ( .A(n35851), .Z(n35849) );
  HS65_LH_BFX2 U20110 ( .A(n35852), .Z(n35850) );
  HS65_LH_BFX2 U20111 ( .A(n35853), .Z(n35851) );
  HS65_LH_BFX2 U20112 ( .A(n35854), .Z(n35852) );
  HS65_LH_BFX2 U20113 ( .A(n35855), .Z(n35853) );
  HS65_LH_BFX2 U20114 ( .A(n35856), .Z(n35854) );
  HS65_LH_BFX2 U20115 ( .A(n35857), .Z(n35855) );
  HS65_LH_BFX2 U20116 ( .A(n35858), .Z(n35856) );
  HS65_LH_BFX2 U20117 ( .A(n35859), .Z(n35857) );
  HS65_LH_BFX2 U20118 ( .A(n35860), .Z(n35858) );
  HS65_LH_BFX2 U20119 ( .A(n35861), .Z(n35859) );
  HS65_LH_BFX2 U20120 ( .A(n35862), .Z(n35860) );
  HS65_LH_BFX2 U20121 ( .A(n35863), .Z(n35861) );
  HS65_LH_BFX2 U20122 ( .A(n35864), .Z(n35862) );
  HS65_LH_BFX2 U20123 ( .A(n35865), .Z(n35863) );
  HS65_LH_BFX2 U20124 ( .A(n35866), .Z(n35864) );
  HS65_LH_BFX2 U20125 ( .A(n35867), .Z(n35865) );
  HS65_LH_BFX2 U20126 ( .A(n35868), .Z(n35866) );
  HS65_LH_BFX2 U20127 ( .A(n35869), .Z(n35867) );
  HS65_LH_BFX2 U20128 ( .A(n35870), .Z(n35868) );
  HS65_LH_BFX2 U20129 ( .A(n35871), .Z(n35869) );
  HS65_LH_BFX2 U20130 ( .A(n35872), .Z(n35870) );
  HS65_LH_BFX2 U20131 ( .A(n35873), .Z(n35871) );
  HS65_LH_BFX2 U20132 ( .A(n35874), .Z(n35872) );
  HS65_LH_BFX2 U20133 ( .A(n35875), .Z(n35873) );
  HS65_LH_BFX2 U20134 ( .A(n2237), .Z(n35874) );
  HS65_LH_BFX2 U20135 ( .A(n2238), .Z(n35875) );
  HS65_LH_BFX2 U20136 ( .A(n35878), .Z(n35876) );
  HS65_LH_BFX2 U20137 ( .A(n35879), .Z(n35877) );
  HS65_LH_BFX2 U20138 ( .A(n35880), .Z(n35878) );
  HS65_LH_BFX2 U20139 ( .A(n35881), .Z(n35879) );
  HS65_LH_BFX2 U20140 ( .A(n35882), .Z(n35880) );
  HS65_LH_BFX2 U20141 ( .A(n35883), .Z(n35881) );
  HS65_LH_BFX2 U20142 ( .A(n35884), .Z(n35882) );
  HS65_LH_BFX2 U20143 ( .A(n35885), .Z(n35883) );
  HS65_LH_BFX2 U20144 ( .A(n35886), .Z(n35884) );
  HS65_LH_BFX2 U20145 ( .A(n35887), .Z(n35885) );
  HS65_LH_BFX2 U20146 ( .A(n35888), .Z(n35886) );
  HS65_LH_BFX2 U20147 ( .A(n35889), .Z(n35887) );
  HS65_LH_BFX2 U20148 ( .A(n35890), .Z(n35888) );
  HS65_LH_BFX2 U20149 ( .A(n35891), .Z(n35889) );
  HS65_LH_BFX2 U20150 ( .A(n35892), .Z(n35890) );
  HS65_LH_BFX2 U20151 ( .A(n35893), .Z(n35891) );
  HS65_LH_BFX2 U20152 ( .A(n35894), .Z(n35892) );
  HS65_LH_BFX2 U20153 ( .A(n35895), .Z(n35893) );
  HS65_LH_BFX2 U20154 ( .A(n35896), .Z(n35894) );
  HS65_LH_BFX2 U20155 ( .A(n35897), .Z(n35895) );
  HS65_LH_BFX2 U20156 ( .A(n35898), .Z(n35896) );
  HS65_LH_BFX2 U20157 ( .A(n35899), .Z(n35897) );
  HS65_LH_BFX2 U20158 ( .A(n35900), .Z(n35898) );
  HS65_LH_BFX2 U20159 ( .A(n35901), .Z(n35899) );
  HS65_LH_BFX2 U20160 ( .A(n35902), .Z(n35900) );
  HS65_LH_BFX2 U20161 ( .A(n35903), .Z(n35901) );
  HS65_LH_BFX2 U20162 ( .A(n35904), .Z(n35902) );
  HS65_LH_BFX2 U20163 ( .A(n35905), .Z(n35903) );
  HS65_LH_BFX2 U20164 ( .A(n1997), .Z(n35904) );
  HS65_LH_BFX2 U20165 ( .A(n1998), .Z(n35905) );
  HS65_LH_BFX2 U20166 ( .A(n35909), .Z(n35906) );
  HS65_LH_BFX2 U20167 ( .A(n37717), .Z(n35907) );
  HS65_LH_BFX2 U20168 ( .A(n35940), .Z(n35908) );
  HS65_LH_BFX2 U20169 ( .A(n35911), .Z(n35909) );
  HS65_LH_BFX2 U20170 ( .A(n2117), .Z(n35910) );
  HS65_LH_BFX2 U20171 ( .A(n35913), .Z(n35911) );
  HS65_LH_BFX2 U20172 ( .A(n35910), .Z(n35912) );
  HS65_LH_BFX2 U20173 ( .A(n35915), .Z(n35913) );
  HS65_LH_BFX2 U20174 ( .A(n35912), .Z(n35914) );
  HS65_LH_BFX2 U20175 ( .A(n35917), .Z(n35915) );
  HS65_LH_BFX2 U20176 ( .A(n35914), .Z(n35916) );
  HS65_LH_BFX2 U20177 ( .A(n35919), .Z(n35917) );
  HS65_LH_BFX2 U20178 ( .A(n35916), .Z(n35918) );
  HS65_LH_BFX2 U20179 ( .A(n35921), .Z(n35919) );
  HS65_LH_BFX2 U20180 ( .A(n35918), .Z(n35920) );
  HS65_LH_BFX2 U20181 ( .A(n35923), .Z(n35921) );
  HS65_LH_BFX2 U20182 ( .A(n35920), .Z(n35922) );
  HS65_LH_BFX2 U20183 ( .A(n35925), .Z(n35923) );
  HS65_LH_BFX2 U20184 ( .A(n35922), .Z(n35924) );
  HS65_LH_BFX2 U20185 ( .A(n35927), .Z(n35925) );
  HS65_LH_BFX2 U20186 ( .A(n35924), .Z(n35926) );
  HS65_LH_BFX2 U20187 ( .A(n35929), .Z(n35927) );
  HS65_LH_BFX2 U20188 ( .A(n35926), .Z(n35928) );
  HS65_LH_BFX2 U20189 ( .A(n35931), .Z(n35929) );
  HS65_LH_BFX2 U20190 ( .A(n35928), .Z(n35930) );
  HS65_LH_BFX2 U20191 ( .A(n35934), .Z(n35931) );
  HS65_LH_BFX2 U20192 ( .A(n35930), .Z(n35932) );
  HS65_LH_IVX2 U20193 ( .A(n35938), .Z(n35933) );
  HS65_LH_IVX2 U20194 ( .A(n35933), .Z(n35934) );
  HS65_LH_IVX2 U20195 ( .A(n16262), .Z(n35935) );
  HS65_LH_IVX2 U20196 ( .A(n35935), .Z(n35936) );
  HS65_LH_IVX2 U20197 ( .A(n2118), .Z(n35937) );
  HS65_LH_IVX2 U20198 ( .A(n35937), .Z(n35938) );
  HS65_LH_IVX2 U20199 ( .A(n35932), .Z(n35939) );
  HS65_LH_IVX2 U20200 ( .A(n35939), .Z(n35940) );
  HS65_LH_BFX2 U20201 ( .A(n35946), .Z(n35941) );
  HS65_LH_BFX2 U20202 ( .A(n37666), .Z(n35942) );
  HS65_LH_BFX2 U20203 ( .A(n2190), .Z(n35943) );
  HS65_LH_IVX2 U20204 ( .A(n35948), .Z(n35944) );
  HS65_LH_IVX2 U20205 ( .A(n35944), .Z(n35945) );
  HS65_LH_BFX2 U20206 ( .A(n35947), .Z(n35946) );
  HS65_LH_BFX2 U20207 ( .A(n35949), .Z(n35947) );
  HS65_LH_BFX2 U20208 ( .A(n35950), .Z(n35948) );
  HS65_LH_BFX2 U20209 ( .A(n35951), .Z(n35949) );
  HS65_LH_BFX2 U20210 ( .A(n35952), .Z(n35950) );
  HS65_LH_BFX2 U20211 ( .A(n35953), .Z(n35951) );
  HS65_LH_BFX2 U20212 ( .A(n35954), .Z(n35952) );
  HS65_LH_BFX2 U20213 ( .A(n35955), .Z(n35953) );
  HS65_LH_BFX2 U20214 ( .A(n35956), .Z(n35954) );
  HS65_LH_BFX2 U20215 ( .A(n35957), .Z(n35955) );
  HS65_LH_BFX2 U20216 ( .A(n35958), .Z(n35956) );
  HS65_LH_BFX2 U20217 ( .A(n35959), .Z(n35957) );
  HS65_LH_BFX2 U20218 ( .A(n35960), .Z(n35958) );
  HS65_LH_BFX2 U20219 ( .A(n35961), .Z(n35959) );
  HS65_LH_BFX2 U20220 ( .A(n35962), .Z(n35960) );
  HS65_LH_BFX2 U20221 ( .A(n35963), .Z(n35961) );
  HS65_LH_BFX2 U20222 ( .A(n35964), .Z(n35962) );
  HS65_LH_BFX2 U20223 ( .A(n35965), .Z(n35963) );
  HS65_LH_BFX2 U20224 ( .A(n35966), .Z(n35964) );
  HS65_LH_BFX2 U20225 ( .A(n35967), .Z(n35965) );
  HS65_LH_BFX2 U20226 ( .A(n35968), .Z(n35966) );
  HS65_LH_BFX2 U20227 ( .A(n35969), .Z(n35967) );
  HS65_LH_BFX2 U20228 ( .A(n35970), .Z(n35968) );
  HS65_LH_BFX2 U20229 ( .A(n35971), .Z(n35969) );
  HS65_LH_BFX2 U20230 ( .A(n35972), .Z(n35970) );
  HS65_LH_BFX2 U20231 ( .A(n35973), .Z(n35971) );
  HS65_LH_BFX2 U20232 ( .A(n35943), .Z(n35972) );
  HS65_LH_BFX2 U20233 ( .A(n2189), .Z(n35973) );
  HS65_LH_BFX2 U20234 ( .A(n35976), .Z(n35974) );
  HS65_LH_BFX2 U20235 ( .A(n2021), .Z(n35975) );
  HS65_LH_BFX2 U20236 ( .A(n35978), .Z(n35976) );
  HS65_LH_BFX2 U20237 ( .A(n35975), .Z(n35977) );
  HS65_LH_BFX2 U20238 ( .A(n35980), .Z(n35978) );
  HS65_LH_BFX2 U20239 ( .A(n35977), .Z(n35979) );
  HS65_LH_BFX2 U20240 ( .A(n35982), .Z(n35980) );
  HS65_LH_BFX2 U20241 ( .A(n35979), .Z(n35981) );
  HS65_LH_BFX2 U20242 ( .A(n35984), .Z(n35982) );
  HS65_LH_BFX2 U20243 ( .A(n35981), .Z(n35983) );
  HS65_LH_BFX2 U20244 ( .A(n35986), .Z(n35984) );
  HS65_LH_BFX2 U20245 ( .A(n35983), .Z(n35985) );
  HS65_LH_BFX2 U20246 ( .A(n35988), .Z(n35986) );
  HS65_LH_BFX2 U20247 ( .A(n35985), .Z(n35987) );
  HS65_LH_BFX2 U20248 ( .A(n35990), .Z(n35988) );
  HS65_LH_BFX2 U20249 ( .A(n35987), .Z(n35989) );
  HS65_LH_BFX2 U20250 ( .A(n35992), .Z(n35990) );
  HS65_LH_BFX2 U20251 ( .A(n35989), .Z(n35991) );
  HS65_LH_BFX2 U20252 ( .A(n35994), .Z(n35992) );
  HS65_LH_BFX2 U20253 ( .A(n35991), .Z(n35993) );
  HS65_LH_BFX2 U20254 ( .A(n35996), .Z(n35994) );
  HS65_LH_BFX2 U20255 ( .A(n35993), .Z(n35995) );
  HS65_LH_BFX2 U20256 ( .A(n35998), .Z(n35996) );
  HS65_LH_BFX2 U20257 ( .A(n35995), .Z(n35997) );
  HS65_LH_BFX2 U20258 ( .A(n36001), .Z(n35998) );
  HS65_LH_BFX2 U20259 ( .A(n35997), .Z(n35999) );
  HS65_LH_IVX2 U20260 ( .A(n36006), .Z(n36000) );
  HS65_LH_IVX2 U20261 ( .A(n36000), .Z(n36001) );
  HS65_LH_BFX2 U20262 ( .A(n35999), .Z(n36002) );
  HS65_LH_IVX2 U20263 ( .A(n36002), .Z(n36003) );
  HS65_LH_IVX2 U20264 ( .A(n36003), .Z(n36004) );
  HS65_LH_IVX2 U20265 ( .A(n2022), .Z(n36005) );
  HS65_LH_IVX2 U20266 ( .A(n36005), .Z(n36006) );
  HS65_LH_BFX2 U20267 ( .A(n36010), .Z(n36007) );
  HS65_LH_BFX2 U20268 ( .A(n36013), .Z(n36008) );
  HS65_LH_IVX2 U20269 ( .A(n36015), .Z(n36009) );
  HS65_LH_IVX2 U20270 ( .A(n36009), .Z(n36010) );
  HS65_LH_BFX2 U20271 ( .A(n2141), .Z(n36011) );
  HS65_LH_IVX2 U20272 ( .A(n37424), .Z(n36012) );
  HS65_LH_IVX2 U20273 ( .A(n36012), .Z(n36013) );
  HS65_LH_BFX2 U20274 ( .A(n36011), .Z(n36014) );
  HS65_LH_BFX2 U20275 ( .A(n36017), .Z(n36015) );
  HS65_LH_BFX2 U20276 ( .A(n36014), .Z(n36016) );
  HS65_LH_BFX2 U20277 ( .A(n36019), .Z(n36017) );
  HS65_LH_BFX2 U20278 ( .A(n36016), .Z(n36018) );
  HS65_LH_BFX2 U20279 ( .A(n36021), .Z(n36019) );
  HS65_LH_BFX2 U20280 ( .A(n36018), .Z(n36020) );
  HS65_LH_BFX2 U20281 ( .A(n36023), .Z(n36021) );
  HS65_LH_BFX2 U20282 ( .A(n36020), .Z(n36022) );
  HS65_LH_BFX2 U20283 ( .A(n36025), .Z(n36023) );
  HS65_LH_BFX2 U20284 ( .A(n36022), .Z(n36024) );
  HS65_LH_BFX2 U20285 ( .A(n36027), .Z(n36025) );
  HS65_LH_BFX2 U20286 ( .A(n36024), .Z(n36026) );
  HS65_LH_BFX2 U20287 ( .A(n36029), .Z(n36027) );
  HS65_LH_BFX2 U20288 ( .A(n36026), .Z(n36028) );
  HS65_LH_BFX2 U20289 ( .A(n36031), .Z(n36029) );
  HS65_LH_BFX2 U20290 ( .A(n36028), .Z(n36030) );
  HS65_LH_BFX2 U20291 ( .A(n36033), .Z(n36031) );
  HS65_LH_BFX2 U20292 ( .A(n36030), .Z(n36032) );
  HS65_LH_BFX2 U20293 ( .A(n36036), .Z(n36033) );
  HS65_LH_BFX2 U20294 ( .A(n36032), .Z(n36034) );
  HS65_LH_IVX2 U20295 ( .A(n36041), .Z(n36035) );
  HS65_LH_IVX2 U20296 ( .A(n36035), .Z(n36036) );
  HS65_LH_BFX2 U20297 ( .A(n36034), .Z(n36037) );
  HS65_LH_IVX2 U20298 ( .A(n36044), .Z(n36038) );
  HS65_LH_IVX2 U20299 ( .A(n36038), .Z(n36039) );
  HS65_LH_IVX2 U20300 ( .A(n36043), .Z(n36040) );
  HS65_LH_IVX2 U20301 ( .A(n36040), .Z(n36041) );
  HS65_LH_IVX2 U20302 ( .A(n2142), .Z(n36042) );
  HS65_LH_IVX2 U20303 ( .A(n36042), .Z(n36043) );
  HS65_LH_BFX2 U20304 ( .A(n36037), .Z(n36044) );
  HS65_LH_BFX2 U20305 ( .A(n36049), .Z(n36046) );
  HS65_LH_BFX2 U20306 ( .A(n36052), .Z(n36047) );
  HS65_LH_IVX2 U20307 ( .A(n36057), .Z(n36048) );
  HS65_LH_IVX2 U20308 ( .A(n36048), .Z(n36049) );
  HS65_LH_BFX2 U20309 ( .A(n2477), .Z(n36050) );
  HS65_LH_IVX2 U20310 ( .A(n36058), .Z(n36051) );
  HS65_LH_IVX2 U20311 ( .A(n36051), .Z(n36052) );
  HS65_LH_IVX2 U20312 ( .A(n36056), .Z(n36053) );
  HS65_LH_IVX2 U20313 ( .A(n36053), .Z(n36054) );
  HS65_LH_IVX2 U20314 ( .A(n36064), .Z(n36055) );
  HS65_LH_IVX2 U20315 ( .A(n36055), .Z(n36056) );
  HS65_LH_BFX2 U20316 ( .A(n36060), .Z(n36057) );
  HS65_LH_BFX2 U20317 ( .A(n36062), .Z(n36058) );
  HS65_LH_IVX2 U20318 ( .A(n36066), .Z(n36059) );
  HS65_LH_IVX2 U20319 ( .A(n36059), .Z(n36060) );
  HS65_LH_IVX2 U20320 ( .A(n36068), .Z(n36061) );
  HS65_LH_IVX2 U20321 ( .A(n36061), .Z(n36062) );
  HS65_LH_IVX2 U20322 ( .A(n36070), .Z(n36063) );
  HS65_LH_IVX2 U20323 ( .A(n36063), .Z(n36064) );
  HS65_LH_IVX2 U20324 ( .A(n36072), .Z(n36065) );
  HS65_LH_IVX2 U20325 ( .A(n36065), .Z(n36066) );
  HS65_LH_IVX2 U20326 ( .A(n36074), .Z(n36067) );
  HS65_LH_IVX2 U20327 ( .A(n36067), .Z(n36068) );
  HS65_LH_IVX2 U20328 ( .A(n36076), .Z(n36069) );
  HS65_LH_IVX2 U20329 ( .A(n36069), .Z(n36070) );
  HS65_LH_IVX2 U20330 ( .A(n36078), .Z(n36071) );
  HS65_LH_IVX2 U20331 ( .A(n36071), .Z(n36072) );
  HS65_LH_IVX2 U20332 ( .A(n36080), .Z(n36073) );
  HS65_LH_IVX2 U20333 ( .A(n36073), .Z(n36074) );
  HS65_LH_IVX2 U20334 ( .A(n36082), .Z(n36075) );
  HS65_LH_IVX2 U20335 ( .A(n36075), .Z(n36076) );
  HS65_LH_IVX2 U20336 ( .A(n36084), .Z(n36077) );
  HS65_LH_IVX2 U20337 ( .A(n36077), .Z(n36078) );
  HS65_LH_IVX2 U20338 ( .A(n36086), .Z(n36079) );
  HS65_LH_IVX2 U20339 ( .A(n36079), .Z(n36080) );
  HS65_LH_IVX2 U20340 ( .A(n36093), .Z(n36081) );
  HS65_LH_IVX2 U20341 ( .A(n36081), .Z(n36082) );
  HS65_LH_IVX2 U20342 ( .A(n36088), .Z(n36083) );
  HS65_LH_IVX2 U20343 ( .A(n36083), .Z(n36084) );
  HS65_LH_IVX2 U20344 ( .A(n36091), .Z(n36085) );
  HS65_LH_IVX2 U20345 ( .A(n36085), .Z(n36086) );
  HS65_LH_IVX2 U20346 ( .A(n36098), .Z(n36087) );
  HS65_LH_IVX2 U20347 ( .A(n36087), .Z(n36088) );
  HS65_LH_BFX2 U20348 ( .A(n36050), .Z(n36089) );
  HS65_LH_IVX2 U20349 ( .A(n36095), .Z(n36090) );
  HS65_LH_IVX2 U20350 ( .A(n36090), .Z(n36091) );
  HS65_LH_IVX2 U20351 ( .A(n36097), .Z(n36092) );
  HS65_LH_IVX2 U20352 ( .A(n36092), .Z(n36093) );
  HS65_LH_IVX2 U20353 ( .A(n36100), .Z(n36094) );
  HS65_LH_IVX2 U20354 ( .A(n36094), .Z(n36095) );
  HS65_LH_IVX2 U20355 ( .A(n36102), .Z(n36096) );
  HS65_LH_IVX2 U20356 ( .A(n36096), .Z(n36097) );
  HS65_LH_BFX2 U20357 ( .A(n36103), .Z(n36098) );
  HS65_LH_IVX2 U20358 ( .A(n36105), .Z(n36099) );
  HS65_LH_IVX2 U20359 ( .A(n36099), .Z(n36100) );
  HS65_LH_IVX2 U20360 ( .A(n36107), .Z(n36101) );
  HS65_LH_IVX2 U20361 ( .A(n36101), .Z(n36102) );
  HS65_LH_BFX2 U20362 ( .A(n36108), .Z(n36103) );
  HS65_LH_IVX2 U20363 ( .A(n36110), .Z(n36104) );
  HS65_LH_IVX2 U20364 ( .A(n36104), .Z(n36105) );
  HS65_LH_IVX2 U20365 ( .A(n36114), .Z(n36106) );
  HS65_LH_IVX2 U20366 ( .A(n36106), .Z(n36107) );
  HS65_LH_BFX2 U20367 ( .A(n36111), .Z(n36108) );
  HS65_LH_IVX2 U20368 ( .A(n36116), .Z(n36109) );
  HS65_LH_IVX2 U20369 ( .A(n36109), .Z(n36110) );
  HS65_LH_BFX2 U20370 ( .A(n36117), .Z(n36111) );
  HS65_LH_BFX2 U20371 ( .A(n36089), .Z(n36112) );
  HS65_LH_IVX2 U20372 ( .A(n36121), .Z(n36113) );
  HS65_LH_IVX2 U20373 ( .A(n36113), .Z(n36114) );
  HS65_LH_IVX2 U20374 ( .A(n36119), .Z(n36115) );
  HS65_LH_IVX2 U20375 ( .A(n36115), .Z(n36116) );
  HS65_LH_BFX2 U20376 ( .A(n36120), .Z(n36117) );
  HS65_LH_IVX2 U20377 ( .A(n36123), .Z(n36118) );
  HS65_LH_IVX2 U20378 ( .A(n36118), .Z(n36119) );
  HS65_LH_BFX2 U20379 ( .A(n2478), .Z(n36120) );
  HS65_LH_BFX2 U20380 ( .A(n36112), .Z(n36121) );
  HS65_LH_IVX2 U20381 ( .A(n36124), .Z(n36122) );
  HS65_LH_IVX2 U20382 ( .A(n36122), .Z(n36123) );
  HS65_LH_BFX2 U20383 ( .A(n36125), .Z(n36124) );
  HS65_LH_BFX2 U20384 ( .A(n36126), .Z(n36125) );
  HS65_LH_BFX2 U20385 ( .A(n17923), .Z(n36126) );
  HS65_LH_BFX2 U20386 ( .A(n36129), .Z(n36127) );
  HS65_LH_IVX2 U20387 ( .A(n36136), .Z(n36128) );
  HS65_LH_IVX2 U20388 ( .A(n36128), .Z(n36129) );
  HS65_LH_BFX2 U20389 ( .A(n36133), .Z(n36130) );
  HS65_LH_BFX2 U20390 ( .A(n2574), .Z(n36131) );
  HS65_LH_IVX2 U20391 ( .A(n37211), .Z(n36132) );
  HS65_LH_IVX2 U20392 ( .A(n36132), .Z(n36133) );
  HS65_LH_IVX2 U20393 ( .A(n36137), .Z(n36134) );
  HS65_LH_IVX2 U20394 ( .A(n36134), .Z(n36135) );
  HS65_LH_BFX2 U20395 ( .A(n36138), .Z(n36136) );
  HS65_LH_BFX2 U20396 ( .A(n36139), .Z(n36137) );
  HS65_LH_BFX2 U20397 ( .A(n36140), .Z(n36138) );
  HS65_LH_BFX2 U20398 ( .A(n36141), .Z(n36139) );
  HS65_LH_BFX2 U20399 ( .A(n36142), .Z(n36140) );
  HS65_LH_BFX2 U20400 ( .A(n36143), .Z(n36141) );
  HS65_LH_BFX2 U20401 ( .A(n36144), .Z(n36142) );
  HS65_LH_BFX2 U20402 ( .A(n36145), .Z(n36143) );
  HS65_LH_BFX2 U20403 ( .A(n36146), .Z(n36144) );
  HS65_LH_BFX2 U20404 ( .A(n36147), .Z(n36145) );
  HS65_LH_BFX2 U20405 ( .A(n36148), .Z(n36146) );
  HS65_LH_BFX2 U20406 ( .A(n36149), .Z(n36147) );
  HS65_LH_BFX2 U20407 ( .A(n36150), .Z(n36148) );
  HS65_LH_BFX2 U20408 ( .A(n36151), .Z(n36149) );
  HS65_LH_BFX2 U20409 ( .A(n36152), .Z(n36150) );
  HS65_LH_BFX2 U20410 ( .A(n36153), .Z(n36151) );
  HS65_LH_BFX2 U20411 ( .A(n36154), .Z(n36152) );
  HS65_LH_BFX2 U20412 ( .A(n36155), .Z(n36153) );
  HS65_LH_BFX2 U20413 ( .A(n36156), .Z(n36154) );
  HS65_LH_BFX2 U20414 ( .A(n36157), .Z(n36155) );
  HS65_LH_BFX2 U20415 ( .A(n36160), .Z(n36156) );
  HS65_LH_BFX2 U20416 ( .A(n36159), .Z(n36157) );
  HS65_LH_BFX2 U20417 ( .A(n15885), .Z(n36158) );
  HS65_LH_BFX2 U20418 ( .A(n36161), .Z(n36159) );
  HS65_LH_BFX2 U20419 ( .A(n2573), .Z(n36160) );
  HS65_LH_BFX2 U20420 ( .A(n36131), .Z(n36161) );
  HS65_LH_BFX2 U20421 ( .A(n36168), .Z(n36162) );
  HS65_LH_IVX2 U20422 ( .A(n36170), .Z(n36163) );
  HS65_LH_IVX2 U20423 ( .A(n36163), .Z(n36164) );
  HS65_LH_BFX2 U20424 ( .A(n36169), .Z(n36165) );
  HS65_LH_BFX2 U20425 ( .A(n1973), .Z(n36166) );
  HS65_LH_IVX2 U20426 ( .A(n36180), .Z(n36167) );
  HS65_LH_IVX2 U20427 ( .A(n36167), .Z(n36168) );
  HS65_LH_BFX2 U20428 ( .A(n36173), .Z(n36169) );
  HS65_LH_BFX2 U20429 ( .A(n36172), .Z(n36170) );
  HS65_LH_IVX2 U20430 ( .A(n36176), .Z(n36171) );
  HS65_LH_IVX2 U20431 ( .A(n36171), .Z(n36172) );
  HS65_LH_BFX2 U20432 ( .A(n36177), .Z(n36173) );
  HS65_LH_BFX2 U20433 ( .A(n36166), .Z(n36174) );
  HS65_LH_IVX2 U20434 ( .A(n36182), .Z(n36175) );
  HS65_LH_IVX2 U20435 ( .A(n36175), .Z(n36176) );
  HS65_LH_BFX2 U20436 ( .A(n36183), .Z(n36177) );
  HS65_LH_BFX2 U20437 ( .A(n36174), .Z(n36178) );
  HS65_LH_IVX2 U20438 ( .A(n36185), .Z(n36179) );
  HS65_LH_IVX2 U20439 ( .A(n36179), .Z(n36180) );
  HS65_LH_IVX2 U20440 ( .A(n36895), .Z(n36181) );
  HS65_LH_IVX2 U20441 ( .A(n36181), .Z(n36182) );
  HS65_LH_BFX2 U20442 ( .A(n36184), .Z(n36183) );
  HS65_LH_BFX2 U20443 ( .A(n36187), .Z(n36184) );
  HS65_LH_BFX2 U20444 ( .A(n36188), .Z(n36185) );
  HS65_LH_BFX2 U20445 ( .A(n32445), .Z(n36186) );
  HS65_LH_BFX2 U20446 ( .A(n36190), .Z(n36187) );
  HS65_LH_BFX2 U20447 ( .A(n36191), .Z(n36188) );
  HS65_LH_BFX2 U20448 ( .A(n36186), .Z(n36189) );
  HS65_LH_BFX2 U20449 ( .A(n36192), .Z(n36190) );
  HS65_LH_BFX2 U20450 ( .A(n36193), .Z(n36191) );
  HS65_LH_BFX2 U20451 ( .A(n36194), .Z(n36192) );
  HS65_LH_BFX2 U20452 ( .A(n36195), .Z(n36193) );
  HS65_LH_BFX2 U20453 ( .A(n36196), .Z(n36194) );
  HS65_LH_BFX2 U20454 ( .A(n36197), .Z(n36195) );
  HS65_LH_BFX2 U20455 ( .A(n36198), .Z(n36196) );
  HS65_LH_BFX2 U20456 ( .A(n36199), .Z(n36197) );
  HS65_LH_BFX2 U20457 ( .A(n36200), .Z(n36198) );
  HS65_LH_BFX2 U20458 ( .A(n36201), .Z(n36199) );
  HS65_LH_BFX2 U20460 ( .A(n36202), .Z(n36200) );
  HS65_LH_BFX2 U20461 ( .A(n36203), .Z(n36201) );
  HS65_LH_BFX2 U20462 ( .A(n36204), .Z(n36202) );
  HS65_LH_BFX2 U20463 ( .A(n36205), .Z(n36203) );
  HS65_LH_BFX2 U20464 ( .A(n1974), .Z(n36204) );
  HS65_LH_BFX2 U20465 ( .A(n36178), .Z(n36205) );
  HS65_LH_BFX2 U20466 ( .A(n36208), .Z(n36206) );
  HS65_LH_BFX2 U20467 ( .A(n36209), .Z(n36207) );
  HS65_LH_BFX2 U20468 ( .A(n36210), .Z(n36208) );
  HS65_LH_BFX2 U20469 ( .A(n36211), .Z(n36209) );
  HS65_LH_BFX2 U20470 ( .A(n36212), .Z(n36210) );
  HS65_LH_BFX2 U20471 ( .A(n36213), .Z(n36211) );
  HS65_LH_BFX2 U20472 ( .A(n36214), .Z(n36212) );
  HS65_LH_BFX2 U20473 ( .A(n36215), .Z(n36213) );
  HS65_LH_BFX2 U20474 ( .A(n36216), .Z(n36214) );
  HS65_LH_BFX2 U20475 ( .A(n36217), .Z(n36215) );
  HS65_LH_BFX2 U20476 ( .A(n36218), .Z(n36216) );
  HS65_LH_BFX2 U20477 ( .A(n36219), .Z(n36217) );
  HS65_LH_BFX2 U20478 ( .A(n36220), .Z(n36218) );
  HS65_LH_BFX2 U20479 ( .A(n36221), .Z(n36219) );
  HS65_LH_BFX2 U20480 ( .A(n36222), .Z(n36220) );
  HS65_LH_BFX2 U20481 ( .A(n36223), .Z(n36221) );
  HS65_LH_BFX2 U20482 ( .A(n36224), .Z(n36222) );
  HS65_LH_BFX2 U20483 ( .A(n36225), .Z(n36223) );
  HS65_LH_BFX2 U20484 ( .A(n36226), .Z(n36224) );
  HS65_LH_BFX2 U20485 ( .A(n36227), .Z(n36225) );
  HS65_LH_BFX2 U20486 ( .A(n36228), .Z(n36226) );
  HS65_LH_BFX2 U20487 ( .A(n36229), .Z(n36227) );
  HS65_LH_BFX2 U20488 ( .A(n36230), .Z(n36228) );
  HS65_LH_BFX2 U20489 ( .A(n36231), .Z(n36229) );
  HS65_LH_BFX2 U20490 ( .A(n36232), .Z(n36230) );
  HS65_LH_BFX2 U20491 ( .A(n36233), .Z(n36231) );
  HS65_LH_BFX2 U20492 ( .A(n36234), .Z(n36232) );
  HS65_LH_BFX2 U20493 ( .A(n36235), .Z(n36233) );
  HS65_LH_BFX2 U20494 ( .A(n2069), .Z(n36234) );
  HS65_LH_BFX2 U20495 ( .A(n2070), .Z(n36235) );
  HS65_LH_IVX2 U20496 ( .A(n36241), .Z(n36236) );
  HS65_LH_IVX2 U20497 ( .A(n36236), .Z(n36237) );
  HS65_LH_BFX2 U20498 ( .A(n2285), .Z(n36238) );
  HS65_LH_BFX2 U20499 ( .A(n37075), .Z(n36239) );
  HS65_LH_BFX2 U20500 ( .A(n36238), .Z(n36240) );
  HS65_LH_BFX2 U20501 ( .A(n36243), .Z(n36241) );
  HS65_LH_BFX2 U20502 ( .A(n36240), .Z(n36242) );
  HS65_LH_BFX2 U20503 ( .A(n36245), .Z(n36243) );
  HS65_LH_BFX2 U20504 ( .A(n36242), .Z(n36244) );
  HS65_LH_BFX2 U20505 ( .A(n36247), .Z(n36245) );
  HS65_LH_BFX2 U20506 ( .A(n36244), .Z(n36246) );
  HS65_LH_BFX2 U20507 ( .A(n36249), .Z(n36247) );
  HS65_LH_BFX2 U20508 ( .A(n36246), .Z(n36248) );
  HS65_LH_BFX2 U20509 ( .A(n36251), .Z(n36249) );
  HS65_LH_BFX2 U20510 ( .A(n36248), .Z(n36250) );
  HS65_LH_BFX2 U20511 ( .A(n36253), .Z(n36251) );
  HS65_LH_BFX2 U20512 ( .A(n36250), .Z(n36252) );
  HS65_LH_BFX2 U20513 ( .A(n36255), .Z(n36253) );
  HS65_LH_BFX2 U20514 ( .A(n36252), .Z(n36254) );
  HS65_LH_BFX2 U20515 ( .A(n36257), .Z(n36255) );
  HS65_LH_BFX2 U20516 ( .A(n36254), .Z(n36256) );
  HS65_LH_BFX2 U20517 ( .A(n36259), .Z(n36257) );
  HS65_LH_BFX2 U20518 ( .A(n36256), .Z(n36258) );
  HS65_LH_BFX2 U20519 ( .A(n36261), .Z(n36259) );
  HS65_LH_BFX2 U20520 ( .A(n36258), .Z(n36260) );
  HS65_LH_BFX2 U20521 ( .A(n36263), .Z(n36261) );
  HS65_LH_BFX2 U20522 ( .A(n36260), .Z(n36262) );
  HS65_LH_BFX2 U20523 ( .A(n36267), .Z(n36263) );
  HS65_LH_IVX2 U20524 ( .A(n16123), .Z(n36265) );
  HS65_LH_IVX2 U20525 ( .A(n36265), .Z(n36266) );
  HS65_LH_BFX2 U20526 ( .A(n36269), .Z(n36267) );
  HS65_LH_IVX2 U20527 ( .A(n2286), .Z(n36268) );
  HS65_LH_IVX2 U20528 ( .A(n36268), .Z(n36269) );
  HS65_LH_IVX2 U20529 ( .A(n36262), .Z(n36270) );
  HS65_LH_IVX2 U20530 ( .A(n36270), .Z(n36271) );
  HS65_LH_BFX2 U20531 ( .A(n36274), .Z(n36272) );
  HS65_LH_NAND4ABX3 U20532 ( .A(n16185), .B(n16184), .C(n16183), .D(n16182), 
        .Z(n2213) );
  HS65_LH_IVX2 U20533 ( .A(n36277), .Z(n36273) );
  HS65_LH_IVX2 U20534 ( .A(n36273), .Z(n36274) );
  HS65_LH_NAND2X2 U20535 ( .A(n16187), .B(n16186), .Z(n16195) );
  HS65_LH_BFX2 U20536 ( .A(n16195), .Z(n36275) );
  HS65_LH_BFX2 U20537 ( .A(n36278), .Z(n36276) );
  HS65_LH_BFX2 U20538 ( .A(n36279), .Z(n36277) );
  HS65_LH_BFX2 U20539 ( .A(n36280), .Z(n36278) );
  HS65_LH_BFX2 U20540 ( .A(n36281), .Z(n36279) );
  HS65_LH_BFX2 U20541 ( .A(n36282), .Z(n36280) );
  HS65_LH_BFX2 U20542 ( .A(n36283), .Z(n36281) );
  HS65_LH_BFX2 U20543 ( .A(n36284), .Z(n36282) );
  HS65_LH_BFX2 U20544 ( .A(n36285), .Z(n36283) );
  HS65_LH_BFX2 U20545 ( .A(n36286), .Z(n36284) );
  HS65_LH_BFX2 U20546 ( .A(n36287), .Z(n36285) );
  HS65_LH_BFX2 U20547 ( .A(n36288), .Z(n36286) );
  HS65_LH_BFX2 U20548 ( .A(n36289), .Z(n36287) );
  HS65_LH_BFX2 U20549 ( .A(n36290), .Z(n36288) );
  HS65_LH_BFX2 U20550 ( .A(n36291), .Z(n36289) );
  HS65_LH_BFX2 U20551 ( .A(n36292), .Z(n36290) );
  HS65_LH_BFX2 U20552 ( .A(n36293), .Z(n36291) );
  HS65_LH_BFX2 U20553 ( .A(n36294), .Z(n36292) );
  HS65_LH_BFX2 U20554 ( .A(n36295), .Z(n36293) );
  HS65_LH_BFX2 U20555 ( .A(n36296), .Z(n36294) );
  HS65_LH_BFX2 U20556 ( .A(n36297), .Z(n36295) );
  HS65_LH_BFX2 U20557 ( .A(n36298), .Z(n36296) );
  HS65_LH_BFX2 U20558 ( .A(n36299), .Z(n36297) );
  HS65_LH_BFX2 U20559 ( .A(n36300), .Z(n36298) );
  HS65_LH_BFX2 U20560 ( .A(n36301), .Z(n36299) );
  HS65_LH_BFX2 U20561 ( .A(n36302), .Z(n36300) );
  HS65_LH_BFX2 U20562 ( .A(n36303), .Z(n36301) );
  HS65_LH_BFX2 U20563 ( .A(n2214), .Z(n36302) );
  HS65_LH_BFX2 U20564 ( .A(n2213), .Z(n36303) );
  HS65_LH_BFX2 U20565 ( .A(n36308), .Z(n36304) );
  HS65_LH_BFX2 U20566 ( .A(n36310), .Z(n36305) );
  HS65_LH_BFX2 U20567 ( .A(n36312), .Z(n36306) );
  HS65_LH_IVX2 U20568 ( .A(n36314), .Z(n36307) );
  HS65_LH_IVX2 U20569 ( .A(n36307), .Z(n36308) );
  HS65_LH_IVX2 U20570 ( .A(n36316), .Z(n36309) );
  HS65_LH_IVX2 U20571 ( .A(n36309), .Z(n36310) );
  HS65_LH_IVX2 U20572 ( .A(n36318), .Z(n36311) );
  HS65_LH_IVX2 U20573 ( .A(n36311), .Z(n36312) );
  HS65_LH_IVX2 U20574 ( .A(n36320), .Z(n36313) );
  HS65_LH_IVX2 U20575 ( .A(n36313), .Z(n36314) );
  HS65_LH_IVX2 U20576 ( .A(n36322), .Z(n36315) );
  HS65_LH_IVX2 U20577 ( .A(n36315), .Z(n36316) );
  HS65_LH_IVX2 U20578 ( .A(n36324), .Z(n36317) );
  HS65_LH_IVX2 U20579 ( .A(n36317), .Z(n36318) );
  HS65_LH_IVX2 U20580 ( .A(n36326), .Z(n36319) );
  HS65_LH_IVX2 U20582 ( .A(n36319), .Z(n36320) );
  HS65_LH_IVX2 U20583 ( .A(n36328), .Z(n36321) );
  HS65_LH_IVX2 U20584 ( .A(n36321), .Z(n36322) );
  HS65_LH_IVX2 U20585 ( .A(n36330), .Z(n36323) );
  HS65_LH_IVX2 U20586 ( .A(n36323), .Z(n36324) );
  HS65_LH_IVX2 U20587 ( .A(n36332), .Z(n36325) );
  HS65_LH_IVX2 U20588 ( .A(n36325), .Z(n36326) );
  HS65_LH_IVX2 U20589 ( .A(n36334), .Z(n36327) );
  HS65_LH_IVX2 U20590 ( .A(n36327), .Z(n36328) );
  HS65_LH_IVX2 U20591 ( .A(n36336), .Z(n36329) );
  HS65_LH_IVX2 U20592 ( .A(n36329), .Z(n36330) );
  HS65_LH_IVX2 U20593 ( .A(n36338), .Z(n36331) );
  HS65_LH_IVX2 U20594 ( .A(n36331), .Z(n36332) );
  HS65_LH_IVX2 U20595 ( .A(n36340), .Z(n36333) );
  HS65_LH_IVX2 U20596 ( .A(n36333), .Z(n36334) );
  HS65_LH_IVX2 U20597 ( .A(n36342), .Z(n36335) );
  HS65_LH_IVX2 U20598 ( .A(n36335), .Z(n36336) );
  HS65_LH_IVX2 U20599 ( .A(n36344), .Z(n36337) );
  HS65_LH_IVX2 U20600 ( .A(n36337), .Z(n36338) );
  HS65_LH_IVX2 U20601 ( .A(n36346), .Z(n36339) );
  HS65_LH_IVX2 U20602 ( .A(n36339), .Z(n36340) );
  HS65_LH_IVX2 U20603 ( .A(n36348), .Z(n36341) );
  HS65_LH_IVX2 U20604 ( .A(n36341), .Z(n36342) );
  HS65_LH_IVX2 U20605 ( .A(n36350), .Z(n36343) );
  HS65_LH_IVX2 U20606 ( .A(n36343), .Z(n36344) );
  HS65_LH_IVX2 U20607 ( .A(n36352), .Z(n36345) );
  HS65_LH_IVX2 U20608 ( .A(n36345), .Z(n36346) );
  HS65_LH_IVX2 U20609 ( .A(n36354), .Z(n36347) );
  HS65_LH_IVX2 U20610 ( .A(n36347), .Z(n36348) );
  HS65_LH_IVX2 U20611 ( .A(n36356), .Z(n36349) );
  HS65_LH_IVX2 U20612 ( .A(n36349), .Z(n36350) );
  HS65_LH_IVX2 U20613 ( .A(n36358), .Z(n36351) );
  HS65_LH_IVX2 U20614 ( .A(n36351), .Z(n36352) );
  HS65_LH_IVX2 U20615 ( .A(n36360), .Z(n36353) );
  HS65_LH_IVX2 U20616 ( .A(n36353), .Z(n36354) );
  HS65_LH_IVX2 U20617 ( .A(n36362), .Z(n36355) );
  HS65_LH_IVX2 U20618 ( .A(n36355), .Z(n36356) );
  HS65_LH_IVX2 U20619 ( .A(n36364), .Z(n36357) );
  HS65_LH_IVX2 U20620 ( .A(n36357), .Z(n36358) );
  HS65_LH_IVX2 U20621 ( .A(n36366), .Z(n36359) );
  HS65_LH_IVX2 U20622 ( .A(n36359), .Z(n36360) );
  HS65_LH_IVX2 U20623 ( .A(n36368), .Z(n36361) );
  HS65_LH_IVX2 U20624 ( .A(n36361), .Z(n36362) );
  HS65_LH_IVX2 U20625 ( .A(n36370), .Z(n36363) );
  HS65_LH_IVX2 U20626 ( .A(n36363), .Z(n36364) );
  HS65_LH_IVX2 U20627 ( .A(n36372), .Z(n36365) );
  HS65_LH_IVX2 U20628 ( .A(n36365), .Z(n36366) );
  HS65_LH_IVX2 U20629 ( .A(n36374), .Z(n36367) );
  HS65_LH_IVX2 U20630 ( .A(n36367), .Z(n36368) );
  HS65_LH_IVX2 U20631 ( .A(n36376), .Z(n36369) );
  HS65_LH_IVX2 U20632 ( .A(n36369), .Z(n36370) );
  HS65_LH_IVX2 U20633 ( .A(n36378), .Z(n36371) );
  HS65_LH_IVX2 U20634 ( .A(n36371), .Z(n36372) );
  HS65_LH_IVX2 U20635 ( .A(n36383), .Z(n36373) );
  HS65_LH_IVX2 U20636 ( .A(n36373), .Z(n36374) );
  HS65_LH_IVX2 U20637 ( .A(n36380), .Z(n36375) );
  HS65_LH_IVX2 U20638 ( .A(n36375), .Z(n36376) );
  HS65_LH_IVX2 U20639 ( .A(n36382), .Z(n36377) );
  HS65_LH_IVX2 U20640 ( .A(n36377), .Z(n36378) );
  HS65_LH_IVX2 U20641 ( .A(n2333), .Z(n36379) );
  HS65_LH_IVX2 U20642 ( .A(n36379), .Z(n36380) );
  HS65_LH_IVX2 U20643 ( .A(n2334), .Z(n36381) );
  HS65_LH_IVX2 U20644 ( .A(n36381), .Z(n36382) );
  HS65_LH_BFX2 U20645 ( .A(n36388), .Z(n36383) );
  HS65_LH_IVX2 U20646 ( .A(n36384), .Z(n36385) );
  HS65_LH_IVX2 U20647 ( .A(n16083), .Z(n36386) );
  HS65_LH_IVX2 U20648 ( .A(n36386), .Z(n36387) );
  HS65_LH_BFX2 U20649 ( .A(n36389), .Z(n36388) );
  HS65_LH_BFX2 U20650 ( .A(n36390), .Z(n36389) );
  HS65_LH_BFX2 U20651 ( .A(n36391), .Z(n36390) );
  HS65_LH_BFX2 U20652 ( .A(n36392), .Z(n36391) );
  HS65_LH_BFX2 U20653 ( .A(n17984), .Z(n36392) );
  HS65_LH_IVX2 U20654 ( .A(n37585), .Z(n36393) );
  HS65_LH_IVX2 U20655 ( .A(n36393), .Z(n36394) );
  HS65_LH_BFX2 U20656 ( .A(n36397), .Z(n36395) );
  HS65_LH_BFX2 U20657 ( .A(n36398), .Z(n36396) );
  HS65_LH_BFX2 U20658 ( .A(n36399), .Z(n36397) );
  HS65_LH_BFX2 U20659 ( .A(n36400), .Z(n36398) );
  HS65_LH_BFX2 U20660 ( .A(n36401), .Z(n36399) );
  HS65_LH_BFX2 U20661 ( .A(n36402), .Z(n36400) );
  HS65_LH_BFX2 U20662 ( .A(n36403), .Z(n36401) );
  HS65_LH_BFX2 U20663 ( .A(n36404), .Z(n36402) );
  HS65_LH_BFX2 U20664 ( .A(n36405), .Z(n36403) );
  HS65_LH_BFX2 U20665 ( .A(n36406), .Z(n36404) );
  HS65_LH_BFX2 U20666 ( .A(n36407), .Z(n36405) );
  HS65_LH_BFX2 U20667 ( .A(n36408), .Z(n36406) );
  HS65_LH_BFX2 U20668 ( .A(n36409), .Z(n36407) );
  HS65_LH_BFX2 U20669 ( .A(n36410), .Z(n36408) );
  HS65_LH_BFX2 U20670 ( .A(n36411), .Z(n36409) );
  HS65_LH_BFX2 U20671 ( .A(n36412), .Z(n36410) );
  HS65_LH_BFX2 U20672 ( .A(n36413), .Z(n36411) );
  HS65_LH_BFX2 U20673 ( .A(n36414), .Z(n36412) );
  HS65_LH_BFX2 U20674 ( .A(n36415), .Z(n36413) );
  HS65_LH_BFX2 U20675 ( .A(n36416), .Z(n36414) );
  HS65_LH_BFX2 U20676 ( .A(n36417), .Z(n36415) );
  HS65_LH_BFX2 U20677 ( .A(n36418), .Z(n36416) );
  HS65_LH_BFX2 U20678 ( .A(n36419), .Z(n36417) );
  HS65_LH_BFX2 U20679 ( .A(n36420), .Z(n36418) );
  HS65_LH_BFX2 U20680 ( .A(n36421), .Z(n36419) );
  HS65_LH_BFX2 U20681 ( .A(n36422), .Z(n36420) );
  HS65_LH_BFX2 U20682 ( .A(n36426), .Z(n36421) );
  HS65_LH_BFX2 U20683 ( .A(n36424), .Z(n36422) );
  HS65_LH_BFX2 U20684 ( .A(n36425), .Z(n36423) );
  HS65_LH_BFX2 U20685 ( .A(n2166), .Z(n36424) );
  HS65_LH_BFX2 U20686 ( .A(n16223), .Z(n36425) );
  HS65_LH_BFX2 U20687 ( .A(n2165), .Z(n36426) );
  HS65_LH_BFX2 U20688 ( .A(n36429), .Z(n36427) );
  HS65_LH_IVX2 U20689 ( .A(n36434), .Z(n36428) );
  HS65_LH_IVX2 U20690 ( .A(n36428), .Z(n36429) );
  HS65_LH_BFX2 U20691 ( .A(n36432), .Z(n36430) );
  HS65_LH_BFX2 U20692 ( .A(n2406), .Z(n36431) );
  HS65_LH_BFX2 U20693 ( .A(n36435), .Z(n36432) );
  HS65_LH_BFX2 U20694 ( .A(n36431), .Z(n36433) );
  HS65_LH_BFX2 U20695 ( .A(n36437), .Z(n36434) );
  HS65_LH_BFX2 U20696 ( .A(n36438), .Z(n36435) );
  HS65_LH_BFX2 U20697 ( .A(n36433), .Z(n36436) );
  HS65_LH_BFX2 U20698 ( .A(n36440), .Z(n36437) );
  HS65_LH_BFX2 U20699 ( .A(n36441), .Z(n36438) );
  HS65_LH_BFX2 U20700 ( .A(n36436), .Z(n36439) );
  HS65_LH_BFX2 U20701 ( .A(n36443), .Z(n36440) );
  HS65_LH_BFX2 U20702 ( .A(n36444), .Z(n36441) );
  HS65_LH_BFX2 U20703 ( .A(n36439), .Z(n36442) );
  HS65_LH_BFX2 U20704 ( .A(n36446), .Z(n36443) );
  HS65_LH_BFX2 U20705 ( .A(n36447), .Z(n36444) );
  HS65_LH_BFX2 U20706 ( .A(n36442), .Z(n36445) );
  HS65_LH_BFX2 U20707 ( .A(n36449), .Z(n36446) );
  HS65_LH_BFX2 U20708 ( .A(n36450), .Z(n36447) );
  HS65_LH_BFX2 U20709 ( .A(n36445), .Z(n36448) );
  HS65_LH_BFX2 U20710 ( .A(n36452), .Z(n36449) );
  HS65_LH_BFX2 U20711 ( .A(n36453), .Z(n36450) );
  HS65_LH_BFX2 U20712 ( .A(n36448), .Z(n36451) );
  HS65_LH_BFX2 U20713 ( .A(n36455), .Z(n36452) );
  HS65_LH_BFX2 U20714 ( .A(n36456), .Z(n36453) );
  HS65_LH_BFX2 U20715 ( .A(n36451), .Z(n36454) );
  HS65_LH_BFX2 U20716 ( .A(n36458), .Z(n36455) );
  HS65_LH_BFX2 U20717 ( .A(n36459), .Z(n36456) );
  HS65_LH_BFX2 U20718 ( .A(n36454), .Z(n36457) );
  HS65_LH_BFX2 U20719 ( .A(n36461), .Z(n36458) );
  HS65_LH_BFX2 U20720 ( .A(n36462), .Z(n36459) );
  HS65_LH_BFX2 U20721 ( .A(n36457), .Z(n36460) );
  HS65_LH_BFX2 U20722 ( .A(n36464), .Z(n36461) );
  HS65_LH_BFX2 U20723 ( .A(n36465), .Z(n36462) );
  HS65_LH_BFX2 U20724 ( .A(n36460), .Z(n36463) );
  HS65_LH_BFX2 U20725 ( .A(n36467), .Z(n36464) );
  HS65_LH_BFX2 U20726 ( .A(n36468), .Z(n36465) );
  HS65_LH_BFX2 U20727 ( .A(n36463), .Z(n36466) );
  HS65_LH_BFX2 U20728 ( .A(n36475), .Z(n36467) );
  HS65_LH_BFX2 U20729 ( .A(n36471), .Z(n36468) );
  HS65_LH_BFX2 U20730 ( .A(n16033), .Z(n36469) );
  HS65_LH_IVX2 U20731 ( .A(n36477), .Z(n36470) );
  HS65_LH_IVX2 U20732 ( .A(n36470), .Z(n36471) );
  HS65_LH_BFX2 U20733 ( .A(n16032), .Z(n36472) );
  HS65_LH_IVX2 U20734 ( .A(n36466), .Z(n36473) );
  HS65_LH_IVX2 U20735 ( .A(n36473), .Z(n36474) );
  HS65_LH_BFX2 U20736 ( .A(n36476), .Z(n36475) );
  HS65_LH_BFX2 U20737 ( .A(n2405), .Z(n36476) );
  HS65_LH_BFX2 U20738 ( .A(n36479), .Z(n36477) );
  HS65_LH_BFX2 U20739 ( .A(n16022), .Z(n36478) );
  HS65_LH_BFX2 U20740 ( .A(n36480), .Z(n36479) );
  HS65_LH_BFX2 U20741 ( .A(n36481), .Z(n36480) );
  HS65_LH_BFX2 U20742 ( .A(n36482), .Z(n36481) );
  HS65_LH_BFX2 U20743 ( .A(n17950), .Z(n36482) );
  HS65_LH_BFX2 U20744 ( .A(n36486), .Z(n36483) );
  HS65_LH_BFX2 U20745 ( .A(n36491), .Z(n36484) );
  HS65_LH_IVX2 U20746 ( .A(n36495), .Z(n36485) );
  HS65_LH_IVX2 U20747 ( .A(n36485), .Z(n36486) );
  HS65_LH_BFX2 U20748 ( .A(n2430), .Z(n36487) );
  HS65_LH_NAND4ABX3 U20749 ( .A(n16011), .B(n16010), .C(n16009), .D(n16008), 
        .Z(n16014) );
  HS65_LH_BFX2 U20750 ( .A(n16014), .Z(n36488) );
  HS65_LH_BFX2 U20751 ( .A(n2429), .Z(n36489) );
  HS65_LH_IVX2 U20752 ( .A(n36499), .Z(n36490) );
  HS65_LH_IVX2 U20753 ( .A(n36490), .Z(n36491) );
  HS65_LH_BFX2 U20754 ( .A(n36487), .Z(n36492) );
  HS65_LH_IVX2 U20755 ( .A(n36501), .Z(n36493) );
  HS65_LH_IVX2 U20756 ( .A(n36493), .Z(n36494) );
  HS65_LH_BFX2 U20757 ( .A(n36497), .Z(n36495) );
  HS65_LH_IVX2 U20758 ( .A(n36503), .Z(n36496) );
  HS65_LH_IVX2 U20759 ( .A(n36496), .Z(n36497) );
  HS65_LH_IVX2 U20760 ( .A(n36505), .Z(n36498) );
  HS65_LH_IVX2 U20761 ( .A(n36498), .Z(n36499) );
  HS65_LH_IVX2 U20762 ( .A(n36507), .Z(n36500) );
  HS65_LH_IVX2 U20763 ( .A(n36500), .Z(n36501) );
  HS65_LH_IVX2 U20764 ( .A(n36509), .Z(n36502) );
  HS65_LH_IVX2 U20765 ( .A(n36502), .Z(n36503) );
  HS65_LH_IVX2 U20766 ( .A(n36511), .Z(n36504) );
  HS65_LH_IVX2 U20767 ( .A(n36504), .Z(n36505) );
  HS65_LH_IVX2 U20768 ( .A(n36513), .Z(n36506) );
  HS65_LH_IVX2 U20769 ( .A(n36506), .Z(n36507) );
  HS65_LH_IVX2 U20770 ( .A(n36515), .Z(n36508) );
  HS65_LH_IVX2 U20771 ( .A(n36508), .Z(n36509) );
  HS65_LH_IVX2 U20772 ( .A(n36517), .Z(n36510) );
  HS65_LH_IVX2 U20773 ( .A(n36510), .Z(n36511) );
  HS65_LH_IVX2 U20774 ( .A(n36519), .Z(n36512) );
  HS65_LH_IVX2 U20775 ( .A(n36512), .Z(n36513) );
  HS65_LH_IVX2 U20776 ( .A(n36521), .Z(n36514) );
  HS65_LH_IVX2 U20777 ( .A(n36514), .Z(n36515) );
  HS65_LH_IVX2 U20778 ( .A(n36523), .Z(n36516) );
  HS65_LH_IVX2 U20779 ( .A(n36516), .Z(n36517) );
  HS65_LH_IVX2 U20780 ( .A(n36525), .Z(n36518) );
  HS65_LH_IVX2 U20781 ( .A(n36518), .Z(n36519) );
  HS65_LH_IVX2 U20782 ( .A(n36527), .Z(n36520) );
  HS65_LH_IVX2 U20783 ( .A(n36520), .Z(n36521) );
  HS65_LH_IVX2 U20784 ( .A(n36529), .Z(n36522) );
  HS65_LH_IVX2 U20785 ( .A(n36522), .Z(n36523) );
  HS65_LH_IVX2 U20786 ( .A(n36531), .Z(n36524) );
  HS65_LH_IVX2 U20787 ( .A(n36524), .Z(n36525) );
  HS65_LH_IVX2 U20788 ( .A(n36533), .Z(n36526) );
  HS65_LH_IVX2 U20789 ( .A(n36526), .Z(n36527) );
  HS65_LH_IVX2 U20790 ( .A(n36535), .Z(n36528) );
  HS65_LH_IVX2 U20791 ( .A(n36528), .Z(n36529) );
  HS65_LH_IVX2 U20792 ( .A(n36542), .Z(n36530) );
  HS65_LH_IVX2 U20793 ( .A(n36530), .Z(n36531) );
  HS65_LH_IVX2 U20794 ( .A(n36537), .Z(n36532) );
  HS65_LH_IVX2 U20795 ( .A(n36532), .Z(n36533) );
  HS65_LH_IVX2 U20796 ( .A(n36540), .Z(n36534) );
  HS65_LH_IVX2 U20797 ( .A(n36534), .Z(n36535) );
  HS65_LH_IVX2 U20798 ( .A(n36547), .Z(n36536) );
  HS65_LH_IVX2 U20799 ( .A(n36536), .Z(n36537) );
  HS65_LH_BFX2 U20800 ( .A(n36492), .Z(n36538) );
  HS65_LH_IVX2 U20801 ( .A(n36544), .Z(n36539) );
  HS65_LH_IVX2 U20802 ( .A(n36539), .Z(n36540) );
  HS65_LH_IVX2 U20803 ( .A(n36546), .Z(n36541) );
  HS65_LH_IVX2 U20804 ( .A(n36541), .Z(n36542) );
  HS65_LH_IVX2 U20805 ( .A(n36549), .Z(n36543) );
  HS65_LH_IVX2 U20806 ( .A(n36543), .Z(n36544) );
  HS65_LH_IVX2 U20807 ( .A(n36551), .Z(n36545) );
  HS65_LH_IVX2 U20808 ( .A(n36545), .Z(n36546) );
  HS65_LH_BFX2 U20809 ( .A(n36552), .Z(n36547) );
  HS65_LH_IVX2 U20810 ( .A(n36554), .Z(n36548) );
  HS65_LH_IVX2 U20811 ( .A(n36548), .Z(n36549) );
  HS65_LH_IVX2 U20812 ( .A(n36556), .Z(n36550) );
  HS65_LH_IVX2 U20813 ( .A(n36550), .Z(n36551) );
  HS65_LH_BFX2 U20814 ( .A(n36557), .Z(n36552) );
  HS65_LH_IVX2 U20815 ( .A(n36559), .Z(n36553) );
  HS65_LH_IVX2 U20816 ( .A(n36553), .Z(n36554) );
  HS65_LH_IVX2 U20817 ( .A(n36538), .Z(n36555) );
  HS65_LH_IVX2 U20818 ( .A(n36555), .Z(n36556) );
  HS65_LH_BFX2 U20819 ( .A(n36562), .Z(n36557) );
  HS65_LH_IVX2 U20820 ( .A(n36489), .Z(n36558) );
  HS65_LH_IVX2 U20821 ( .A(n36558), .Z(n36559) );
  HS65_LH_IVX2 U20822 ( .A(n36560), .Z(n36561) );
  HS65_LH_BFX2 U20823 ( .A(n36564), .Z(n36562) );
  HS65_LH_BFX2 U20824 ( .A(n16013), .Z(n36563) );
  HS65_LH_BFX2 U20825 ( .A(n36565), .Z(n36564) );
  HS65_LH_BFX2 U20826 ( .A(n36566), .Z(n36565) );
  HS65_LH_BFX2 U20827 ( .A(n36567), .Z(n36566) );
  HS65_LH_BFX2 U20828 ( .A(n36568), .Z(n36567) );
  HS65_LH_BFX2 U20829 ( .A(n17981), .Z(n36568) );
  HS65_LH_BFX2 U20830 ( .A(n36577), .Z(n36569) );
  HS65_LH_IVX2 U20831 ( .A(n36570), .Z(n36571) );
  HS65_LH_IVX2 U20832 ( .A(n36579), .Z(n36572) );
  HS65_LH_IVX2 U20833 ( .A(n36572), .Z(n36573) );
  HS65_LH_IVX2 U20834 ( .A(n36581), .Z(n36574) );
  HS65_LH_IVX2 U20835 ( .A(n36574), .Z(n36575) );
  HS65_LH_IVX2 U20836 ( .A(n36582), .Z(n36576) );
  HS65_LH_IVX2 U20837 ( .A(n36576), .Z(n36577) );
  HS65_LH_IVX2 U20838 ( .A(n36586), .Z(n36578) );
  HS65_LH_IVX2 U20839 ( .A(n36578), .Z(n36579) );
  HS65_LH_IVX2 U20840 ( .A(n36588), .Z(n36580) );
  HS65_LH_IVX2 U20841 ( .A(n36580), .Z(n36581) );
  HS65_LH_BFX2 U20842 ( .A(n36584), .Z(n36582) );
  HS65_LH_IVX2 U20843 ( .A(n36590), .Z(n36583) );
  HS65_LH_IVX2 U20844 ( .A(n36583), .Z(n36584) );
  HS65_LH_IVX2 U20845 ( .A(n36592), .Z(n36585) );
  HS65_LH_IVX2 U20846 ( .A(n36585), .Z(n36586) );
  HS65_LH_IVX2 U20847 ( .A(n36594), .Z(n36587) );
  HS65_LH_IVX2 U20848 ( .A(n36587), .Z(n36588) );
  HS65_LH_IVX2 U20849 ( .A(n36596), .Z(n36589) );
  HS65_LH_IVX2 U20850 ( .A(n36589), .Z(n36590) );
  HS65_LH_IVX2 U20851 ( .A(n36598), .Z(n36591) );
  HS65_LH_IVX2 U20852 ( .A(n36591), .Z(n36592) );
  HS65_LH_IVX2 U20853 ( .A(n36600), .Z(n36593) );
  HS65_LH_IVX2 U20854 ( .A(n36593), .Z(n36594) );
  HS65_LH_IVX2 U20855 ( .A(n36602), .Z(n36595) );
  HS65_LH_IVX2 U20856 ( .A(n36595), .Z(n36596) );
  HS65_LH_IVX2 U20857 ( .A(n36604), .Z(n36597) );
  HS65_LH_IVX2 U20858 ( .A(n36597), .Z(n36598) );
  HS65_LH_IVX2 U20859 ( .A(n36606), .Z(n36599) );
  HS65_LH_IVX2 U20860 ( .A(n36599), .Z(n36600) );
  HS65_LH_IVX2 U20861 ( .A(n36608), .Z(n36601) );
  HS65_LH_IVX2 U20862 ( .A(n36601), .Z(n36602) );
  HS65_LH_IVX2 U20863 ( .A(n36610), .Z(n36603) );
  HS65_LH_IVX2 U20864 ( .A(n36603), .Z(n36604) );
  HS65_LH_IVX2 U20865 ( .A(n36612), .Z(n36605) );
  HS65_LH_IVX2 U20866 ( .A(n36605), .Z(n36606) );
  HS65_LH_IVX2 U20867 ( .A(n36614), .Z(n36607) );
  HS65_LH_IVX2 U20868 ( .A(n36607), .Z(n36608) );
  HS65_LH_IVX2 U20869 ( .A(n36616), .Z(n36609) );
  HS65_LH_IVX2 U20870 ( .A(n36609), .Z(n36610) );
  HS65_LH_IVX2 U20871 ( .A(n36618), .Z(n36611) );
  HS65_LH_IVX2 U20872 ( .A(n36611), .Z(n36612) );
  HS65_LH_IVX2 U20873 ( .A(n36620), .Z(n36613) );
  HS65_LH_IVX2 U20874 ( .A(n36613), .Z(n36614) );
  HS65_LH_IVX2 U20875 ( .A(n36622), .Z(n36615) );
  HS65_LH_IVX2 U20876 ( .A(n36615), .Z(n36616) );
  HS65_LH_IVX2 U20877 ( .A(n36624), .Z(n36617) );
  HS65_LH_IVX2 U20878 ( .A(n36617), .Z(n36618) );
  HS65_LH_IVX2 U20879 ( .A(n36626), .Z(n36619) );
  HS65_LH_IVX2 U20880 ( .A(n36619), .Z(n36620) );
  HS65_LH_IVX2 U20881 ( .A(n36628), .Z(n36621) );
  HS65_LH_IVX2 U20882 ( .A(n36621), .Z(n36622) );
  HS65_LH_IVX2 U20883 ( .A(n36630), .Z(n36623) );
  HS65_LH_IVX2 U20884 ( .A(n36623), .Z(n36624) );
  HS65_LH_IVX2 U20885 ( .A(n36635), .Z(n36625) );
  HS65_LH_IVX2 U20886 ( .A(n36625), .Z(n36626) );
  HS65_LH_IVX2 U20887 ( .A(n36632), .Z(n36627) );
  HS65_LH_IVX2 U20888 ( .A(n36627), .Z(n36628) );
  HS65_LH_IVX2 U20889 ( .A(n36634), .Z(n36629) );
  HS65_LH_IVX2 U20890 ( .A(n36629), .Z(n36630) );
  HS65_LH_IVX2 U20891 ( .A(n36637), .Z(n36631) );
  HS65_LH_IVX2 U20892 ( .A(n36631), .Z(n36632) );
  HS65_LH_IVX2 U20893 ( .A(n36639), .Z(n36633) );
  HS65_LH_IVX2 U20894 ( .A(n36633), .Z(n36634) );
  HS65_LH_BFX2 U20895 ( .A(n36640), .Z(n36635) );
  HS65_LH_IVX2 U20896 ( .A(n36642), .Z(n36636) );
  HS65_LH_IVX2 U20897 ( .A(n36636), .Z(n36637) );
  HS65_LH_IVX2 U20898 ( .A(n36644), .Z(n36638) );
  HS65_LH_IVX2 U20899 ( .A(n36638), .Z(n36639) );
  HS65_LH_BFX2 U20900 ( .A(n36645), .Z(n36640) );
  HS65_LH_IVX2 U20901 ( .A(n36648), .Z(n36641) );
  HS65_LH_IVX2 U20902 ( .A(n36641), .Z(n36642) );
  HS65_LH_IVX2 U20903 ( .A(n2382), .Z(n36643) );
  HS65_LH_IVX2 U20904 ( .A(n36643), .Z(n36644) );
  HS65_LH_BFX2 U20905 ( .A(n36651), .Z(n36645) );
  HS65_LH_BFX2 U20906 ( .A(n16042), .Z(n36646) );
  HS65_LH_IVX2 U20907 ( .A(n2381), .Z(n36647) );
  HS65_LH_IVX2 U20908 ( .A(n36647), .Z(n36648) );
  HS65_LH_IVX2 U20909 ( .A(n16053), .Z(n36649) );
  HS65_LH_IVX2 U20910 ( .A(n36649), .Z(n36650) );
  HS65_LH_BFX2 U20911 ( .A(n36652), .Z(n36651) );
  HS65_LH_BFX2 U20912 ( .A(n36653), .Z(n36652) );
  HS65_LH_BFX2 U20913 ( .A(n36654), .Z(n36653) );
  HS65_LH_BFX2 U20914 ( .A(n36655), .Z(n36654) );
  HS65_LH_BFX2 U20915 ( .A(n36656), .Z(n36655) );
  HS65_LH_BFX2 U20916 ( .A(n17944), .Z(n36656) );
  HS65_LH_BFX2 U20917 ( .A(n36660), .Z(n36657) );
  HS65_LH_BFX2 U20918 ( .A(n36661), .Z(n36658) );
  HS65_LH_BFX2 U20919 ( .A(n2526), .Z(n36659) );
  HS65_LH_BFX2 U20920 ( .A(n36663), .Z(n36660) );
  HS65_LH_BFX2 U20921 ( .A(n36664), .Z(n36661) );
  HS65_LH_BFX2 U20922 ( .A(n36659), .Z(n36662) );
  HS65_LH_BFX2 U20923 ( .A(n36666), .Z(n36663) );
  HS65_LH_BFX2 U20924 ( .A(n36667), .Z(n36664) );
  HS65_LH_BFX2 U20925 ( .A(n36662), .Z(n36665) );
  HS65_LH_BFX2 U20926 ( .A(n36669), .Z(n36666) );
  HS65_LH_BFX2 U20927 ( .A(n36670), .Z(n36667) );
  HS65_LH_BFX2 U20928 ( .A(n36665), .Z(n36668) );
  HS65_LH_BFX2 U20929 ( .A(n36672), .Z(n36669) );
  HS65_LH_BFX2 U20930 ( .A(n36673), .Z(n36670) );
  HS65_LH_BFX2 U20931 ( .A(n36668), .Z(n36671) );
  HS65_LH_BFX2 U20932 ( .A(n36675), .Z(n36672) );
  HS65_LH_BFX2 U20933 ( .A(n36676), .Z(n36673) );
  HS65_LH_BFX2 U20934 ( .A(n36671), .Z(n36674) );
  HS65_LH_BFX2 U20935 ( .A(n36678), .Z(n36675) );
  HS65_LH_BFX2 U20936 ( .A(n36679), .Z(n36676) );
  HS65_LH_BFX2 U20937 ( .A(n36674), .Z(n36677) );
  HS65_LH_BFX2 U20938 ( .A(n36681), .Z(n36678) );
  HS65_LH_BFX2 U20939 ( .A(n36682), .Z(n36679) );
  HS65_LH_BFX2 U20940 ( .A(n36677), .Z(n36680) );
  HS65_LH_BFX2 U20941 ( .A(n36684), .Z(n36681) );
  HS65_LH_BFX2 U20942 ( .A(n36685), .Z(n36682) );
  HS65_LH_BFX2 U20943 ( .A(n36680), .Z(n36683) );
  HS65_LH_BFX2 U20944 ( .A(n36687), .Z(n36684) );
  HS65_LH_BFX2 U20945 ( .A(n36688), .Z(n36685) );
  HS65_LH_BFX2 U20946 ( .A(n36683), .Z(n36686) );
  HS65_LH_BFX2 U20947 ( .A(n36690), .Z(n36687) );
  HS65_LH_BFX2 U20948 ( .A(n36691), .Z(n36688) );
  HS65_LH_BFX2 U20949 ( .A(n36686), .Z(n36689) );
  HS65_LH_BFX2 U20950 ( .A(n36693), .Z(n36690) );
  HS65_LH_BFX2 U20951 ( .A(n36694), .Z(n36691) );
  HS65_LH_BFX2 U20952 ( .A(n36689), .Z(n36692) );
  HS65_LH_BFX2 U20953 ( .A(n36699), .Z(n36693) );
  HS65_LH_BFX2 U20954 ( .A(n36697), .Z(n36694) );
  HS65_LH_BFX2 U20955 ( .A(n15934), .Z(n36695) );
  HS65_LH_IVX2 U20956 ( .A(n36702), .Z(n36696) );
  HS65_LH_IVX2 U20957 ( .A(n36696), .Z(n36697) );
  HS65_LH_BFX2 U20958 ( .A(n15933), .Z(n36698) );
  HS65_LH_BFX2 U20959 ( .A(n36705), .Z(n36699) );
  HS65_LH_BFX2 U20960 ( .A(n36692), .Z(n36700) );
  HS65_LH_IVX2 U20961 ( .A(n36707), .Z(n36701) );
  HS65_LH_IVX2 U20962 ( .A(n36701), .Z(n36702) );
  HS65_LH_IVX2 U20963 ( .A(n36700), .Z(n36703) );
  HS65_LH_IVX2 U20964 ( .A(n36703), .Z(n36704) );
  HS65_LH_BFX2 U20965 ( .A(n36706), .Z(n36705) );
  HS65_LH_BFX2 U20966 ( .A(n2525), .Z(n36706) );
  HS65_LH_BFX2 U20967 ( .A(n36708), .Z(n36707) );
  HS65_LH_BFX2 U20968 ( .A(n36709), .Z(n36708) );
  HS65_LH_BFX2 U20969 ( .A(n36710), .Z(n36709) );
  HS65_LH_BFX2 U20970 ( .A(n36711), .Z(n36710) );
  HS65_LH_BFX2 U20971 ( .A(n17947), .Z(n36711) );
  HS65_LH_BFX2 U20972 ( .A(n36761), .Z(n36712) );
  HS65_LH_BFX2 U20973 ( .A(n2501), .Z(n36713) );
  HS65_LH_BFX2 U20974 ( .A(n36717), .Z(n36714) );
  HS65_LH_BFX2 U20975 ( .A(n2502), .Z(n36715) );
  HS65_LH_BFX2 U20976 ( .A(n36713), .Z(n36716) );
  HS65_LH_BFX2 U20977 ( .A(n36720), .Z(n36717) );
  HS65_LH_BFX2 U20978 ( .A(n36715), .Z(n36718) );
  HS65_LH_BFX2 U20979 ( .A(n36716), .Z(n36719) );
  HS65_LH_BFX2 U20980 ( .A(n36723), .Z(n36720) );
  HS65_LH_BFX2 U20981 ( .A(n36718), .Z(n36721) );
  HS65_LH_BFX2 U20982 ( .A(n36719), .Z(n36722) );
  HS65_LH_BFX2 U20983 ( .A(n36726), .Z(n36723) );
  HS65_LH_BFX2 U20984 ( .A(n36721), .Z(n36724) );
  HS65_LH_BFX2 U20985 ( .A(n36722), .Z(n36725) );
  HS65_LH_BFX2 U20986 ( .A(n36729), .Z(n36726) );
  HS65_LH_BFX2 U20987 ( .A(n36724), .Z(n36727) );
  HS65_LH_BFX2 U20988 ( .A(n36725), .Z(n36728) );
  HS65_LH_BFX2 U20989 ( .A(n36732), .Z(n36729) );
  HS65_LH_BFX2 U20990 ( .A(n36727), .Z(n36730) );
  HS65_LH_BFX2 U20991 ( .A(n36728), .Z(n36731) );
  HS65_LH_BFX2 U20992 ( .A(n36735), .Z(n36732) );
  HS65_LH_BFX2 U20993 ( .A(n36730), .Z(n36733) );
  HS65_LH_BFX2 U20994 ( .A(n36731), .Z(n36734) );
  HS65_LH_BFX2 U20995 ( .A(n36738), .Z(n36735) );
  HS65_LH_BFX2 U20996 ( .A(n36733), .Z(n36736) );
  HS65_LH_BFX2 U20997 ( .A(n36734), .Z(n36737) );
  HS65_LH_BFX2 U20998 ( .A(n36741), .Z(n36738) );
  HS65_LH_BFX2 U20999 ( .A(n36736), .Z(n36739) );
  HS65_LH_BFX2 U21000 ( .A(n36737), .Z(n36740) );
  HS65_LH_BFX2 U21001 ( .A(n36744), .Z(n36741) );
  HS65_LH_BFX2 U21002 ( .A(n36739), .Z(n36742) );
  HS65_LH_BFX2 U21003 ( .A(n36740), .Z(n36743) );
  HS65_LH_BFX2 U21004 ( .A(n36747), .Z(n36744) );
  HS65_LH_BFX2 U21005 ( .A(n36742), .Z(n36745) );
  HS65_LH_BFX2 U21006 ( .A(n36743), .Z(n36746) );
  HS65_LH_BFX2 U21007 ( .A(n36750), .Z(n36747) );
  HS65_LH_BFX2 U21008 ( .A(n36745), .Z(n36748) );
  HS65_LH_BFX2 U21009 ( .A(n36746), .Z(n36749) );
  HS65_LH_BFX2 U21010 ( .A(n36753), .Z(n36750) );
  HS65_LH_BFX2 U21011 ( .A(n36748), .Z(n36751) );
  HS65_LH_BFX2 U21012 ( .A(n36749), .Z(n36752) );
  HS65_LH_BFX2 U21013 ( .A(n36762), .Z(n36753) );
  HS65_LH_BFX2 U21014 ( .A(n36751), .Z(n36754) );
  HS65_LH_BFX2 U21015 ( .A(n15942), .Z(n36755) );
  HS65_LH_IVX2 U21016 ( .A(n36752), .Z(n36756) );
  HS65_LH_IVX2 U21017 ( .A(n36756), .Z(n36757) );
  HS65_LH_IVX2 U21018 ( .A(n36758), .Z(n36759) );
  HS65_LH_IVX2 U21019 ( .A(n36754), .Z(n36760) );
  HS65_LH_IVX2 U21020 ( .A(n36760), .Z(n36761) );
  HS65_LH_BFX2 U21021 ( .A(n36763), .Z(n36762) );
  HS65_LH_BFX2 U21022 ( .A(n36764), .Z(n36763) );
  HS65_LH_BFX2 U21023 ( .A(n36765), .Z(n36764) );
  HS65_LH_BFX2 U21024 ( .A(n36766), .Z(n36765) );
  HS65_LH_BFX2 U21025 ( .A(n36767), .Z(n36766) );
  HS65_LH_BFX2 U21026 ( .A(n17898), .Z(n36767) );
  HS65_LH_BFX2 U21027 ( .A(n36771), .Z(n36768) );
  HS65_LH_BFX2 U21028 ( .A(n36772), .Z(n36769) );
  HS65_LH_BFX2 U21029 ( .A(n36773), .Z(n36770) );
  HS65_LH_BFX2 U21030 ( .A(n36774), .Z(n36771) );
  HS65_LH_BFX2 U21031 ( .A(n36775), .Z(n36772) );
  HS65_LH_BFX2 U21032 ( .A(n36776), .Z(n36773) );
  HS65_LH_BFX2 U21033 ( .A(n36777), .Z(n36774) );
  HS65_LH_BFX2 U21034 ( .A(n36778), .Z(n36775) );
  HS65_LH_BFX2 U21035 ( .A(n36779), .Z(n36776) );
  HS65_LH_BFX2 U21036 ( .A(n36780), .Z(n36777) );
  HS65_LH_BFX2 U21037 ( .A(n36781), .Z(n36778) );
  HS65_LH_BFX2 U21038 ( .A(n36782), .Z(n36779) );
  HS65_LH_BFX2 U21039 ( .A(n36783), .Z(n36780) );
  HS65_LH_BFX2 U21040 ( .A(n36784), .Z(n36781) );
  HS65_LH_BFX2 U21041 ( .A(n36785), .Z(n36782) );
  HS65_LH_BFX2 U21042 ( .A(n36786), .Z(n36783) );
  HS65_LH_BFX2 U21043 ( .A(n36787), .Z(n36784) );
  HS65_LH_BFX2 U21044 ( .A(n36788), .Z(n36785) );
  HS65_LH_BFX2 U21045 ( .A(n36789), .Z(n36786) );
  HS65_LH_BFX2 U21046 ( .A(n36790), .Z(n36787) );
  HS65_LH_BFX2 U21047 ( .A(n36791), .Z(n36788) );
  HS65_LH_BFX2 U21048 ( .A(n36792), .Z(n36789) );
  HS65_LH_BFX2 U21049 ( .A(n36793), .Z(n36790) );
  HS65_LH_BFX2 U21050 ( .A(n36794), .Z(n36791) );
  HS65_LH_BFX2 U21051 ( .A(n36795), .Z(n36792) );
  HS65_LH_BFX2 U21052 ( .A(n36796), .Z(n36793) );
  HS65_LH_BFX2 U21053 ( .A(n36797), .Z(n36794) );
  HS65_LH_BFX2 U21054 ( .A(n36798), .Z(n36795) );
  HS65_LH_BFX2 U21055 ( .A(n36799), .Z(n36796) );
  HS65_LH_BFX2 U21056 ( .A(n36800), .Z(n36797) );
  HS65_LH_BFX2 U21057 ( .A(n36801), .Z(n36798) );
  HS65_LH_BFX2 U21058 ( .A(n36802), .Z(n36799) );
  HS65_LH_BFX2 U21059 ( .A(n36803), .Z(n36800) );
  HS65_LH_BFX2 U21060 ( .A(n36804), .Z(n36801) );
  HS65_LH_BFX2 U21061 ( .A(n36805), .Z(n36802) );
  HS65_LH_BFX2 U21062 ( .A(n36806), .Z(n36803) );
  HS65_LH_BFX2 U21063 ( .A(n36807), .Z(n36804) );
  HS65_LH_BFX2 U21064 ( .A(n36808), .Z(n36805) );
  HS65_LH_BFX2 U21065 ( .A(n36809), .Z(n36806) );
  HS65_LH_BFX2 U21066 ( .A(n36810), .Z(n36807) );
  HS65_LH_BFX2 U21067 ( .A(n36811), .Z(n36808) );
  HS65_LH_BFX2 U21068 ( .A(n36812), .Z(n36809) );
  HS65_LH_BFX2 U21069 ( .A(n36813), .Z(n36810) );
  HS65_LH_BFX2 U21070 ( .A(n36814), .Z(n36811) );
  HS65_LH_BFX2 U21071 ( .A(n36815), .Z(n36812) );
  HS65_LH_BFX2 U21072 ( .A(n2453), .Z(n36813) );
  HS65_LH_BFX2 U21073 ( .A(n2454), .Z(n36814) );
  HS65_LH_BFX2 U21074 ( .A(n36816), .Z(n36815) );
  HS65_LH_BFX2 U21075 ( .A(n36817), .Z(n36816) );
  HS65_LH_BFX2 U21076 ( .A(n36818), .Z(n36817) );
  HS65_LH_BFX2 U21077 ( .A(n36819), .Z(n36818) );
  HS65_LH_BFX2 U21078 ( .A(n17969), .Z(n36819) );
  HS65_LH_IVX2 U21079 ( .A(n36831), .Z(n36820) );
  HS65_LH_IVX2 U21080 ( .A(n36820), .Z(n36821) );
  HS65_LH_BFX2 U21081 ( .A(n36825), .Z(n36822) );
  HS65_LH_BFX2 U21082 ( .A(n2094), .Z(n36823) );
  HS65_LH_IVX2 U21083 ( .A(n36830), .Z(n36824) );
  HS65_LH_IVX2 U21084 ( .A(n36824), .Z(n36825) );
  HS65_LH_BFX2 U21085 ( .A(n36823), .Z(n36826) );
  HS65_LH_IVX2 U21086 ( .A(n36833), .Z(n36827) );
  HS65_LH_IVX2 U21087 ( .A(n36827), .Z(n36828) );
  HS65_LH_IVX2 U21088 ( .A(n36920), .Z(n36829) );
  HS65_LH_IVX2 U21089 ( .A(n36829), .Z(n36830) );
  HS65_LH_BFX2 U21090 ( .A(n36832), .Z(n36831) );
  HS65_LH_BFX2 U21091 ( .A(n36835), .Z(n36832) );
  HS65_LH_BFX2 U21092 ( .A(n36836), .Z(n36833) );
  HS65_LH_BFX2 U21093 ( .A(n36189), .Z(n36834) );
  HS65_LH_BFX2 U21094 ( .A(n36861), .Z(n36835) );
  HS65_LH_BFX2 U21095 ( .A(n36839), .Z(n36836) );
  HS65_LH_BFX2 U21096 ( .A(n36834), .Z(n36837) );
  HS65_LH_IVX2 U21097 ( .A(n36842), .Z(n36838) );
  HS65_LH_IVX2 U21098 ( .A(n36838), .Z(n36839) );
  HS65_LH_BFX2 U21099 ( .A(n2093), .Z(n36840) );
  HS65_LH_BFX2 U21100 ( .A(n36840), .Z(n36841) );
  HS65_LH_BFX2 U21101 ( .A(n36844), .Z(n36842) );
  HS65_LH_BFX2 U21102 ( .A(n36841), .Z(n36843) );
  HS65_LH_BFX2 U21103 ( .A(n36846), .Z(n36844) );
  HS65_LH_BFX2 U21104 ( .A(n36843), .Z(n36845) );
  HS65_LH_BFX2 U21105 ( .A(n36848), .Z(n36846) );
  HS65_LH_BFX2 U21106 ( .A(n36845), .Z(n36847) );
  HS65_LH_BFX2 U21107 ( .A(n36850), .Z(n36848) );
  HS65_LH_BFX2 U21108 ( .A(n36847), .Z(n36849) );
  HS65_LH_BFX2 U21109 ( .A(n36852), .Z(n36850) );
  HS65_LH_BFX2 U21110 ( .A(n36849), .Z(n36851) );
  HS65_LH_BFX2 U21111 ( .A(n36854), .Z(n36852) );
  HS65_LH_BFX2 U21112 ( .A(n36851), .Z(n36853) );
  HS65_LH_BFX2 U21113 ( .A(n36856), .Z(n36854) );
  HS65_LH_BFX2 U21114 ( .A(n36853), .Z(n36855) );
  HS65_LH_BFX2 U21115 ( .A(n36859), .Z(n36856) );
  HS65_LH_BFX2 U21116 ( .A(n16285), .Z(n36857) );
  HS65_LH_IVX2 U21117 ( .A(n36826), .Z(n36858) );
  HS65_LH_IVX2 U21118 ( .A(n36858), .Z(n36859) );
  HS65_LH_IVX2 U21119 ( .A(n36855), .Z(n36860) );
  HS65_LH_IVX2 U21120 ( .A(n36860), .Z(n36861) );
  HS65_LH_BFX2 U21121 ( .A(n36865), .Z(n36862) );
  HS65_LH_BFX2 U21122 ( .A(n36866), .Z(n36863) );
  HS65_LH_BFX2 U21123 ( .A(n37125), .Z(n36864) );
  HS65_LH_BFX2 U21124 ( .A(n36867), .Z(n36865) );
  HS65_LH_BFX2 U21125 ( .A(n36868), .Z(n36866) );
  HS65_LH_BFX2 U21126 ( .A(n36869), .Z(n36867) );
  HS65_LH_BFX2 U21127 ( .A(n36870), .Z(n36868) );
  HS65_LH_BFX2 U21128 ( .A(n36871), .Z(n36869) );
  HS65_LH_BFX2 U21129 ( .A(n36872), .Z(n36870) );
  HS65_LH_BFX2 U21130 ( .A(n36873), .Z(n36871) );
  HS65_LH_BFX2 U21131 ( .A(n36874), .Z(n36872) );
  HS65_LH_BFX2 U21132 ( .A(n36875), .Z(n36873) );
  HS65_LH_BFX2 U21133 ( .A(n36876), .Z(n36874) );
  HS65_LH_BFX2 U21134 ( .A(n36877), .Z(n36875) );
  HS65_LH_BFX2 U21135 ( .A(n36878), .Z(n36876) );
  HS65_LH_BFX2 U21136 ( .A(n36879), .Z(n36877) );
  HS65_LH_BFX2 U21137 ( .A(n36880), .Z(n36878) );
  HS65_LH_BFX2 U21138 ( .A(n36881), .Z(n36879) );
  HS65_LH_BFX2 U21139 ( .A(n36882), .Z(n36880) );
  HS65_LH_BFX2 U21140 ( .A(n36883), .Z(n36881) );
  HS65_LH_BFX2 U21141 ( .A(n36884), .Z(n36882) );
  HS65_LH_BFX2 U21142 ( .A(n36885), .Z(n36883) );
  HS65_LH_BFX2 U21143 ( .A(n36886), .Z(n36884) );
  HS65_LH_BFX2 U21144 ( .A(n36887), .Z(n36885) );
  HS65_LH_BFX2 U21145 ( .A(n36888), .Z(n36886) );
  HS65_LH_BFX2 U21146 ( .A(n36889), .Z(n36887) );
  HS65_LH_BFX2 U21147 ( .A(n36890), .Z(n36888) );
  HS65_LH_BFX2 U21148 ( .A(n36891), .Z(n36889) );
  HS65_LH_BFX2 U21149 ( .A(n36892), .Z(n36890) );
  HS65_LH_BFX2 U21150 ( .A(n36893), .Z(n36891) );
  HS65_LH_BFX2 U21151 ( .A(n36894), .Z(n36892) );
  HS65_LH_BFX2 U21152 ( .A(n2262), .Z(n36893) );
  HS65_LH_BFX2 U21153 ( .A(n2261), .Z(n36894) );
  HS65_LH_BFX2 U21154 ( .A(n36898), .Z(n36895) );
  HS65_LH_BFX2 U21155 ( .A(n36900), .Z(n36896) );
  HS65_LH_IVX2 U21156 ( .A(n36903), .Z(n36897) );
  HS65_LH_IVX2 U21157 ( .A(n36897), .Z(n36898) );
  HS65_LH_IVX2 U21158 ( .A(n36905), .Z(n36899) );
  HS65_LH_IVX2 U21159 ( .A(n36899), .Z(n36900) );
  HS65_LH_BFX2 U21160 ( .A(n1949), .Z(n36901) );
  HS65_LH_IVX2 U21161 ( .A(n36908), .Z(n36902) );
  HS65_LH_IVX2 U21162 ( .A(n36902), .Z(n36903) );
  HS65_LH_IVX2 U21163 ( .A(n36910), .Z(n36904) );
  HS65_LH_IVX2 U21164 ( .A(n36904), .Z(n36905) );
  HS65_LH_BFX2 U21165 ( .A(n36901), .Z(n36906) );
  HS65_LH_IVX2 U21166 ( .A(n36913), .Z(n36907) );
  HS65_LH_IVX2 U21167 ( .A(n36907), .Z(n36908) );
  HS65_LH_IVX2 U21168 ( .A(n36915), .Z(n36909) );
  HS65_LH_IVX2 U21169 ( .A(n36909), .Z(n36910) );
  HS65_LH_BFX2 U21170 ( .A(n36906), .Z(n36911) );
  HS65_LH_IVX2 U21171 ( .A(n36939), .Z(n36912) );
  HS65_LH_IVX2 U21172 ( .A(n36912), .Z(n36913) );
  HS65_LH_IVX2 U21173 ( .A(n36922), .Z(n36914) );
  HS65_LH_IVX2 U21174 ( .A(n36914), .Z(n36915) );
  HS65_LH_IVX2 U21175 ( .A(n36935), .Z(n36916) );
  HS65_LH_IVX2 U21176 ( .A(n36916), .Z(n36917) );
  HS65_LH_BFX2 U21177 ( .A(n36911), .Z(n36918) );
  HS65_LH_IVX2 U21178 ( .A(n36895), .Z(n36919) );
  HS65_LH_IVX2 U21179 ( .A(n36919), .Z(n36920) );
  HS65_LH_IVX2 U21180 ( .A(n36927), .Z(n36921) );
  HS65_LH_IVX2 U21181 ( .A(n36921), .Z(n36922) );
  HS65_LH_IVX2 U21182 ( .A(n36930), .Z(n36923) );
  HS65_LH_IVX2 U21183 ( .A(n36923), .Z(n36924) );
  HS65_LH_BFX2 U21184 ( .A(n36918), .Z(n36925) );
  HS65_LH_IVX2 U21185 ( .A(n36932), .Z(n36926) );
  HS65_LH_IVX2 U21186 ( .A(n36926), .Z(n36927) );
  HS65_LH_BFX2 U21187 ( .A(n36925), .Z(n36928) );
  HS65_LH_IVX2 U21188 ( .A(n36917), .Z(n36929) );
  HS65_LH_IVX2 U21189 ( .A(n36929), .Z(n36930) );
  HS65_LH_BFX2 U21190 ( .A(n36928), .Z(n36931) );
  HS65_LH_BFX2 U21191 ( .A(n36936), .Z(n36932) );
  HS65_LH_BFX2 U21192 ( .A(n36931), .Z(n36933) );
  HS65_LH_IVX2 U21193 ( .A(n36941), .Z(n36934) );
  HS65_LH_IVX2 U21194 ( .A(n36934), .Z(n36935) );
  HS65_LH_BFX2 U21195 ( .A(n36942), .Z(n36936) );
  HS65_LH_BFX2 U21196 ( .A(n36933), .Z(n36937) );
  HS65_LH_IVX2 U21197 ( .A(n36948), .Z(n36938) );
  HS65_LH_IVX2 U21198 ( .A(n36938), .Z(n36939) );
  HS65_LH_IVX2 U21199 ( .A(n36895), .Z(n36940) );
  HS65_LH_IVX2 U21200 ( .A(n36940), .Z(n36941) );
  HS65_LH_BFX2 U21201 ( .A(n36944), .Z(n36942) );
  HS65_LH_BFX2 U21202 ( .A(n36937), .Z(n36943) );
  HS65_LH_BFX2 U21203 ( .A(n36946), .Z(n36944) );
  HS65_LH_BFX2 U21204 ( .A(n36943), .Z(n36945) );
  HS65_LH_BFX2 U21205 ( .A(n36952), .Z(n36946) );
  HS65_LH_BFX2 U21206 ( .A(n36945), .Z(n36947) );
  HS65_LH_BFX2 U21207 ( .A(n36837), .Z(n36948) );
  HS65_LH_BFX2 U21208 ( .A(n1950), .Z(n36949) );
  HS65_LH_BFX2 U21209 ( .A(n36947), .Z(n36950) );
  HS65_LH_IVX2 U21210 ( .A(n36957), .Z(n36951) );
  HS65_LH_IVX2 U21211 ( .A(n36951), .Z(n36952) );
  HS65_LH_BFX2 U21212 ( .A(n36950), .Z(n36953) );
  HS65_LH_IVX2 U21213 ( .A(n36953), .Z(n36954) );
  HS65_LH_IVX2 U21214 ( .A(n36954), .Z(n36955) );
  HS65_LH_IVX2 U21215 ( .A(n36949), .Z(n36956) );
  HS65_LH_IVX2 U21216 ( .A(n36956), .Z(n36957) );
  HS65_LH_BFX2 U21217 ( .A(n17419), .Z(n36958) );
  HS65_LH_BFX2 U21218 ( .A(n36960), .Z(n36959) );
  HS65_LH_BFX2 U21219 ( .A(n36961), .Z(n36960) );
  HS65_LH_BFX2 U21220 ( .A(n36962), .Z(n36961) );
  HS65_LH_BFX2 U21221 ( .A(n36963), .Z(n36962) );
  HS65_LH_BFX2 U21222 ( .A(n36964), .Z(n36963) );
  HS65_LH_BFX2 U21223 ( .A(n36965), .Z(n36964) );
  HS65_LH_BFX2 U21224 ( .A(n36966), .Z(n36965) );
  HS65_LH_BFX2 U21225 ( .A(n36967), .Z(n36966) );
  HS65_LH_BFX2 U21226 ( .A(n36968), .Z(n36967) );
  HS65_LH_BFX2 U21227 ( .A(n36969), .Z(n36968) );
  HS65_LH_BFX2 U21228 ( .A(n36970), .Z(n36969) );
  HS65_LH_BFX2 U21229 ( .A(n36971), .Z(n36970) );
  HS65_LH_BFX2 U21230 ( .A(n36972), .Z(n36971) );
  HS65_LH_BFX2 U21231 ( .A(n36973), .Z(n36972) );
  HS65_LH_BFX2 U21232 ( .A(n36974), .Z(n36973) );
  HS65_LH_BFX2 U21233 ( .A(n36975), .Z(n36974) );
  HS65_LH_BFX2 U21234 ( .A(n17780), .Z(n36975) );
  HS65_LH_BFX2 U21235 ( .A(n40160), .Z(n36976) );
  HS65_LH_BFX2 U21236 ( .A(n36980), .Z(n36977) );
  HS65_LH_BFX2 U21237 ( .A(n36981), .Z(n36978) );
  HS65_LH_BFX2 U21238 ( .A(n30897), .Z(n36979) );
  HS65_LH_BFX2 U21239 ( .A(n36983), .Z(n36980) );
  HS65_LH_BFX2 U21240 ( .A(n36984), .Z(n36981) );
  HS65_LH_BFX2 U21241 ( .A(n36979), .Z(n36982) );
  HS65_LH_BFX2 U21242 ( .A(n36986), .Z(n36983) );
  HS65_LH_BFX2 U21243 ( .A(n36987), .Z(n36984) );
  HS65_LH_BFX2 U21244 ( .A(n36982), .Z(n36985) );
  HS65_LH_BFX2 U21245 ( .A(n36989), .Z(n36986) );
  HS65_LH_BFX2 U21246 ( .A(n36990), .Z(n36987) );
  HS65_LH_BFX2 U21247 ( .A(n36985), .Z(n36988) );
  HS65_LH_BFX2 U21248 ( .A(n36992), .Z(n36989) );
  HS65_LH_BFX2 U21249 ( .A(n36993), .Z(n36990) );
  HS65_LH_BFX2 U21250 ( .A(n36988), .Z(n36991) );
  HS65_LH_BFX2 U21251 ( .A(n36995), .Z(n36992) );
  HS65_LH_BFX2 U21252 ( .A(n36996), .Z(n36993) );
  HS65_LH_BFX2 U21253 ( .A(n36991), .Z(n36994) );
  HS65_LH_BFX2 U21254 ( .A(n36998), .Z(n36995) );
  HS65_LH_BFX2 U21255 ( .A(n36999), .Z(n36996) );
  HS65_LH_BFX2 U21256 ( .A(n36994), .Z(n36997) );
  HS65_LH_BFX2 U21257 ( .A(n37001), .Z(n36998) );
  HS65_LH_BFX2 U21258 ( .A(n37002), .Z(n36999) );
  HS65_LH_BFX2 U21259 ( .A(n36997), .Z(n37000) );
  HS65_LH_BFX2 U21260 ( .A(n37004), .Z(n37001) );
  HS65_LH_BFX2 U21261 ( .A(n37005), .Z(n37002) );
  HS65_LH_BFX2 U21262 ( .A(n37000), .Z(n37003) );
  HS65_LH_BFX2 U21263 ( .A(n37007), .Z(n37004) );
  HS65_LH_BFX2 U21264 ( .A(n37008), .Z(n37005) );
  HS65_LH_BFX2 U21265 ( .A(n37003), .Z(n37006) );
  HS65_LH_BFX2 U21266 ( .A(n37010), .Z(n37007) );
  HS65_LH_BFX2 U21267 ( .A(n37011), .Z(n37008) );
  HS65_LH_BFX2 U21268 ( .A(n37006), .Z(n37009) );
  HS65_LH_BFX2 U21269 ( .A(n37013), .Z(n37010) );
  HS65_LH_BFX2 U21270 ( .A(n37014), .Z(n37011) );
  HS65_LH_BFX2 U21271 ( .A(n37009), .Z(n37012) );
  HS65_LH_BFX2 U21272 ( .A(n37016), .Z(n37013) );
  HS65_LH_BFX2 U21273 ( .A(n37017), .Z(n37014) );
  HS65_LH_BFX2 U21274 ( .A(n37012), .Z(n37015) );
  HS65_LH_BFX2 U21275 ( .A(n37019), .Z(n37016) );
  HS65_LH_BFX2 U21276 ( .A(n37020), .Z(n37017) );
  HS65_LH_BFX2 U21277 ( .A(n37015), .Z(n37018) );
  HS65_LH_BFX2 U21278 ( .A(n37022), .Z(n37019) );
  HS65_LH_BFX2 U21279 ( .A(n37023), .Z(n37020) );
  HS65_LH_BFX2 U21280 ( .A(n37018), .Z(n37021) );
  HS65_LH_BFX2 U21281 ( .A(n37025), .Z(n37022) );
  HS65_LH_BFX2 U21282 ( .A(n37026), .Z(n37023) );
  HS65_LH_BFX2 U21283 ( .A(n37021), .Z(n37024) );
  HS65_LH_BFX2 U21284 ( .A(n37028), .Z(n37025) );
  HS65_LH_BFX2 U21285 ( .A(n37029), .Z(n37026) );
  HS65_LH_BFX2 U21286 ( .A(n37024), .Z(n37027) );
  HS65_LH_BFX2 U21287 ( .A(n37035), .Z(n37028) );
  HS65_LH_BFX2 U21288 ( .A(n37032), .Z(n37029) );
  HS65_LH_BFX2 U21289 ( .A(n37027), .Z(n37030) );
  HS65_LH_IVX2 U21290 ( .A(n18041), .Z(n37031) );
  HS65_LH_IVX2 U21291 ( .A(n37031), .Z(n37032) );
  HS65_LH_IVX2 U21292 ( .A(n37030), .Z(n37033) );
  HS65_LH_IVX2 U21293 ( .A(n37033), .Z(n37034) );
  HS65_LH_BFX2 U21294 ( .A(n14099), .Z(n37035) );
  HS65_LH_BFX2 U21295 ( .A(n37037), .Z(n37036) );
  HS65_LH_BFX2 U21296 ( .A(n37038), .Z(n37037) );
  HS65_LH_BFX2 U21297 ( .A(n37039), .Z(n37038) );
  HS65_LH_BFX2 U21298 ( .A(n37040), .Z(n37039) );
  HS65_LH_BFX2 U21299 ( .A(n37041), .Z(n37040) );
  HS65_LH_BFX2 U21300 ( .A(n37042), .Z(n37041) );
  HS65_LH_BFX2 U21301 ( .A(n37043), .Z(n37042) );
  HS65_LH_BFX2 U21302 ( .A(n37044), .Z(n37043) );
  HS65_LH_BFX2 U21303 ( .A(n37045), .Z(n37044) );
  HS65_LH_BFX2 U21304 ( .A(n37046), .Z(n37045) );
  HS65_LH_BFX2 U21305 ( .A(n37048), .Z(n37046) );
  HS65_LH_BFX2 U21306 ( .A(n17647), .Z(n37047) );
  HS65_LH_BFX2 U21307 ( .A(n37049), .Z(n37048) );
  HS65_LH_BFX2 U21308 ( .A(n15491), .Z(n37049) );
  HS65_LH_BFX2 U21309 ( .A(n37051), .Z(n37050) );
  HS65_LH_BFX2 U21310 ( .A(n37052), .Z(n37051) );
  HS65_LH_BFX2 U21311 ( .A(n37053), .Z(n37052) );
  HS65_LH_BFX2 U21312 ( .A(n37054), .Z(n37053) );
  HS65_LH_BFX2 U21313 ( .A(n37055), .Z(n37054) );
  HS65_LH_BFX2 U21314 ( .A(n37056), .Z(n37055) );
  HS65_LH_BFX2 U21315 ( .A(n37057), .Z(n37056) );
  HS65_LH_BFX2 U21316 ( .A(n37058), .Z(n37057) );
  HS65_LH_BFX2 U21317 ( .A(n37059), .Z(n37058) );
  HS65_LH_BFX2 U21318 ( .A(n37060), .Z(n37059) );
  HS65_LH_BFX2 U21319 ( .A(n37061), .Z(n37060) );
  HS65_LH_BFX2 U21320 ( .A(n37062), .Z(n37061) );
  HS65_LH_BFX2 U21321 ( .A(n37063), .Z(n37062) );
  HS65_LH_BFX2 U21322 ( .A(n37064), .Z(n37063) );
  HS65_LH_BFX2 U21323 ( .A(n37065), .Z(n37064) );
  HS65_LH_BFX2 U21324 ( .A(n37066), .Z(n37065) );
  HS65_LH_BFX2 U21325 ( .A(n37067), .Z(n37066) );
  HS65_LH_BFX2 U21326 ( .A(n37068), .Z(n37067) );
  HS65_LH_BFX2 U21327 ( .A(n37069), .Z(n37068) );
  HS65_LH_BFX2 U21328 ( .A(n40990), .Z(n37069) );
  HS65_LH_BFX2 U21329 ( .A(n17301), .Z(n37070) );
  HS65_LH_BFX2 U21330 ( .A(n37073), .Z(n37071) );
  HS65_LH_IVX2 U21331 ( .A(n37078), .Z(n37072) );
  HS65_LH_IVX2 U21332 ( .A(n37072), .Z(n37073) );
  HS65_LH_BFX2 U21333 ( .A(n37076), .Z(n37074) );
  HS65_LH_BFX2 U21334 ( .A(n37077), .Z(n37075) );
  HS65_LH_BFX2 U21335 ( .A(n37079), .Z(n37076) );
  HS65_LH_BFX2 U21336 ( .A(n37080), .Z(n37077) );
  HS65_LH_BFX2 U21337 ( .A(n37081), .Z(n37078) );
  HS65_LH_BFX2 U21338 ( .A(n37082), .Z(n37079) );
  HS65_LH_BFX2 U21339 ( .A(n37083), .Z(n37080) );
  HS65_LH_BFX2 U21340 ( .A(n37084), .Z(n37081) );
  HS65_LH_BFX2 U21341 ( .A(n37085), .Z(n37082) );
  HS65_LH_BFX2 U21342 ( .A(n37086), .Z(n37083) );
  HS65_LH_BFX2 U21343 ( .A(n37087), .Z(n37084) );
  HS65_LH_BFX2 U21344 ( .A(n37088), .Z(n37085) );
  HS65_LH_BFX2 U21345 ( .A(n37089), .Z(n37086) );
  HS65_LH_BFX2 U21346 ( .A(n37090), .Z(n37087) );
  HS65_LH_BFX2 U21347 ( .A(n37091), .Z(n37088) );
  HS65_LH_BFX2 U21348 ( .A(n37092), .Z(n37089) );
  HS65_LH_BFX2 U21349 ( .A(n37093), .Z(n37090) );
  HS65_LH_BFX2 U21350 ( .A(n37094), .Z(n37091) );
  HS65_LH_BFX2 U21351 ( .A(n37095), .Z(n37092) );
  HS65_LH_BFX2 U21352 ( .A(n37096), .Z(n37093) );
  HS65_LH_BFX2 U21353 ( .A(n37097), .Z(n37094) );
  HS65_LH_BFX2 U21354 ( .A(n37098), .Z(n37095) );
  HS65_LH_BFX2 U21355 ( .A(n37099), .Z(n37096) );
  HS65_LH_BFX2 U21356 ( .A(n37100), .Z(n37097) );
  HS65_LH_BFX2 U21357 ( .A(n37101), .Z(n37098) );
  HS65_LH_BFX2 U21358 ( .A(n37102), .Z(n37099) );
  HS65_LH_BFX2 U21359 ( .A(n37103), .Z(n37100) );
  HS65_LH_BFX2 U21360 ( .A(n37104), .Z(n37101) );
  HS65_LH_BFX2 U21361 ( .A(n37105), .Z(n37102) );
  HS65_LH_BFX2 U21362 ( .A(n37106), .Z(n37103) );
  HS65_LH_BFX2 U21363 ( .A(n37107), .Z(n37104) );
  HS65_LH_BFX2 U21364 ( .A(n37108), .Z(n37105) );
  HS65_LH_BFX2 U21365 ( .A(n37109), .Z(n37106) );
  HS65_LH_BFX2 U21366 ( .A(n37110), .Z(n37107) );
  HS65_LH_BFX2 U21367 ( .A(n37111), .Z(n37108) );
  HS65_LH_BFX2 U21368 ( .A(n37112), .Z(n37109) );
  HS65_LH_BFX2 U21369 ( .A(n37113), .Z(n37110) );
  HS65_LH_BFX2 U21370 ( .A(n37114), .Z(n37111) );
  HS65_LH_BFX2 U21371 ( .A(n37118), .Z(n37112) );
  HS65_LH_BFX2 U21372 ( .A(n37116), .Z(n37113) );
  HS65_LH_BFX2 U21373 ( .A(n37117), .Z(n37114) );
  HS65_LH_BFX2 U21374 ( .A(n40987), .Z(n37115) );
  HS65_LH_BFX2 U21375 ( .A(n37119), .Z(n37116) );
  HS65_LH_BFX2 U21376 ( .A(n1473), .Z(n37117) );
  HS65_LH_BFX2 U21377 ( .A(n1472), .Z(n37118) );
  HS65_LH_BFX2 U21378 ( .A(n37120), .Z(n37119) );
  HS65_LH_BFX2 U21379 ( .A(n37121), .Z(n37120) );
  HS65_LH_BFX2 U21380 ( .A(n37122), .Z(n37121) );
  HS65_LH_BFX2 U21381 ( .A(n17885), .Z(n37122) );
  HS65_LH_IVX2 U21382 ( .A(n37132), .Z(n37123) );
  HS65_LH_IVX2 U21383 ( .A(n37123), .Z(n37124) );
  HS65_LH_BFX2 U21384 ( .A(n37128), .Z(n37125) );
  HS65_LH_BFX2 U21385 ( .A(n37130), .Z(n37126) );
  HS65_LH_IVX2 U21386 ( .A(n37134), .Z(n37127) );
  HS65_LH_IVX2 U21387 ( .A(n37127), .Z(n37128) );
  HS65_LH_IVX2 U21388 ( .A(n37136), .Z(n37129) );
  HS65_LH_IVX2 U21389 ( .A(n37129), .Z(n37130) );
  HS65_LH_IVX2 U21390 ( .A(n37138), .Z(n37131) );
  HS65_LH_IVX2 U21391 ( .A(n37131), .Z(n37132) );
  HS65_LH_IVX2 U21392 ( .A(n37140), .Z(n37133) );
  HS65_LH_IVX2 U21393 ( .A(n37133), .Z(n37134) );
  HS65_LH_IVX2 U21394 ( .A(n37142), .Z(n37135) );
  HS65_LH_IVX2 U21395 ( .A(n37135), .Z(n37136) );
  HS65_LH_IVX2 U21396 ( .A(n37144), .Z(n37137) );
  HS65_LH_IVX2 U21397 ( .A(n37137), .Z(n37138) );
  HS65_LH_IVX2 U21398 ( .A(n37146), .Z(n37139) );
  HS65_LH_IVX2 U21399 ( .A(n37139), .Z(n37140) );
  HS65_LH_IVX2 U21400 ( .A(n37148), .Z(n37141) );
  HS65_LH_IVX2 U21401 ( .A(n37141), .Z(n37142) );
  HS65_LH_IVX2 U21402 ( .A(n37150), .Z(n37143) );
  HS65_LH_IVX2 U21403 ( .A(n37143), .Z(n37144) );
  HS65_LH_IVX2 U21404 ( .A(n37152), .Z(n37145) );
  HS65_LH_IVX2 U21405 ( .A(n37145), .Z(n37146) );
  HS65_LH_IVX2 U21406 ( .A(n37154), .Z(n37147) );
  HS65_LH_IVX2 U21407 ( .A(n37147), .Z(n37148) );
  HS65_LH_IVX2 U21408 ( .A(n37156), .Z(n37149) );
  HS65_LH_IVX2 U21409 ( .A(n37149), .Z(n37150) );
  HS65_LH_IVX2 U21410 ( .A(n37158), .Z(n37151) );
  HS65_LH_IVX2 U21411 ( .A(n37151), .Z(n37152) );
  HS65_LH_IVX2 U21412 ( .A(n37160), .Z(n37153) );
  HS65_LH_IVX2 U21413 ( .A(n37153), .Z(n37154) );
  HS65_LH_IVX2 U21414 ( .A(n37162), .Z(n37155) );
  HS65_LH_IVX2 U21415 ( .A(n37155), .Z(n37156) );
  HS65_LH_IVX2 U21416 ( .A(n37164), .Z(n37157) );
  HS65_LH_IVX2 U21417 ( .A(n37157), .Z(n37158) );
  HS65_LH_IVX2 U21418 ( .A(n37166), .Z(n37159) );
  HS65_LH_IVX2 U21419 ( .A(n37159), .Z(n37160) );
  HS65_LH_IVX2 U21420 ( .A(n37168), .Z(n37161) );
  HS65_LH_IVX2 U21421 ( .A(n37161), .Z(n37162) );
  HS65_LH_IVX2 U21422 ( .A(n37170), .Z(n37163) );
  HS65_LH_IVX2 U21423 ( .A(n37163), .Z(n37164) );
  HS65_LH_IVX2 U21424 ( .A(n37172), .Z(n37165) );
  HS65_LH_IVX2 U21425 ( .A(n37165), .Z(n37166) );
  HS65_LH_IVX2 U21426 ( .A(n37174), .Z(n37167) );
  HS65_LH_IVX2 U21427 ( .A(n37167), .Z(n37168) );
  HS65_LH_IVX2 U21428 ( .A(n37176), .Z(n37169) );
  HS65_LH_IVX2 U21429 ( .A(n37169), .Z(n37170) );
  HS65_LH_IVX2 U21430 ( .A(n37178), .Z(n37171) );
  HS65_LH_IVX2 U21431 ( .A(n37171), .Z(n37172) );
  HS65_LH_IVX2 U21432 ( .A(n37180), .Z(n37173) );
  HS65_LH_IVX2 U21433 ( .A(n37173), .Z(n37174) );
  HS65_LH_IVX2 U21434 ( .A(n37182), .Z(n37175) );
  HS65_LH_IVX2 U21435 ( .A(n37175), .Z(n37176) );
  HS65_LH_IVX2 U21436 ( .A(n37184), .Z(n37177) );
  HS65_LH_IVX2 U21437 ( .A(n37177), .Z(n37178) );
  HS65_LH_IVX2 U21438 ( .A(n37186), .Z(n37179) );
  HS65_LH_IVX2 U21439 ( .A(n37179), .Z(n37180) );
  HS65_LH_IVX2 U21440 ( .A(n37188), .Z(n37181) );
  HS65_LH_IVX2 U21441 ( .A(n37181), .Z(n37182) );
  HS65_LH_IVX2 U21442 ( .A(n37190), .Z(n37183) );
  HS65_LH_IVX2 U21443 ( .A(n37183), .Z(n37184) );
  HS65_LH_IVX2 U21444 ( .A(n37192), .Z(n37185) );
  HS65_LH_IVX2 U21445 ( .A(n37185), .Z(n37186) );
  HS65_LH_IVX2 U21446 ( .A(n37197), .Z(n37187) );
  HS65_LH_IVX2 U21447 ( .A(n37187), .Z(n37188) );
  HS65_LH_IVX2 U21448 ( .A(n37194), .Z(n37189) );
  HS65_LH_IVX2 U21449 ( .A(n37189), .Z(n37190) );
  HS65_LH_IVX2 U21450 ( .A(n37196), .Z(n37191) );
  HS65_LH_IVX2 U21451 ( .A(n37191), .Z(n37192) );
  HS65_LH_IVX2 U21452 ( .A(n37199), .Z(n37193) );
  HS65_LH_IVX2 U21453 ( .A(n37193), .Z(n37194) );
  HS65_LH_IVX2 U21454 ( .A(n37201), .Z(n37195) );
  HS65_LH_IVX2 U21455 ( .A(n37195), .Z(n37196) );
  HS65_LH_BFX2 U21456 ( .A(n37202), .Z(n37197) );
  HS65_LH_IVX2 U21457 ( .A(n1449), .Z(n37198) );
  HS65_LH_IVX2 U21458 ( .A(n37198), .Z(n37199) );
  HS65_LH_IVX2 U21459 ( .A(n1450), .Z(n37200) );
  HS65_LH_IVX2 U21460 ( .A(n37200), .Z(n37201) );
  HS65_LH_BFX2 U21461 ( .A(n37203), .Z(n37202) );
  HS65_LH_BFX2 U21462 ( .A(n37204), .Z(n37203) );
  HS65_LH_BFX2 U21463 ( .A(n37205), .Z(n37204) );
  HS65_LH_BFX2 U21464 ( .A(n37206), .Z(n37205) );
  HS65_LH_BFX2 U21465 ( .A(n17875), .Z(n37206) );
  HS65_LH_BFX2 U21466 ( .A(n37209), .Z(n37207) );
  HS65_LH_BFX2 U21467 ( .A(n1748), .Z(n37208) );
  HS65_LH_BFX2 U21468 ( .A(n37212), .Z(n37209) );
  HS65_LH_BFX2 U21469 ( .A(n37208), .Z(n37210) );
  HS65_LH_BFX2 U21470 ( .A(n37214), .Z(n37211) );
  HS65_LH_BFX2 U21471 ( .A(n37215), .Z(n37212) );
  HS65_LH_BFX2 U21472 ( .A(n37210), .Z(n37213) );
  HS65_LH_BFX2 U21473 ( .A(n37217), .Z(n37214) );
  HS65_LH_BFX2 U21474 ( .A(n37218), .Z(n37215) );
  HS65_LH_BFX2 U21475 ( .A(n37213), .Z(n37216) );
  HS65_LH_BFX2 U21476 ( .A(n37220), .Z(n37217) );
  HS65_LH_BFX2 U21477 ( .A(n37221), .Z(n37218) );
  HS65_LH_BFX2 U21478 ( .A(n37216), .Z(n37219) );
  HS65_LH_BFX2 U21479 ( .A(n37223), .Z(n37220) );
  HS65_LH_BFX2 U21480 ( .A(n37224), .Z(n37221) );
  HS65_LH_BFX2 U21481 ( .A(n37219), .Z(n37222) );
  HS65_LH_BFX2 U21482 ( .A(n37226), .Z(n37223) );
  HS65_LH_BFX2 U21483 ( .A(n37227), .Z(n37224) );
  HS65_LH_BFX2 U21484 ( .A(n37222), .Z(n37225) );
  HS65_LH_BFX2 U21485 ( .A(n37229), .Z(n37226) );
  HS65_LH_BFX2 U21486 ( .A(n37230), .Z(n37227) );
  HS65_LH_BFX2 U21487 ( .A(n37225), .Z(n37228) );
  HS65_LH_BFX2 U21488 ( .A(n37232), .Z(n37229) );
  HS65_LH_BFX2 U21489 ( .A(n37233), .Z(n37230) );
  HS65_LH_BFX2 U21490 ( .A(n37228), .Z(n37231) );
  HS65_LH_BFX2 U21491 ( .A(n37235), .Z(n37232) );
  HS65_LH_BFX2 U21492 ( .A(n37236), .Z(n37233) );
  HS65_LH_BFX2 U21493 ( .A(n37231), .Z(n37234) );
  HS65_LH_BFX2 U21494 ( .A(n37238), .Z(n37235) );
  HS65_LH_BFX2 U21495 ( .A(n37239), .Z(n37236) );
  HS65_LH_BFX2 U21496 ( .A(n37234), .Z(n37237) );
  HS65_LH_BFX2 U21497 ( .A(n37241), .Z(n37238) );
  HS65_LH_BFX2 U21498 ( .A(n37242), .Z(n37239) );
  HS65_LH_BFX2 U21499 ( .A(n37237), .Z(n37240) );
  HS65_LH_BFX2 U21500 ( .A(n37244), .Z(n37241) );
  HS65_LH_BFX2 U21501 ( .A(n37245), .Z(n37242) );
  HS65_LH_BFX2 U21502 ( .A(n37240), .Z(n37243) );
  HS65_LH_BFX2 U21503 ( .A(n37247), .Z(n37244) );
  HS65_LH_BFX2 U21504 ( .A(n37248), .Z(n37245) );
  HS65_LH_BFX2 U21505 ( .A(n37243), .Z(n37246) );
  HS65_LH_BFX2 U21506 ( .A(n37252), .Z(n37247) );
  HS65_LH_BFX2 U21507 ( .A(n37253), .Z(n37248) );
  HS65_LH_BFX2 U21508 ( .A(n16600), .Z(n37249) );
  HS65_LH_IVX2 U21509 ( .A(n37246), .Z(n37250) );
  HS65_LH_IVX2 U21510 ( .A(n37250), .Z(n37251) );
  HS65_LH_BFX2 U21511 ( .A(n37254), .Z(n37252) );
  HS65_LH_BFX2 U21512 ( .A(n1749), .Z(n37253) );
  HS65_LH_BFX2 U21513 ( .A(n37255), .Z(n37254) );
  HS65_LH_BFX2 U21514 ( .A(n37256), .Z(n37255) );
  HS65_LH_BFX2 U21515 ( .A(n37257), .Z(n37256) );
  HS65_LH_BFX2 U21516 ( .A(n17931), .Z(n37257) );
  HS65_LH_BFX2 U21517 ( .A(n37263), .Z(n37258) );
  HS65_LH_BFX2 U21518 ( .A(n37265), .Z(n37259) );
  HS65_LH_IVX2 U21519 ( .A(n37267), .Z(n37260) );
  HS65_LH_IVX2 U21520 ( .A(n37260), .Z(n37261) );
  HS65_LH_IVX2 U21521 ( .A(n37269), .Z(n37262) );
  HS65_LH_IVX2 U21522 ( .A(n37262), .Z(n37263) );
  HS65_LH_IVX2 U21523 ( .A(n37271), .Z(n37264) );
  HS65_LH_IVX2 U21524 ( .A(n37264), .Z(n37265) );
  HS65_LH_IVX2 U21525 ( .A(n37273), .Z(n37266) );
  HS65_LH_IVX2 U21526 ( .A(n37266), .Z(n37267) );
  HS65_LH_IVX2 U21527 ( .A(n37275), .Z(n37268) );
  HS65_LH_IVX2 U21528 ( .A(n37268), .Z(n37269) );
  HS65_LH_IVX2 U21529 ( .A(n37277), .Z(n37270) );
  HS65_LH_IVX2 U21530 ( .A(n37270), .Z(n37271) );
  HS65_LH_IVX2 U21531 ( .A(n37279), .Z(n37272) );
  HS65_LH_IVX2 U21532 ( .A(n37272), .Z(n37273) );
  HS65_LH_IVX2 U21533 ( .A(n37281), .Z(n37274) );
  HS65_LH_IVX2 U21534 ( .A(n37274), .Z(n37275) );
  HS65_LH_IVX2 U21535 ( .A(n37283), .Z(n37276) );
  HS65_LH_IVX2 U21536 ( .A(n37276), .Z(n37277) );
  HS65_LH_IVX2 U21537 ( .A(n37285), .Z(n37278) );
  HS65_LH_IVX2 U21538 ( .A(n37278), .Z(n37279) );
  HS65_LH_IVX2 U21539 ( .A(n37287), .Z(n37280) );
  HS65_LH_IVX2 U21540 ( .A(n37280), .Z(n37281) );
  HS65_LH_IVX2 U21541 ( .A(n37289), .Z(n37282) );
  HS65_LH_IVX2 U21542 ( .A(n37282), .Z(n37283) );
  HS65_LH_IVX2 U21543 ( .A(n37291), .Z(n37284) );
  HS65_LH_IVX2 U21544 ( .A(n37284), .Z(n37285) );
  HS65_LH_IVX2 U21545 ( .A(n37293), .Z(n37286) );
  HS65_LH_IVX2 U21546 ( .A(n37286), .Z(n37287) );
  HS65_LH_IVX2 U21547 ( .A(n37295), .Z(n37288) );
  HS65_LH_IVX2 U21548 ( .A(n37288), .Z(n37289) );
  HS65_LH_IVX2 U21549 ( .A(n37297), .Z(n37290) );
  HS65_LH_IVX2 U21550 ( .A(n37290), .Z(n37291) );
  HS65_LH_IVX2 U21551 ( .A(n37299), .Z(n37292) );
  HS65_LH_IVX2 U21552 ( .A(n37292), .Z(n37293) );
  HS65_LH_IVX2 U21553 ( .A(n37301), .Z(n37294) );
  HS65_LH_IVX2 U21554 ( .A(n37294), .Z(n37295) );
  HS65_LH_IVX2 U21555 ( .A(n37303), .Z(n37296) );
  HS65_LH_IVX2 U21556 ( .A(n37296), .Z(n37297) );
  HS65_LH_IVX2 U21557 ( .A(n37305), .Z(n37298) );
  HS65_LH_IVX2 U21558 ( .A(n37298), .Z(n37299) );
  HS65_LH_IVX2 U21559 ( .A(n37307), .Z(n37300) );
  HS65_LH_IVX2 U21560 ( .A(n37300), .Z(n37301) );
  HS65_LH_IVX2 U21561 ( .A(n37312), .Z(n37302) );
  HS65_LH_IVX2 U21562 ( .A(n37302), .Z(n37303) );
  HS65_LH_IVX2 U21563 ( .A(n37309), .Z(n37304) );
  HS65_LH_IVX2 U21564 ( .A(n37304), .Z(n37305) );
  HS65_LH_IVX2 U21565 ( .A(n37311), .Z(n37306) );
  HS65_LH_IVX2 U21566 ( .A(n37306), .Z(n37307) );
  HS65_LH_IVX2 U21567 ( .A(n37314), .Z(n37308) );
  HS65_LH_IVX2 U21568 ( .A(n37308), .Z(n37309) );
  HS65_LH_IVX2 U21569 ( .A(n37316), .Z(n37310) );
  HS65_LH_IVX2 U21570 ( .A(n37310), .Z(n37311) );
  HS65_LH_BFX2 U21571 ( .A(n37317), .Z(n37312) );
  HS65_LH_IVX2 U21572 ( .A(n37319), .Z(n37313) );
  HS65_LH_IVX2 U21573 ( .A(n37313), .Z(n37314) );
  HS65_LH_IVX2 U21574 ( .A(n37321), .Z(n37315) );
  HS65_LH_IVX2 U21575 ( .A(n37315), .Z(n37316) );
  HS65_LH_BFX2 U21576 ( .A(n37322), .Z(n37317) );
  HS65_LH_IVX2 U21577 ( .A(n37326), .Z(n37318) );
  HS65_LH_IVX2 U21578 ( .A(n37318), .Z(n37319) );
  HS65_LH_IVX2 U21579 ( .A(n37324), .Z(n37320) );
  HS65_LH_IVX2 U21580 ( .A(n37320), .Z(n37321) );
  HS65_LH_BFX2 U21581 ( .A(n37325), .Z(n37322) );
  HS65_LH_IVX2 U21582 ( .A(n37328), .Z(n37323) );
  HS65_LH_IVX2 U21583 ( .A(n37323), .Z(n37324) );
  HS65_LH_BFX2 U21584 ( .A(n37329), .Z(n37325) );
  HS65_LH_BFX2 U21585 ( .A(n37330), .Z(n37326) );
  HS65_LH_IVX2 U21586 ( .A(n1496), .Z(n37327) );
  HS65_LH_IVX2 U21587 ( .A(n37327), .Z(n37328) );
  HS65_LH_BFX2 U21588 ( .A(n37331), .Z(n37329) );
  HS65_LH_BFX2 U21589 ( .A(n37332), .Z(n37330) );
  HS65_LH_BFX2 U21590 ( .A(n37333), .Z(n37331) );
  HS65_LH_BFX2 U21591 ( .A(n1495), .Z(n37332) );
  HS65_LH_BFX2 U21592 ( .A(n37334), .Z(n37333) );
  HS65_LH_BFX2 U21593 ( .A(n37335), .Z(n37334) );
  HS65_LH_BFX2 U21594 ( .A(n37336), .Z(n37335) );
  HS65_LH_BFX2 U21595 ( .A(n17890), .Z(n37336) );
  HS65_LH_BFX2 U21596 ( .A(n17927), .Z(n37337) );
  HS65_LH_NAND4ABX3 U21597 ( .A(n17002), .B(n17001), .C(n17000), .D(n16999), 
        .Z(n1288) );
  HS65_LH_BFX2 U21598 ( .A(n37343), .Z(n37338) );
  HS65_LH_IVX2 U21599 ( .A(n37347), .Z(n37339) );
  HS65_LH_IVX2 U21600 ( .A(n37339), .Z(n37340) );
  HS65_LH_BFX2 U21601 ( .A(n37345), .Z(n37341) );
  HS65_LH_IVX2 U21602 ( .A(n37349), .Z(n37342) );
  HS65_LH_IVX2 U21603 ( .A(n37342), .Z(n37343) );
  HS65_LH_IVX2 U21604 ( .A(n37351), .Z(n37344) );
  HS65_LH_IVX2 U21605 ( .A(n37344), .Z(n37345) );
  HS65_LH_IVX2 U21606 ( .A(n37353), .Z(n37346) );
  HS65_LH_IVX2 U21607 ( .A(n37346), .Z(n37347) );
  HS65_LH_IVX2 U21608 ( .A(n37355), .Z(n37348) );
  HS65_LH_IVX2 U21609 ( .A(n37348), .Z(n37349) );
  HS65_LH_IVX2 U21610 ( .A(n37357), .Z(n37350) );
  HS65_LH_IVX2 U21611 ( .A(n37350), .Z(n37351) );
  HS65_LH_IVX2 U21612 ( .A(n37359), .Z(n37352) );
  HS65_LH_IVX2 U21613 ( .A(n37352), .Z(n37353) );
  HS65_LH_IVX2 U21614 ( .A(n37361), .Z(n37354) );
  HS65_LH_IVX2 U21615 ( .A(n37354), .Z(n37355) );
  HS65_LH_IVX2 U21616 ( .A(n37363), .Z(n37356) );
  HS65_LH_IVX2 U21617 ( .A(n37356), .Z(n37357) );
  HS65_LH_IVX2 U21618 ( .A(n37365), .Z(n37358) );
  HS65_LH_IVX2 U21619 ( .A(n37358), .Z(n37359) );
  HS65_LH_IVX2 U21620 ( .A(n37367), .Z(n37360) );
  HS65_LH_IVX2 U21621 ( .A(n37360), .Z(n37361) );
  HS65_LH_IVX2 U21622 ( .A(n37369), .Z(n37362) );
  HS65_LH_IVX2 U21623 ( .A(n37362), .Z(n37363) );
  HS65_LH_IVX2 U21624 ( .A(n37371), .Z(n37364) );
  HS65_LH_IVX2 U21625 ( .A(n37364), .Z(n37365) );
  HS65_LH_IVX2 U21626 ( .A(n37373), .Z(n37366) );
  HS65_LH_IVX2 U21627 ( .A(n37366), .Z(n37367) );
  HS65_LH_IVX2 U21628 ( .A(n37375), .Z(n37368) );
  HS65_LH_IVX2 U21629 ( .A(n37368), .Z(n37369) );
  HS65_LH_IVX2 U21630 ( .A(n37377), .Z(n37370) );
  HS65_LH_IVX2 U21631 ( .A(n37370), .Z(n37371) );
  HS65_LH_IVX2 U21632 ( .A(n37379), .Z(n37372) );
  HS65_LH_IVX2 U21633 ( .A(n37372), .Z(n37373) );
  HS65_LH_IVX2 U21634 ( .A(n37381), .Z(n37374) );
  HS65_LH_IVX2 U21635 ( .A(n37374), .Z(n37375) );
  HS65_LH_IVX2 U21636 ( .A(n37383), .Z(n37376) );
  HS65_LH_IVX2 U21637 ( .A(n37376), .Z(n37377) );
  HS65_LH_IVX2 U21638 ( .A(n37385), .Z(n37378) );
  HS65_LH_IVX2 U21639 ( .A(n37378), .Z(n37379) );
  HS65_LH_IVX2 U21640 ( .A(n37387), .Z(n37380) );
  HS65_LH_IVX2 U21641 ( .A(n37380), .Z(n37381) );
  HS65_LH_IVX2 U21642 ( .A(n37389), .Z(n37382) );
  HS65_LH_IVX2 U21643 ( .A(n37382), .Z(n37383) );
  HS65_LH_IVX2 U21644 ( .A(n37391), .Z(n37384) );
  HS65_LH_IVX2 U21645 ( .A(n37384), .Z(n37385) );
  HS65_LH_IVX2 U21646 ( .A(n37393), .Z(n37386) );
  HS65_LH_IVX2 U21647 ( .A(n37386), .Z(n37387) );
  HS65_LH_IVX2 U21648 ( .A(n37398), .Z(n37388) );
  HS65_LH_IVX2 U21649 ( .A(n37388), .Z(n37389) );
  HS65_LH_IVX2 U21650 ( .A(n37395), .Z(n37390) );
  HS65_LH_IVX2 U21651 ( .A(n37390), .Z(n37391) );
  HS65_LH_IVX2 U21652 ( .A(n37397), .Z(n37392) );
  HS65_LH_IVX2 U21653 ( .A(n37392), .Z(n37393) );
  HS65_LH_IVX2 U21654 ( .A(n37400), .Z(n37394) );
  HS65_LH_IVX2 U21657 ( .A(n37394), .Z(n37395) );
  HS65_LH_IVX2 U21658 ( .A(n37402), .Z(n37396) );
  HS65_LH_IVX2 U21659 ( .A(n37396), .Z(n37397) );
  HS65_LH_BFX2 U21660 ( .A(n37403), .Z(n37398) );
  HS65_LH_IVX2 U21661 ( .A(n37405), .Z(n37399) );
  HS65_LH_IVX2 U21662 ( .A(n37399), .Z(n37400) );
  HS65_LH_IVX2 U21663 ( .A(n37407), .Z(n37401) );
  HS65_LH_IVX2 U21664 ( .A(n37401), .Z(n37402) );
  HS65_LH_BFX2 U21665 ( .A(n37408), .Z(n37403) );
  HS65_LH_IVX2 U21666 ( .A(n37410), .Z(n37404) );
  HS65_LH_IVX2 U21667 ( .A(n37404), .Z(n37405) );
  HS65_LH_IVX2 U21668 ( .A(n37412), .Z(n37406) );
  HS65_LH_IVX2 U21669 ( .A(n37406), .Z(n37407) );
  HS65_LH_BFX2 U21670 ( .A(n37413), .Z(n37408) );
  HS65_LH_IVX2 U21671 ( .A(n37415), .Z(n37409) );
  HS65_LH_IVX2 U21672 ( .A(n37409), .Z(n37410) );
  HS65_LH_IVX2 U21673 ( .A(n1289), .Z(n37411) );
  HS65_LH_IVX2 U21674 ( .A(n37411), .Z(n37412) );
  HS65_LH_BFX2 U21675 ( .A(n37416), .Z(n37413) );
  HS65_LH_IVX2 U21676 ( .A(n1288), .Z(n37414) );
  HS65_LH_IVX2 U21677 ( .A(n37414), .Z(n37415) );
  HS65_LH_BFX2 U21678 ( .A(n37417), .Z(n37416) );
  HS65_LH_BFX2 U21679 ( .A(n37418), .Z(n37417) );
  HS65_LH_BFX2 U21680 ( .A(n37419), .Z(n37418) );
  HS65_LH_BFX2 U21681 ( .A(n37420), .Z(n37419) );
  HS65_LH_BFX2 U21682 ( .A(n37337), .Z(n37420) );
  HS65_LH_BFX2 U21683 ( .A(n37426), .Z(n37421) );
  HS65_LH_BFX2 U21684 ( .A(n37428), .Z(n37422) );
  HS65_LH_IVX2 U21685 ( .A(n37430), .Z(n37423) );
  HS65_LH_IVX2 U21686 ( .A(n37423), .Z(n37424) );
  HS65_LH_IVX2 U21687 ( .A(n37432), .Z(n37425) );
  HS65_LH_IVX2 U21688 ( .A(n37425), .Z(n37426) );
  HS65_LH_IVX2 U21689 ( .A(n37434), .Z(n37427) );
  HS65_LH_IVX2 U21690 ( .A(n37427), .Z(n37428) );
  HS65_LH_IVX2 U21691 ( .A(n37436), .Z(n37429) );
  HS65_LH_IVX2 U21692 ( .A(n37429), .Z(n37430) );
  HS65_LH_IVX2 U21693 ( .A(n37438), .Z(n37431) );
  HS65_LH_IVX2 U21694 ( .A(n37431), .Z(n37432) );
  HS65_LH_IVX2 U21695 ( .A(n37440), .Z(n37433) );
  HS65_LH_IVX2 U21696 ( .A(n37433), .Z(n37434) );
  HS65_LH_IVX2 U21697 ( .A(n37442), .Z(n37435) );
  HS65_LH_IVX2 U21698 ( .A(n37435), .Z(n37436) );
  HS65_LH_IVX2 U21699 ( .A(n37444), .Z(n37437) );
  HS65_LH_IVX2 U21700 ( .A(n37437), .Z(n37438) );
  HS65_LH_IVX2 U21701 ( .A(n37446), .Z(n37439) );
  HS65_LH_IVX2 U21702 ( .A(n37439), .Z(n37440) );
  HS65_LH_IVX2 U21703 ( .A(n37448), .Z(n37441) );
  HS65_LH_IVX2 U21704 ( .A(n37441), .Z(n37442) );
  HS65_LH_IVX2 U21705 ( .A(n37450), .Z(n37443) );
  HS65_LH_IVX2 U21706 ( .A(n37443), .Z(n37444) );
  HS65_LH_IVX2 U21707 ( .A(n37452), .Z(n37445) );
  HS65_LH_IVX2 U21708 ( .A(n37445), .Z(n37446) );
  HS65_LH_IVX2 U21709 ( .A(n37454), .Z(n37447) );
  HS65_LH_IVX2 U21710 ( .A(n37447), .Z(n37448) );
  HS65_LH_IVX2 U21711 ( .A(n37459), .Z(n37449) );
  HS65_LH_IVX2 U21712 ( .A(n37449), .Z(n37450) );
  HS65_LH_IVX2 U21713 ( .A(n37456), .Z(n37451) );
  HS65_LH_IVX2 U21714 ( .A(n37451), .Z(n37452) );
  HS65_LH_IVX2 U21715 ( .A(n37461), .Z(n37453) );
  HS65_LH_IVX2 U21716 ( .A(n37453), .Z(n37454) );
  HS65_LH_IVX2 U21717 ( .A(n37463), .Z(n37455) );
  HS65_LH_IVX2 U21718 ( .A(n37455), .Z(n37456) );
  HS65_LH_BFX2 U21719 ( .A(n1334), .Z(n37457) );
  HS65_LH_IVX2 U21720 ( .A(n37468), .Z(n37458) );
  HS65_LH_IVX2 U21721 ( .A(n37458), .Z(n37459) );
  HS65_LH_IVX2 U21722 ( .A(n37465), .Z(n37460) );
  HS65_LH_IVX2 U21723 ( .A(n37460), .Z(n37461) );
  HS65_LH_IVX2 U21724 ( .A(n37467), .Z(n37462) );
  HS65_LH_IVX2 U21725 ( .A(n37462), .Z(n37463) );
  HS65_LH_IVX2 U21726 ( .A(n37470), .Z(n37464) );
  HS65_LH_IVX2 U21727 ( .A(n37464), .Z(n37465) );
  HS65_LH_IVX2 U21729 ( .A(n37472), .Z(n37466) );
  HS65_LH_IVX2 U21730 ( .A(n37466), .Z(n37467) );
  HS65_LH_BFX2 U21731 ( .A(n37473), .Z(n37468) );
  HS65_LH_IVX2 U21732 ( .A(n37475), .Z(n37469) );
  HS65_LH_IVX2 U21733 ( .A(n37469), .Z(n37470) );
  HS65_LH_IVX2 U21734 ( .A(n37477), .Z(n37471) );
  HS65_LH_IVX2 U21735 ( .A(n37471), .Z(n37472) );
  HS65_LH_BFX2 U21736 ( .A(n37478), .Z(n37473) );
  HS65_LH_IVX2 U21737 ( .A(n37480), .Z(n37474) );
  HS65_LH_IVX2 U21738 ( .A(n37474), .Z(n37475) );
  HS65_LH_IVX2 U21739 ( .A(n37482), .Z(n37476) );
  HS65_LH_IVX2 U21740 ( .A(n37476), .Z(n37477) );
  HS65_LH_BFX2 U21741 ( .A(n37483), .Z(n37478) );
  HS65_LH_IVX2 U21742 ( .A(n37485), .Z(n37479) );
  HS65_LH_IVX2 U21743 ( .A(n37479), .Z(n37480) );
  HS65_LH_IVX2 U21744 ( .A(n37487), .Z(n37481) );
  HS65_LH_IVX2 U21745 ( .A(n37481), .Z(n37482) );
  HS65_LH_BFX2 U21746 ( .A(n37488), .Z(n37483) );
  HS65_LH_IVX2 U21747 ( .A(n37490), .Z(n37484) );
  HS65_LH_IVX2 U21748 ( .A(n37484), .Z(n37485) );
  HS65_LH_IVX2 U21749 ( .A(n37492), .Z(n37486) );
  HS65_LH_IVX2 U21750 ( .A(n37486), .Z(n37487) );
  HS65_LH_BFX2 U21751 ( .A(n37493), .Z(n37488) );
  HS65_LH_IVX2 U21752 ( .A(n37495), .Z(n37489) );
  HS65_LH_IVX2 U21753 ( .A(n37489), .Z(n37490) );
  HS65_LH_IVX2 U21754 ( .A(n1335), .Z(n37491) );
  HS65_LH_IVX2 U21755 ( .A(n37491), .Z(n37492) );
  HS65_LH_BFX2 U21756 ( .A(n37494), .Z(n37493) );
  HS65_LH_BFX2 U21757 ( .A(n37457), .Z(n37494) );
  HS65_LH_BFX2 U21758 ( .A(n37496), .Z(n37495) );
  HS65_LH_BFX2 U21759 ( .A(n37497), .Z(n37496) );
  HS65_LH_BFX2 U21760 ( .A(n37498), .Z(n37497) );
  HS65_LH_BFX2 U21761 ( .A(n17958), .Z(n37498) );
  HS65_LH_BFX2 U21762 ( .A(n17916), .Z(n37499) );
  HS65_LH_NAND4ABX3 U21763 ( .A(n17070), .B(n17069), .C(n17068), .D(n37575), 
        .Z(n1219) );
  HS65_LH_BFX2 U21764 ( .A(n37505), .Z(n37500) );
  HS65_LH_BFX2 U21765 ( .A(n37507), .Z(n37501) );
  HS65_LH_IVX2 U21766 ( .A(n37509), .Z(n37502) );
  HS65_LH_IVX2 U21767 ( .A(n37502), .Z(n37503) );
  HS65_LH_NAND2X7 U21768 ( .A(n17072), .B(n17071), .Z(n17082) );
  HS65_LH_IVX2 U21769 ( .A(n37511), .Z(n37504) );
  HS65_LH_IVX2 U21770 ( .A(n37504), .Z(n37505) );
  HS65_LH_IVX2 U21771 ( .A(n37513), .Z(n37506) );
  HS65_LH_IVX2 U21772 ( .A(n37506), .Z(n37507) );
  HS65_LH_IVX2 U21773 ( .A(n37515), .Z(n37508) );
  HS65_LH_IVX2 U21774 ( .A(n37508), .Z(n37509) );
  HS65_LH_IVX2 U21775 ( .A(n37517), .Z(n37510) );
  HS65_LH_IVX2 U21776 ( .A(n37510), .Z(n37511) );
  HS65_LH_IVX2 U21777 ( .A(n37519), .Z(n37512) );
  HS65_LH_IVX2 U21778 ( .A(n37512), .Z(n37513) );
  HS65_LH_IVX2 U21779 ( .A(n37521), .Z(n37514) );
  HS65_LH_IVX2 U21780 ( .A(n37514), .Z(n37515) );
  HS65_LH_IVX2 U21781 ( .A(n37523), .Z(n37516) );
  HS65_LH_IVX2 U21782 ( .A(n37516), .Z(n37517) );
  HS65_LH_IVX2 U21783 ( .A(n37525), .Z(n37518) );
  HS65_LH_IVX2 U21784 ( .A(n37518), .Z(n37519) );
  HS65_LH_IVX2 U21785 ( .A(n37527), .Z(n37520) );
  HS65_LH_IVX2 U21786 ( .A(n37520), .Z(n37521) );
  HS65_LH_IVX2 U21787 ( .A(n37529), .Z(n37522) );
  HS65_LH_IVX2 U21788 ( .A(n37522), .Z(n37523) );
  HS65_LH_IVX2 U21789 ( .A(n37531), .Z(n37524) );
  HS65_LH_IVX2 U21790 ( .A(n37524), .Z(n37525) );
  HS65_LH_IVX2 U21791 ( .A(n37533), .Z(n37526) );
  HS65_LH_IVX2 U21792 ( .A(n37526), .Z(n37527) );
  HS65_LH_IVX2 U21793 ( .A(n37535), .Z(n37528) );
  HS65_LH_IVX2 U21794 ( .A(n37528), .Z(n37529) );
  HS65_LH_IVX2 U21795 ( .A(n37537), .Z(n37530) );
  HS65_LH_IVX2 U21796 ( .A(n37530), .Z(n37531) );
  HS65_LH_IVX2 U21797 ( .A(n37539), .Z(n37532) );
  HS65_LH_IVX2 U21798 ( .A(n37532), .Z(n37533) );
  HS65_LH_IVX2 U21799 ( .A(n37541), .Z(n37534) );
  HS65_LH_IVX2 U21800 ( .A(n37534), .Z(n37535) );
  HS65_LH_IVX2 U21801 ( .A(n37543), .Z(n37536) );
  HS65_LH_IVX2 U21802 ( .A(n37536), .Z(n37537) );
  HS65_LH_IVX2 U21803 ( .A(n37545), .Z(n37538) );
  HS65_LH_IVX2 U21804 ( .A(n37538), .Z(n37539) );
  HS65_LH_IVX2 U21805 ( .A(n37547), .Z(n37540) );
  HS65_LH_IVX2 U21806 ( .A(n37540), .Z(n37541) );
  HS65_LH_IVX2 U21807 ( .A(n37549), .Z(n37542) );
  HS65_LH_IVX2 U21808 ( .A(n37542), .Z(n37543) );
  HS65_LH_IVX2 U21809 ( .A(n37551), .Z(n37544) );
  HS65_LH_IVX2 U21810 ( .A(n37544), .Z(n37545) );
  HS65_LH_IVX2 U21811 ( .A(n37553), .Z(n37546) );
  HS65_LH_IVX2 U21812 ( .A(n37546), .Z(n37547) );
  HS65_LH_IVX2 U21813 ( .A(n37555), .Z(n37548) );
  HS65_LH_IVX2 U21814 ( .A(n37548), .Z(n37549) );
  HS65_LH_IVX2 U21815 ( .A(n37560), .Z(n37550) );
  HS65_LH_IVX2 U21816 ( .A(n37550), .Z(n37551) );
  HS65_LH_IVX2 U21817 ( .A(n37557), .Z(n37552) );
  HS65_LH_IVX2 U21818 ( .A(n37552), .Z(n37553) );
  HS65_LH_IVX2 U21819 ( .A(n37559), .Z(n37554) );
  HS65_LH_IVX2 U21820 ( .A(n37554), .Z(n37555) );
  HS65_LH_IVX2 U21821 ( .A(n37562), .Z(n37556) );
  HS65_LH_IVX2 U21822 ( .A(n37556), .Z(n37557) );
  HS65_LH_IVX2 U21823 ( .A(n37564), .Z(n37558) );
  HS65_LH_IVX2 U21824 ( .A(n37558), .Z(n37559) );
  HS65_LH_BFX2 U21825 ( .A(n37565), .Z(n37560) );
  HS65_LH_IVX2 U21826 ( .A(n37567), .Z(n37561) );
  HS65_LH_IVX2 U21827 ( .A(n37561), .Z(n37562) );
  HS65_LH_IVX2 U21828 ( .A(n37569), .Z(n37563) );
  HS65_LH_IVX2 U21829 ( .A(n37563), .Z(n37564) );
  HS65_LH_BFX2 U21830 ( .A(n37570), .Z(n37565) );
  HS65_LH_IVX2 U21831 ( .A(n37574), .Z(n37566) );
  HS65_LH_IVX2 U21832 ( .A(n37566), .Z(n37567) );
  HS65_LH_IVX2 U21833 ( .A(n37572), .Z(n37568) );
  HS65_LH_IVX2 U21834 ( .A(n37568), .Z(n37569) );
  HS65_LH_BFX2 U21835 ( .A(n37573), .Z(n37570) );
  HS65_LH_IVX2 U21836 ( .A(n1220), .Z(n37571) );
  HS65_LH_IVX2 U21837 ( .A(n37571), .Z(n37572) );
  HS65_LH_BFX2 U21838 ( .A(n37578), .Z(n37573) );
  HS65_LH_BFX2 U21839 ( .A(n37577), .Z(n37574) );
  HS65_LH_BFX2 U21840 ( .A(n17067), .Z(n37575) );
  HS65_LH_IVX2 U21841 ( .A(n1219), .Z(n37576) );
  HS65_LH_IVX2 U21842 ( .A(n37576), .Z(n37577) );
  HS65_LH_BFX2 U21843 ( .A(n37579), .Z(n37578) );
  HS65_LH_BFX2 U21844 ( .A(n37580), .Z(n37579) );
  HS65_LH_BFX2 U21845 ( .A(n37581), .Z(n37580) );
  HS65_LH_BFX2 U21846 ( .A(n37582), .Z(n37581) );
  HS65_LH_BFX2 U21847 ( .A(n37499), .Z(n37582) );
  HS65_LH_NAND2X2 U21848 ( .A(n16934), .B(n16933), .Z(n16942) );
  HS65_LH_BFX2 U21849 ( .A(n16942), .Z(n37583) );
  HS65_LH_IVX2 U21850 ( .A(n37592), .Z(n37584) );
  HS65_LH_IVX2 U21851 ( .A(n37584), .Z(n37585) );
  HS65_LH_BFX2 U21852 ( .A(n37590), .Z(n37586) );
  HS65_LH_IVX2 U21853 ( .A(n37594), .Z(n37587) );
  HS65_LH_IVX2 U21854 ( .A(n37587), .Z(n37588) );
  HS65_LH_IVX2 U21855 ( .A(n37596), .Z(n37589) );
  HS65_LH_IVX2 U21856 ( .A(n37589), .Z(n37590) );
  HS65_LH_IVX2 U21857 ( .A(n37598), .Z(n37591) );
  HS65_LH_IVX2 U21858 ( .A(n37591), .Z(n37592) );
  HS65_LH_IVX2 U21859 ( .A(n37600), .Z(n37593) );
  HS65_LH_IVX2 U21860 ( .A(n37593), .Z(n37594) );
  HS65_LH_IVX2 U21861 ( .A(n37602), .Z(n37595) );
  HS65_LH_IVX2 U21862 ( .A(n37595), .Z(n37596) );
  HS65_LH_IVX2 U21863 ( .A(n37604), .Z(n37597) );
  HS65_LH_IVX2 U21864 ( .A(n37597), .Z(n37598) );
  HS65_LH_IVX2 U21865 ( .A(n37606), .Z(n37599) );
  HS65_LH_IVX2 U21866 ( .A(n37599), .Z(n37600) );
  HS65_LH_IVX2 U21867 ( .A(n37608), .Z(n37601) );
  HS65_LH_IVX2 U21868 ( .A(n37601), .Z(n37602) );
  HS65_LH_IVX2 U21869 ( .A(n37610), .Z(n37603) );
  HS65_LH_IVX2 U21870 ( .A(n37603), .Z(n37604) );
  HS65_LH_IVX2 U21871 ( .A(n37612), .Z(n37605) );
  HS65_LH_IVX2 U21872 ( .A(n37605), .Z(n37606) );
  HS65_LH_IVX2 U21873 ( .A(n37614), .Z(n37607) );
  HS65_LH_IVX2 U21874 ( .A(n37607), .Z(n37608) );
  HS65_LH_IVX2 U21875 ( .A(n37616), .Z(n37609) );
  HS65_LH_IVX2 U21876 ( .A(n37609), .Z(n37610) );
  HS65_LH_IVX2 U21877 ( .A(n37618), .Z(n37611) );
  HS65_LH_IVX2 U21878 ( .A(n37611), .Z(n37612) );
  HS65_LH_IVX2 U21879 ( .A(n37620), .Z(n37613) );
  HS65_LH_IVX2 U21880 ( .A(n37613), .Z(n37614) );
  HS65_LH_IVX2 U21881 ( .A(n37622), .Z(n37615) );
  HS65_LH_IVX2 U21882 ( .A(n37615), .Z(n37616) );
  HS65_LH_IVX2 U21883 ( .A(n37624), .Z(n37617) );
  HS65_LH_IVX2 U21884 ( .A(n37617), .Z(n37618) );
  HS65_LH_IVX2 U21885 ( .A(n37626), .Z(n37619) );
  HS65_LH_IVX2 U21886 ( .A(n37619), .Z(n37620) );
  HS65_LH_IVX2 U21887 ( .A(n37628), .Z(n37621) );
  HS65_LH_IVX2 U21888 ( .A(n37621), .Z(n37622) );
  HS65_LH_IVX2 U21889 ( .A(n37630), .Z(n37623) );
  HS65_LH_IVX2 U21890 ( .A(n37623), .Z(n37624) );
  HS65_LH_IVX2 U21891 ( .A(n37632), .Z(n37625) );
  HS65_LH_IVX2 U21892 ( .A(n37625), .Z(n37626) );
  HS65_LH_IVX2 U21893 ( .A(n37637), .Z(n37627) );
  HS65_LH_IVX2 U21894 ( .A(n37627), .Z(n37628) );
  HS65_LH_IVX2 U21895 ( .A(n37634), .Z(n37629) );
  HS65_LH_IVX2 U21896 ( .A(n37629), .Z(n37630) );
  HS65_LH_IVX2 U21897 ( .A(n37636), .Z(n37631) );
  HS65_LH_IVX2 U21898 ( .A(n37631), .Z(n37632) );
  HS65_LH_IVX2 U21899 ( .A(n37639), .Z(n37633) );
  HS65_LH_IVX2 U21900 ( .A(n37633), .Z(n37634) );
  HS65_LH_IVX2 U21901 ( .A(n37641), .Z(n37635) );
  HS65_LH_IVX2 U21902 ( .A(n37635), .Z(n37636) );
  HS65_LH_BFX2 U21903 ( .A(n37642), .Z(n37637) );
  HS65_LH_IVX2 U21904 ( .A(n37644), .Z(n37638) );
  HS65_LH_IVX2 U21905 ( .A(n37638), .Z(n37639) );
  HS65_LH_IVX2 U21906 ( .A(n37646), .Z(n37640) );
  HS65_LH_IVX2 U21907 ( .A(n37640), .Z(n37641) );
  HS65_LH_BFX2 U21908 ( .A(n37647), .Z(n37642) );
  HS65_LH_IVX2 U21909 ( .A(n37651), .Z(n37643) );
  HS65_LH_IVX2 U21910 ( .A(n37643), .Z(n37644) );
  HS65_LH_IVX2 U21911 ( .A(n37649), .Z(n37645) );
  HS65_LH_IVX2 U21912 ( .A(n37645), .Z(n37646) );
  HS65_LH_BFX2 U21913 ( .A(n37650), .Z(n37647) );
  HS65_LH_IVX2 U21914 ( .A(n37654), .Z(n37648) );
  HS65_LH_IVX2 U21915 ( .A(n37648), .Z(n37649) );
  HS65_LH_BFX2 U21916 ( .A(n37657), .Z(n37650) );
  HS65_LH_BFX2 U21917 ( .A(n37656), .Z(n37651) );
  HS65_LH_BFX2 U21918 ( .A(n16941), .Z(n37652) );
  HS65_LH_IVX2 U21919 ( .A(n37659), .Z(n37653) );
  HS65_LH_IVX2 U21920 ( .A(n37653), .Z(n37654) );
  HS65_LH_IVX2 U21921 ( .A(n1357), .Z(n37655) );
  HS65_LH_IVX2 U21922 ( .A(n37655), .Z(n37656) );
  HS65_LH_BFX2 U21923 ( .A(n37658), .Z(n37657) );
  HS65_LH_BFX2 U21924 ( .A(n37660), .Z(n37658) );
  HS65_LH_BFX2 U21925 ( .A(n1358), .Z(n37659) );
  HS65_LH_BFX2 U21926 ( .A(n37661), .Z(n37660) );
  HS65_LH_BFX2 U21927 ( .A(n37662), .Z(n37661) );
  HS65_LH_BFX2 U21928 ( .A(n37663), .Z(n37662) );
  HS65_LH_BFX2 U21929 ( .A(n17909), .Z(n37663) );
  HS65_LH_BFX2 U21930 ( .A(n37667), .Z(n37664) );
  HS65_LH_BFX2 U21931 ( .A(n37668), .Z(n37665) );
  HS65_LH_BFX2 U21932 ( .A(n37669), .Z(n37666) );
  HS65_LH_BFX2 U21933 ( .A(n37670), .Z(n37667) );
  HS65_LH_BFX2 U21934 ( .A(n37671), .Z(n37668) );
  HS65_LH_BFX2 U21935 ( .A(n37672), .Z(n37669) );
  HS65_LH_BFX2 U21936 ( .A(n37673), .Z(n37670) );
  HS65_LH_BFX2 U21937 ( .A(n37674), .Z(n37671) );
  HS65_LH_BFX2 U21938 ( .A(n37675), .Z(n37672) );
  HS65_LH_BFX2 U21939 ( .A(n37676), .Z(n37673) );
  HS65_LH_BFX2 U21940 ( .A(n37677), .Z(n37674) );
  HS65_LH_BFX2 U21941 ( .A(n37678), .Z(n37675) );
  HS65_LH_BFX2 U21942 ( .A(n37679), .Z(n37676) );
  HS65_LH_BFX2 U21943 ( .A(n37680), .Z(n37677) );
  HS65_LH_BFX2 U21944 ( .A(n37681), .Z(n37678) );
  HS65_LH_BFX2 U21945 ( .A(n37682), .Z(n37679) );
  HS65_LH_BFX2 U21946 ( .A(n37683), .Z(n37680) );
  HS65_LH_BFX2 U21947 ( .A(n37684), .Z(n37681) );
  HS65_LH_BFX2 U21948 ( .A(n37685), .Z(n37682) );
  HS65_LH_BFX2 U21949 ( .A(n37686), .Z(n37683) );
  HS65_LH_BFX2 U21950 ( .A(n37687), .Z(n37684) );
  HS65_LH_BFX2 U21951 ( .A(n37688), .Z(n37685) );
  HS65_LH_BFX2 U21952 ( .A(n37689), .Z(n37686) );
  HS65_LH_BFX2 U21953 ( .A(n37690), .Z(n37687) );
  HS65_LH_BFX2 U21954 ( .A(n37691), .Z(n37688) );
  HS65_LH_BFX2 U21955 ( .A(n37692), .Z(n37689) );
  HS65_LH_BFX2 U21956 ( .A(n37693), .Z(n37690) );
  HS65_LH_BFX2 U21957 ( .A(n37694), .Z(n37691) );
  HS65_LH_BFX2 U21958 ( .A(n37695), .Z(n37692) );
  HS65_LH_BFX2 U21959 ( .A(n37696), .Z(n37693) );
  HS65_LH_BFX2 U21960 ( .A(n37697), .Z(n37694) );
  HS65_LH_BFX2 U21961 ( .A(n37698), .Z(n37695) );
  HS65_LH_BFX2 U21962 ( .A(n37699), .Z(n37696) );
  HS65_LH_BFX2 U21963 ( .A(n37700), .Z(n37697) );
  HS65_LH_BFX2 U21964 ( .A(n37701), .Z(n37698) );
  HS65_LH_BFX2 U21965 ( .A(n37702), .Z(n37699) );
  HS65_LH_BFX2 U21966 ( .A(n37703), .Z(n37700) );
  HS65_LH_BFX2 U21967 ( .A(n37704), .Z(n37701) );
  HS65_LH_BFX2 U21968 ( .A(n37705), .Z(n37702) );
  HS65_LH_BFX2 U21969 ( .A(n37706), .Z(n37703) );
  HS65_LH_BFX2 U21970 ( .A(n37707), .Z(n37704) );
  HS65_LH_BFX2 U21971 ( .A(n37708), .Z(n37705) );
  HS65_LH_BFX2 U21972 ( .A(n37709), .Z(n37706) );
  HS65_LH_BFX2 U21973 ( .A(n37710), .Z(n37707) );
  HS65_LH_BFX2 U21974 ( .A(n37711), .Z(n37708) );
  HS65_LH_BFX2 U21975 ( .A(n1380), .Z(n37709) );
  HS65_LH_BFX2 U21976 ( .A(n1381), .Z(n37710) );
  HS65_LH_BFX2 U21977 ( .A(n37712), .Z(n37711) );
  HS65_LH_BFX2 U21978 ( .A(n37713), .Z(n37712) );
  HS65_LH_BFX2 U21979 ( .A(n37714), .Z(n37713) );
  HS65_LH_BFX2 U21980 ( .A(n17935), .Z(n37714) );
  HS65_LH_BFX2 U21981 ( .A(n37720), .Z(n37715) );
  HS65_LH_IVX2 U21982 ( .A(n37724), .Z(n37716) );
  HS65_LH_IVX2 U21983 ( .A(n37716), .Z(n37717) );
  HS65_LH_NAND4ABX3 U21984 ( .A(n16992), .B(n16991), .C(n16990), .D(n16989), 
        .Z(n1312) );
  HS65_LH_BFX2 U21985 ( .A(n37722), .Z(n37718) );
  HS65_LH_NAND4ABX3 U21986 ( .A(n16982), .B(n16981), .C(n16980), .D(n16979), 
        .Z(n1311) );
  HS65_LH_IVX2 U21987 ( .A(n37726), .Z(n37719) );
  HS65_LH_IVX2 U21988 ( .A(n37719), .Z(n37720) );
  HS65_LH_IVX2 U21989 ( .A(n37728), .Z(n37721) );
  HS65_LH_IVX2 U21990 ( .A(n37721), .Z(n37722) );
  HS65_LH_IVX2 U21991 ( .A(n37730), .Z(n37723) );
  HS65_LH_IVX2 U21992 ( .A(n37723), .Z(n37724) );
  HS65_LH_IVX2 U21993 ( .A(n37732), .Z(n37725) );
  HS65_LH_IVX2 U21994 ( .A(n37725), .Z(n37726) );
  HS65_LH_IVX2 U21995 ( .A(n37734), .Z(n37727) );
  HS65_LH_IVX2 U21996 ( .A(n37727), .Z(n37728) );
  HS65_LH_IVX2 U21997 ( .A(n37736), .Z(n37729) );
  HS65_LH_IVX2 U21998 ( .A(n37729), .Z(n37730) );
  HS65_LH_IVX2 U21999 ( .A(n37738), .Z(n37731) );
  HS65_LH_IVX2 U22000 ( .A(n37731), .Z(n37732) );
  HS65_LH_IVX2 U22001 ( .A(n37740), .Z(n37733) );
  HS65_LH_IVX2 U22002 ( .A(n37733), .Z(n37734) );
  HS65_LH_IVX2 U22003 ( .A(n37742), .Z(n37735) );
  HS65_LH_IVX2 U22004 ( .A(n37735), .Z(n37736) );
  HS65_LH_IVX2 U22005 ( .A(n37744), .Z(n37737) );
  HS65_LH_IVX2 U22006 ( .A(n37737), .Z(n37738) );
  HS65_LH_IVX2 U22007 ( .A(n37746), .Z(n37739) );
  HS65_LH_IVX2 U22008 ( .A(n37739), .Z(n37740) );
  HS65_LH_IVX2 U22009 ( .A(n37748), .Z(n37741) );
  HS65_LH_IVX2 U22010 ( .A(n37741), .Z(n37742) );
  HS65_LH_IVX2 U22011 ( .A(n37750), .Z(n37743) );
  HS65_LH_IVX2 U22012 ( .A(n37743), .Z(n37744) );
  HS65_LH_IVX2 U22013 ( .A(n37752), .Z(n37745) );
  HS65_LH_IVX2 U22014 ( .A(n37745), .Z(n37746) );
  HS65_LH_IVX2 U22015 ( .A(n37754), .Z(n37747) );
  HS65_LH_IVX2 U22016 ( .A(n37747), .Z(n37748) );
  HS65_LH_IVX2 U22017 ( .A(n37756), .Z(n37749) );
  HS65_LH_IVX2 U22018 ( .A(n37749), .Z(n37750) );
  HS65_LH_IVX2 U22019 ( .A(n37758), .Z(n37751) );
  HS65_LH_IVX2 U22020 ( .A(n37751), .Z(n37752) );
  HS65_LH_IVX2 U22021 ( .A(n37760), .Z(n37753) );
  HS65_LH_IVX2 U22022 ( .A(n37753), .Z(n37754) );
  HS65_LH_IVX2 U22023 ( .A(n37762), .Z(n37755) );
  HS65_LH_IVX2 U22024 ( .A(n37755), .Z(n37756) );
  HS65_LH_IVX2 U22025 ( .A(n37764), .Z(n37757) );
  HS65_LH_IVX2 U22026 ( .A(n37757), .Z(n37758) );
  HS65_LH_IVX2 U22027 ( .A(n37766), .Z(n37759) );
  HS65_LH_IVX2 U22028 ( .A(n37759), .Z(n37760) );
  HS65_LH_IVX2 U22029 ( .A(n37768), .Z(n37761) );
  HS65_LH_IVX2 U22030 ( .A(n37761), .Z(n37762) );
  HS65_LH_IVX2 U22031 ( .A(n37770), .Z(n37763) );
  HS65_LH_IVX2 U22032 ( .A(n37763), .Z(n37764) );
  HS65_LH_IVX2 U22033 ( .A(n37772), .Z(n37765) );
  HS65_LH_IVX2 U22034 ( .A(n37765), .Z(n37766) );
  HS65_LH_IVX2 U22035 ( .A(n37774), .Z(n37767) );
  HS65_LH_IVX2 U22036 ( .A(n37767), .Z(n37768) );
  HS65_LH_IVX2 U22037 ( .A(n37776), .Z(n37769) );
  HS65_LH_IVX2 U22038 ( .A(n37769), .Z(n37770) );
  HS65_LH_IVX2 U22039 ( .A(n37778), .Z(n37771) );
  HS65_LH_IVX2 U22040 ( .A(n37771), .Z(n37772) );
  HS65_LH_IVX2 U22041 ( .A(n37780), .Z(n37773) );
  HS65_LH_IVX2 U22042 ( .A(n37773), .Z(n37774) );
  HS65_LH_IVX2 U22043 ( .A(n37782), .Z(n37775) );
  HS65_LH_IVX2 U22044 ( .A(n37775), .Z(n37776) );
  HS65_LH_IVX2 U22045 ( .A(n37787), .Z(n37777) );
  HS65_LH_IVX2 U22048 ( .A(n37777), .Z(n37778) );
  HS65_LH_IVX2 U22049 ( .A(n37784), .Z(n37779) );
  HS65_LH_IVX2 U22050 ( .A(n37779), .Z(n37780) );
  HS65_LH_IVX2 U22051 ( .A(n37786), .Z(n37781) );
  HS65_LH_IVX2 U22052 ( .A(n37781), .Z(n37782) );
  HS65_LH_IVX2 U22053 ( .A(n37789), .Z(n37783) );
  HS65_LH_IVX2 U22054 ( .A(n37783), .Z(n37784) );
  HS65_LH_IVX2 U22055 ( .A(n37791), .Z(n37785) );
  HS65_LH_IVX2 U22056 ( .A(n37785), .Z(n37786) );
  HS65_LH_BFX2 U22057 ( .A(n37792), .Z(n37787) );
  HS65_LH_IVX2 U22058 ( .A(n37794), .Z(n37788) );
  HS65_LH_IVX2 U22059 ( .A(n37788), .Z(n37789) );
  HS65_LH_IVX2 U22060 ( .A(n37796), .Z(n37790) );
  HS65_LH_IVX2 U22061 ( .A(n37790), .Z(n37791) );
  HS65_LH_BFX2 U22062 ( .A(n37797), .Z(n37792) );
  HS65_LH_IVX2 U22065 ( .A(n1311), .Z(n37793) );
  HS65_LH_IVX2 U22066 ( .A(n37793), .Z(n37794) );
  HS65_LH_IVX2 U22067 ( .A(n1312), .Z(n37795) );
  HS65_LH_IVX2 U22068 ( .A(n37795), .Z(n37796) );
  HS65_LH_BFX2 U22069 ( .A(n37798), .Z(n37797) );
  HS65_LH_BFX2 U22070 ( .A(n37799), .Z(n37798) );
  HS65_LH_BFX2 U22071 ( .A(n37800), .Z(n37799) );
  HS65_LH_BFX2 U22072 ( .A(n37801), .Z(n37800) );
  HS65_LH_BFX2 U22073 ( .A(n17920), .Z(n37801) );
  HS65_LH_BFX2 U22074 ( .A(n37805), .Z(n37802) );
  HS65_LH_BFX2 U22075 ( .A(n37806), .Z(n37803) );
  HS65_LH_BFX2 U22076 ( .A(n37807), .Z(n37804) );
  HS65_LH_BFX2 U22077 ( .A(n37808), .Z(n37805) );
  HS65_LH_BFX2 U22078 ( .A(n37809), .Z(n37806) );
  HS65_LH_BFX2 U22079 ( .A(n37810), .Z(n37807) );
  HS65_LH_BFX2 U22080 ( .A(n37811), .Z(n37808) );
  HS65_LH_BFX2 U22081 ( .A(n37812), .Z(n37809) );
  HS65_LH_BFX2 U22082 ( .A(n37813), .Z(n37810) );
  HS65_LH_BFX2 U22083 ( .A(n37814), .Z(n37811) );
  HS65_LH_BFX2 U22084 ( .A(n37815), .Z(n37812) );
  HS65_LH_BFX2 U22085 ( .A(n37816), .Z(n37813) );
  HS65_LH_BFX2 U22086 ( .A(n37817), .Z(n37814) );
  HS65_LH_BFX2 U22087 ( .A(n37818), .Z(n37815) );
  HS65_LH_BFX2 U22088 ( .A(n37819), .Z(n37816) );
  HS65_LH_BFX2 U22089 ( .A(n37820), .Z(n37817) );
  HS65_LH_BFX2 U22090 ( .A(n37821), .Z(n37818) );
  HS65_LH_BFX2 U22091 ( .A(n37822), .Z(n37819) );
  HS65_LH_BFX2 U22092 ( .A(n37823), .Z(n37820) );
  HS65_LH_BFX2 U22093 ( .A(n37824), .Z(n37821) );
  HS65_LH_BFX2 U22094 ( .A(n37825), .Z(n37822) );
  HS65_LH_BFX2 U22095 ( .A(n37826), .Z(n37823) );
  HS65_LH_BFX2 U22096 ( .A(n37827), .Z(n37824) );
  HS65_LH_BFX2 U22097 ( .A(n37828), .Z(n37825) );
  HS65_LH_BFX2 U22098 ( .A(n37829), .Z(n37826) );
  HS65_LH_BFX2 U22099 ( .A(n37830), .Z(n37827) );
  HS65_LH_BFX2 U22100 ( .A(n37831), .Z(n37828) );
  HS65_LH_BFX2 U22101 ( .A(n37832), .Z(n37829) );
  HS65_LH_BFX2 U22102 ( .A(n37833), .Z(n37830) );
  HS65_LH_BFX2 U22103 ( .A(n37834), .Z(n37831) );
  HS65_LH_BFX2 U22104 ( .A(n37835), .Z(n37832) );
  HS65_LH_BFX2 U22105 ( .A(n37836), .Z(n37833) );
  HS65_LH_BFX2 U22106 ( .A(n37837), .Z(n37834) );
  HS65_LH_BFX2 U22107 ( .A(n37838), .Z(n37835) );
  HS65_LH_BFX2 U22108 ( .A(n37839), .Z(n37836) );
  HS65_LH_BFX2 U22109 ( .A(n37840), .Z(n37837) );
  HS65_LH_BFX2 U22110 ( .A(n37841), .Z(n37838) );
  HS65_LH_BFX2 U22111 ( .A(n37842), .Z(n37839) );
  HS65_LH_BFX2 U22112 ( .A(n37843), .Z(n37840) );
  HS65_LH_BFX2 U22113 ( .A(n37844), .Z(n37841) );
  HS65_LH_BFX2 U22114 ( .A(n37845), .Z(n37842) );
  HS65_LH_BFX2 U22115 ( .A(n37846), .Z(n37843) );
  HS65_LH_BFX2 U22116 ( .A(n37847), .Z(n37844) );
  HS65_LH_BFX2 U22117 ( .A(n37848), .Z(n37845) );
  HS65_LH_BFX2 U22118 ( .A(n37849), .Z(n37846) );
  HS65_LH_BFX2 U22119 ( .A(n1426), .Z(n37847) );
  HS65_LH_BFX2 U22120 ( .A(n1427), .Z(n37848) );
  HS65_LH_BFX2 U22121 ( .A(n37850), .Z(n37849) );
  HS65_LH_BFX2 U22122 ( .A(n37851), .Z(n37850) );
  HS65_LH_BFX2 U22123 ( .A(n37852), .Z(n37851) );
  HS65_LH_BFX2 U22124 ( .A(n17978), .Z(n37852) );
  HS65_LH_BFX2 U22125 ( .A(n37908), .Z(n37853) );
  HS65_LH_BFX2 U22126 ( .A(n37857), .Z(n37854) );
  HS65_LH_BFX2 U22127 ( .A(n37859), .Z(n37855) );
  HS65_LH_IVX2 U22128 ( .A(n37862), .Z(n37856) );
  HS65_LH_IVX2 U22129 ( .A(n37856), .Z(n37857) );
  HS65_LH_IVX2 U22130 ( .A(n37864), .Z(n37858) );
  HS65_LH_IVX2 U22131 ( .A(n37858), .Z(n37859) );
  HS65_LH_BFX2 U22132 ( .A(n1242), .Z(n37860) );
  HS65_LH_IVX2 U22133 ( .A(n37867), .Z(n37861) );
  HS65_LH_IVX2 U22134 ( .A(n37861), .Z(n37862) );
  HS65_LH_IVX2 U22135 ( .A(n37869), .Z(n37863) );
  HS65_LH_IVX2 U22136 ( .A(n37863), .Z(n37864) );
  HS65_LH_BFX2 U22137 ( .A(n37860), .Z(n37865) );
  HS65_LH_IVX2 U22138 ( .A(n37872), .Z(n37866) );
  HS65_LH_IVX2 U22139 ( .A(n37866), .Z(n37867) );
  HS65_LH_IVX2 U22140 ( .A(n37874), .Z(n37868) );
  HS65_LH_IVX2 U22141 ( .A(n37868), .Z(n37869) );
  HS65_LH_BFX2 U22142 ( .A(n37865), .Z(n37870) );
  HS65_LH_IVX2 U22143 ( .A(n37877), .Z(n37871) );
  HS65_LH_IVX2 U22144 ( .A(n37871), .Z(n37872) );
  HS65_LH_IVX2 U22145 ( .A(n37879), .Z(n37873) );
  HS65_LH_IVX2 U22146 ( .A(n37873), .Z(n37874) );
  HS65_LH_BFX2 U22147 ( .A(n37870), .Z(n37875) );
  HS65_LH_IVX2 U22148 ( .A(n37882), .Z(n37876) );
  HS65_LH_IVX2 U22149 ( .A(n37876), .Z(n37877) );
  HS65_LH_IVX2 U22150 ( .A(n37884), .Z(n37878) );
  HS65_LH_IVX2 U22151 ( .A(n37878), .Z(n37879) );
  HS65_LH_BFX2 U22152 ( .A(n37875), .Z(n37880) );
  HS65_LH_IVX2 U22153 ( .A(n37887), .Z(n37881) );
  HS65_LH_IVX2 U22154 ( .A(n37881), .Z(n37882) );
  HS65_LH_IVX2 U22155 ( .A(n37889), .Z(n37883) );
  HS65_LH_IVX2 U22156 ( .A(n37883), .Z(n37884) );
  HS65_LH_BFX2 U22157 ( .A(n37880), .Z(n37885) );
  HS65_LH_IVX2 U22158 ( .A(n37892), .Z(n37886) );
  HS65_LH_IVX2 U22159 ( .A(n37886), .Z(n37887) );
  HS65_LH_IVX2 U22160 ( .A(n37894), .Z(n37888) );
  HS65_LH_IVX2 U22161 ( .A(n37888), .Z(n37889) );
  HS65_LH_BFX2 U22162 ( .A(n37885), .Z(n37890) );
  HS65_LH_IVX2 U22163 ( .A(n37897), .Z(n37891) );
  HS65_LH_IVX2 U22164 ( .A(n37891), .Z(n37892) );
  HS65_LH_IVX2 U22165 ( .A(n37899), .Z(n37893) );
  HS65_LH_IVX2 U22166 ( .A(n37893), .Z(n37894) );
  HS65_LH_BFX2 U22167 ( .A(n37890), .Z(n37895) );
  HS65_LH_IVX2 U22168 ( .A(n37903), .Z(n37896) );
  HS65_LH_IVX2 U22169 ( .A(n37896), .Z(n37897) );
  HS65_LH_IVX2 U22170 ( .A(n37905), .Z(n37898) );
  HS65_LH_IVX2 U22171 ( .A(n37898), .Z(n37899) );
  HS65_LH_BFX2 U22172 ( .A(n37895), .Z(n37900) );
  HS65_LH_BFX2 U22173 ( .A(n37900), .Z(n37901) );
  HS65_LH_IVX2 U22174 ( .A(n37910), .Z(n37902) );
  HS65_LH_IVX2 U22175 ( .A(n37902), .Z(n37903) );
  HS65_LH_IVX2 U22176 ( .A(n37912), .Z(n37904) );
  HS65_LH_IVX2 U22177 ( .A(n37904), .Z(n37905) );
  HS65_LH_BFX2 U22178 ( .A(n37901), .Z(n37906) );
  HS65_LH_IVX2 U22179 ( .A(n37917), .Z(n37907) );
  HS65_LH_IVX2 U22180 ( .A(n37907), .Z(n37908) );
  HS65_LH_IVX2 U22181 ( .A(n37914), .Z(n37909) );
  HS65_LH_IVX2 U22182 ( .A(n37909), .Z(n37910) );
  HS65_LH_IVX2 U22183 ( .A(n37916), .Z(n37911) );
  HS65_LH_IVX2 U22184 ( .A(n37911), .Z(n37912) );
  HS65_LH_IVX2 U22185 ( .A(n37919), .Z(n37913) );
  HS65_LH_IVX2 U22186 ( .A(n37913), .Z(n37914) );
  HS65_LH_IVX2 U22187 ( .A(n37921), .Z(n37915) );
  HS65_LH_IVX2 U22188 ( .A(n37915), .Z(n37916) );
  HS65_LH_BFX2 U22189 ( .A(n37925), .Z(n37917) );
  HS65_LH_IVX2 U22190 ( .A(n37924), .Z(n37918) );
  HS65_LH_IVX2 U22191 ( .A(n37918), .Z(n37919) );
  HS65_LH_IVX2 U22192 ( .A(n1243), .Z(n37920) );
  HS65_LH_IVX2 U22193 ( .A(n37920), .Z(n37921) );
  HS65_LH_BFX2 U22194 ( .A(n29534), .Z(n37922) );
  HS65_LH_IVX2 U22195 ( .A(n37926), .Z(n37923) );
  HS65_LH_IVX2 U22196 ( .A(n37923), .Z(n37924) );
  HS65_LH_BFX2 U22197 ( .A(n37906), .Z(n37925) );
  HS65_LH_BFX2 U22198 ( .A(n37927), .Z(n37926) );
  HS65_LH_BFX2 U22199 ( .A(n37928), .Z(n37927) );
  HS65_LH_BFX2 U22200 ( .A(n17996), .Z(n37928) );
  HS65_LH_IVX2 U22201 ( .A(n16521), .Z(n37929) );
  HS65_LH_IVX2 U22202 ( .A(n37929), .Z(n37930) );
  HS65_LH_NAND2X2 U22203 ( .A(n16514), .B(n16513), .Z(n16522) );
  HS65_LH_BFX2 U22204 ( .A(n16522), .Z(n37931) );
  HS65_LH_BFX2 U22205 ( .A(n37935), .Z(n37932) );
  HS65_LH_BFX2 U22206 ( .A(n37939), .Z(n37933) );
  HS65_LH_IVX2 U22207 ( .A(n37941), .Z(n37934) );
  HS65_LH_IVX2 U22208 ( .A(n37934), .Z(n37935) );
  HS65_LH_IVX2 U22209 ( .A(n37943), .Z(n37936) );
  HS65_LH_IVX2 U22210 ( .A(n37936), .Z(n37937) );
  HS65_LH_IVX2 U22211 ( .A(n37945), .Z(n37938) );
  HS65_LH_IVX2 U22212 ( .A(n37938), .Z(n37939) );
  HS65_LH_IVX2 U22213 ( .A(n37947), .Z(n37940) );
  HS65_LH_IVX2 U22214 ( .A(n37940), .Z(n37941) );
  HS65_LH_IVX2 U22215 ( .A(n37949), .Z(n37942) );
  HS65_LH_IVX2 U22216 ( .A(n37942), .Z(n37943) );
  HS65_LH_IVX2 U22217 ( .A(n37951), .Z(n37944) );
  HS65_LH_IVX2 U22218 ( .A(n37944), .Z(n37945) );
  HS65_LH_IVX2 U22219 ( .A(n37953), .Z(n37946) );
  HS65_LH_IVX2 U22220 ( .A(n37946), .Z(n37947) );
  HS65_LH_IVX2 U22221 ( .A(n37955), .Z(n37948) );
  HS65_LH_IVX2 U22222 ( .A(n37948), .Z(n37949) );
  HS65_LH_IVX2 U22223 ( .A(n37957), .Z(n37950) );
  HS65_LH_IVX2 U22224 ( .A(n37950), .Z(n37951) );
  HS65_LH_IVX2 U22225 ( .A(n37959), .Z(n37952) );
  HS65_LH_IVX2 U22226 ( .A(n37952), .Z(n37953) );
  HS65_LH_IVX2 U22227 ( .A(n37961), .Z(n37954) );
  HS65_LH_IVX2 U22228 ( .A(n37954), .Z(n37955) );
  HS65_LH_IVX2 U22229 ( .A(n37963), .Z(n37956) );
  HS65_LH_IVX2 U22230 ( .A(n37956), .Z(n37957) );
  HS65_LH_IVX2 U22231 ( .A(n37965), .Z(n37958) );
  HS65_LH_IVX2 U22232 ( .A(n37958), .Z(n37959) );
  HS65_LH_IVX2 U22233 ( .A(n37967), .Z(n37960) );
  HS65_LH_IVX2 U22234 ( .A(n37960), .Z(n37961) );
  HS65_LH_IVX2 U22235 ( .A(n37969), .Z(n37962) );
  HS65_LH_IVX2 U22236 ( .A(n37962), .Z(n37963) );
  HS65_LH_IVX2 U22237 ( .A(n37971), .Z(n37964) );
  HS65_LH_IVX2 U22238 ( .A(n37964), .Z(n37965) );
  HS65_LH_IVX2 U22239 ( .A(n37973), .Z(n37966) );
  HS65_LH_IVX2 U22240 ( .A(n37966), .Z(n37967) );
  HS65_LH_IVX2 U22241 ( .A(n37975), .Z(n37968) );
  HS65_LH_IVX2 U22242 ( .A(n37968), .Z(n37969) );
  HS65_LH_IVX2 U22243 ( .A(n37977), .Z(n37970) );
  HS65_LH_IVX2 U22244 ( .A(n37970), .Z(n37971) );
  HS65_LH_IVX2 U22245 ( .A(n37979), .Z(n37972) );
  HS65_LH_IVX2 U22246 ( .A(n37972), .Z(n37973) );
  HS65_LH_IVX2 U22247 ( .A(n37981), .Z(n37974) );
  HS65_LH_IVX2 U22248 ( .A(n37974), .Z(n37975) );
  HS65_LH_IVX2 U22249 ( .A(n37983), .Z(n37976) );
  HS65_LH_IVX2 U22250 ( .A(n37976), .Z(n37977) );
  HS65_LH_IVX2 U22251 ( .A(n37985), .Z(n37978) );
  HS65_LH_IVX2 U22252 ( .A(n37978), .Z(n37979) );
  HS65_LH_IVX2 U22253 ( .A(n37987), .Z(n37980) );
  HS65_LH_IVX2 U22254 ( .A(n37980), .Z(n37981) );
  HS65_LH_IVX2 U22255 ( .A(n37989), .Z(n37982) );
  HS65_LH_IVX2 U22256 ( .A(n37982), .Z(n37983) );
  HS65_LH_IVX2 U22257 ( .A(n37991), .Z(n37984) );
  HS65_LH_IVX2 U22258 ( .A(n37984), .Z(n37985) );
  HS65_LH_IVX2 U22259 ( .A(n37993), .Z(n37986) );
  HS65_LH_IVX2 U22260 ( .A(n37986), .Z(n37987) );
  HS65_LH_IVX2 U22261 ( .A(n37998), .Z(n37988) );
  HS65_LH_IVX2 U22262 ( .A(n37988), .Z(n37989) );
  HS65_LH_IVX2 U22263 ( .A(n37995), .Z(n37990) );
  HS65_LH_IVX2 U22264 ( .A(n37990), .Z(n37991) );
  HS65_LH_IVX2 U22265 ( .A(n37997), .Z(n37992) );
  HS65_LH_IVX2 U22266 ( .A(n37992), .Z(n37993) );
  HS65_LH_IVX2 U22267 ( .A(n38000), .Z(n37994) );
  HS65_LH_IVX2 U22268 ( .A(n37994), .Z(n37995) );
  HS65_LH_IVX2 U22269 ( .A(n38002), .Z(n37996) );
  HS65_LH_IVX2 U22270 ( .A(n37996), .Z(n37997) );
  HS65_LH_BFX2 U22271 ( .A(n38003), .Z(n37998) );
  HS65_LH_IVX2 U22272 ( .A(n38007), .Z(n37999) );
  HS65_LH_IVX2 U22273 ( .A(n37999), .Z(n38000) );
  HS65_LH_IVX2 U22274 ( .A(n38005), .Z(n38001) );
  HS65_LH_IVX2 U22275 ( .A(n38001), .Z(n38002) );
  HS65_LH_BFX2 U22276 ( .A(n38008), .Z(n38003) );
  HS65_LH_IVX2 U22277 ( .A(n38010), .Z(n38004) );
  HS65_LH_IVX2 U22278 ( .A(n38004), .Z(n38005) );
  HS65_LH_IVX2 U22279 ( .A(n1840), .Z(n38006) );
  HS65_LH_IVX2 U22280 ( .A(n38006), .Z(n38007) );
  HS65_LH_BFX2 U22281 ( .A(n38009), .Z(n38008) );
  HS65_LH_BFX2 U22282 ( .A(n38011), .Z(n38009) );
  HS65_LH_BFX2 U22283 ( .A(n1841), .Z(n38010) );
  HS65_LH_BFX2 U22284 ( .A(n38012), .Z(n38011) );
  HS65_LH_BFX2 U22285 ( .A(n38013), .Z(n38012) );
  HS65_LH_BFX2 U22286 ( .A(n38014), .Z(n38013) );
  HS65_LH_BFX2 U22287 ( .A(n17865), .Z(n38014) );
  HS65_LH_BFX2 U22288 ( .A(n38021), .Z(n38015) );
  HS65_LH_BFX2 U22289 ( .A(n38019), .Z(n38016) );
  HS65_LH_BFX2 U22290 ( .A(n38023), .Z(n38017) );
  HS65_LH_IVX2 U22291 ( .A(n38025), .Z(n38018) );
  HS65_LH_IVX2 U22292 ( .A(n38018), .Z(n38019) );
  HS65_LH_IVX2 U22293 ( .A(n38027), .Z(n38020) );
  HS65_LH_IVX2 U22294 ( .A(n38020), .Z(n38021) );
  HS65_LH_IVX2 U22295 ( .A(n38029), .Z(n38022) );
  HS65_LH_IVX2 U22296 ( .A(n38022), .Z(n38023) );
  HS65_LH_IVX2 U22297 ( .A(n38031), .Z(n38024) );
  HS65_LH_IVX2 U22298 ( .A(n38024), .Z(n38025) );
  HS65_LH_IVX2 U22299 ( .A(n38033), .Z(n38026) );
  HS65_LH_IVX2 U22300 ( .A(n38026), .Z(n38027) );
  HS65_LH_IVX2 U22301 ( .A(n38035), .Z(n38028) );
  HS65_LH_IVX2 U22302 ( .A(n38028), .Z(n38029) );
  HS65_LH_IVX2 U22303 ( .A(n38037), .Z(n38030) );
  HS65_LH_IVX2 U22304 ( .A(n38030), .Z(n38031) );
  HS65_LH_IVX2 U22305 ( .A(n38039), .Z(n38032) );
  HS65_LH_IVX2 U22306 ( .A(n38032), .Z(n38033) );
  HS65_LH_IVX2 U22307 ( .A(n38041), .Z(n38034) );
  HS65_LH_IVX2 U22308 ( .A(n38034), .Z(n38035) );
  HS65_LH_IVX2 U22309 ( .A(n38043), .Z(n38036) );
  HS65_LH_IVX2 U22310 ( .A(n38036), .Z(n38037) );
  HS65_LH_IVX2 U22311 ( .A(n38045), .Z(n38038) );
  HS65_LH_IVX2 U22312 ( .A(n38038), .Z(n38039) );
  HS65_LH_IVX2 U22313 ( .A(n38047), .Z(n38040) );
  HS65_LH_IVX2 U22314 ( .A(n38040), .Z(n38041) );
  HS65_LH_IVX2 U22315 ( .A(n38049), .Z(n38042) );
  HS65_LH_IVX2 U22316 ( .A(n38042), .Z(n38043) );
  HS65_LH_IVX2 U22317 ( .A(n38051), .Z(n38044) );
  HS65_LH_IVX2 U22318 ( .A(n38044), .Z(n38045) );
  HS65_LH_IVX2 U22319 ( .A(n38053), .Z(n38046) );
  HS65_LH_IVX2 U22320 ( .A(n38046), .Z(n38047) );
  HS65_LH_IVX2 U22321 ( .A(n38055), .Z(n38048) );
  HS65_LH_IVX2 U22322 ( .A(n38048), .Z(n38049) );
  HS65_LH_IVX2 U22323 ( .A(n38057), .Z(n38050) );
  HS65_LH_IVX2 U22324 ( .A(n38050), .Z(n38051) );
  HS65_LH_IVX2 U22325 ( .A(n38059), .Z(n38052) );
  HS65_LH_IVX2 U22326 ( .A(n38052), .Z(n38053) );
  HS65_LH_IVX2 U22327 ( .A(n38064), .Z(n38054) );
  HS65_LH_IVX2 U22328 ( .A(n38054), .Z(n38055) );
  HS65_LH_IVX2 U22329 ( .A(n38061), .Z(n38056) );
  HS65_LH_IVX2 U22330 ( .A(n38056), .Z(n38057) );
  HS65_LH_IVX2 U22331 ( .A(n38063), .Z(n38058) );
  HS65_LH_IVX2 U22332 ( .A(n38058), .Z(n38059) );
  HS65_LH_IVX2 U22333 ( .A(n38066), .Z(n38060) );
  HS65_LH_IVX2 U22334 ( .A(n38060), .Z(n38061) );
  HS65_LH_IVX2 U22335 ( .A(n38068), .Z(n38062) );
  HS65_LH_IVX2 U22336 ( .A(n38062), .Z(n38063) );
  HS65_LH_BFX2 U22337 ( .A(n38069), .Z(n38064) );
  HS65_LH_IVX2 U22338 ( .A(n38071), .Z(n38065) );
  HS65_LH_IVX2 U22339 ( .A(n38065), .Z(n38066) );
  HS65_LH_IVX2 U22340 ( .A(n38073), .Z(n38067) );
  HS65_LH_IVX2 U22341 ( .A(n38067), .Z(n38068) );
  HS65_LH_BFX2 U22342 ( .A(n38074), .Z(n38069) );
  HS65_LH_IVX2 U22343 ( .A(n38076), .Z(n38070) );
  HS65_LH_IVX2 U22344 ( .A(n38070), .Z(n38071) );
  HS65_LH_IVX2 U22345 ( .A(n38078), .Z(n38072) );
  HS65_LH_IVX2 U22346 ( .A(n38072), .Z(n38073) );
  HS65_LH_BFX2 U22347 ( .A(n38079), .Z(n38074) );
  HS65_LH_IVX2 U22348 ( .A(n38081), .Z(n38075) );
  HS65_LH_IVX2 U22349 ( .A(n38075), .Z(n38076) );
  HS65_LH_IVX2 U22350 ( .A(n38083), .Z(n38077) );
  HS65_LH_IVX2 U22351 ( .A(n38077), .Z(n38078) );
  HS65_LH_BFX2 U22352 ( .A(n38084), .Z(n38079) );
  HS65_LH_IVX2 U22353 ( .A(n38090), .Z(n38080) );
  HS65_LH_IVX2 U22354 ( .A(n38080), .Z(n38081) );
  HS65_LH_IVX2 U22355 ( .A(n38086), .Z(n38082) );
  HS65_LH_IVX2 U22356 ( .A(n38082), .Z(n38083) );
  HS65_LH_BFX2 U22357 ( .A(n38088), .Z(n38084) );
  HS65_LH_IVX2 U22358 ( .A(n1772), .Z(n38085) );
  HS65_LH_IVX2 U22359 ( .A(n38085), .Z(n38086) );
  HS65_LH_BFX2 U22360 ( .A(n16580), .Z(n38087) );
  HS65_LH_BFX2 U22361 ( .A(n38092), .Z(n38088) );
  HS65_LH_IVX2 U22362 ( .A(n1771), .Z(n38089) );
  HS65_LH_IVX2 U22363 ( .A(n38089), .Z(n38090) );
  HS65_LH_IVX2 U22364 ( .A(n38094), .Z(n38091) );
  HS65_LH_IVX2 U22365 ( .A(n38091), .Z(n38092) );
  HS65_LH_IVX2 U22366 ( .A(n38095), .Z(n38093) );
  HS65_LH_IVX2 U22367 ( .A(n38093), .Z(n38094) );
  HS65_LH_BFX2 U22368 ( .A(n38096), .Z(n38095) );
  HS65_LH_BFX2 U22369 ( .A(n38097), .Z(n38096) );
  HS65_LH_BFX2 U22370 ( .A(n17902), .Z(n38097) );
  HS65_LH_BFX2 U22371 ( .A(n38102), .Z(n38098) );
  HS65_LH_BFX2 U22372 ( .A(n38104), .Z(n38099) );
  HS65_LH_BFX2 U22373 ( .A(n38105), .Z(n38100) );
  HS65_LH_IVX2 U22374 ( .A(n38109), .Z(n38101) );
  HS65_LH_IVX2 U22375 ( .A(n38101), .Z(n38102) );
  HS65_LH_IVX2 U22376 ( .A(n38111), .Z(n38103) );
  HS65_LH_IVX2 U22377 ( .A(n38103), .Z(n38104) );
  HS65_LH_BFX2 U22378 ( .A(n38107), .Z(n38105) );
  HS65_LH_IVX2 U22379 ( .A(n38113), .Z(n38106) );
  HS65_LH_IVX2 U22380 ( .A(n38106), .Z(n38107) );
  HS65_LH_IVX2 U22381 ( .A(n38115), .Z(n38108) );
  HS65_LH_IVX2 U22383 ( .A(n38108), .Z(n38109) );
  HS65_LH_IVX2 U22384 ( .A(n38117), .Z(n38110) );
  HS65_LH_IVX2 U22385 ( .A(n38110), .Z(n38111) );
  HS65_LH_IVX2 U22386 ( .A(n38119), .Z(n38112) );
  HS65_LH_IVX2 U22387 ( .A(n38112), .Z(n38113) );
  HS65_LH_IVX2 U22388 ( .A(n38121), .Z(n38114) );
  HS65_LH_IVX2 U22389 ( .A(n38114), .Z(n38115) );
  HS65_LH_IVX2 U22390 ( .A(n38123), .Z(n38116) );
  HS65_LH_IVX2 U22391 ( .A(n38116), .Z(n38117) );
  HS65_LH_IVX2 U22392 ( .A(n38125), .Z(n38118) );
  HS65_LH_IVX2 U22393 ( .A(n38118), .Z(n38119) );
  HS65_LH_IVX2 U22394 ( .A(n38127), .Z(n38120) );
  HS65_LH_IVX2 U22395 ( .A(n38120), .Z(n38121) );
  HS65_LH_IVX2 U22396 ( .A(n38129), .Z(n38122) );
  HS65_LH_IVX2 U22397 ( .A(n38122), .Z(n38123) );
  HS65_LH_IVX2 U22398 ( .A(n38131), .Z(n38124) );
  HS65_LH_IVX2 U22399 ( .A(n38124), .Z(n38125) );
  HS65_LH_IVX2 U22400 ( .A(n38133), .Z(n38126) );
  HS65_LH_IVX2 U22401 ( .A(n38126), .Z(n38127) );
  HS65_LH_IVX2 U22402 ( .A(n38135), .Z(n38128) );
  HS65_LH_IVX2 U22403 ( .A(n38128), .Z(n38129) );
  HS65_LH_IVX2 U22404 ( .A(n38137), .Z(n38130) );
  HS65_LH_IVX2 U22405 ( .A(n38130), .Z(n38131) );
  HS65_LH_IVX2 U22406 ( .A(n38139), .Z(n38132) );
  HS65_LH_IVX2 U22407 ( .A(n38132), .Z(n38133) );
  HS65_LH_IVX2 U22408 ( .A(n38141), .Z(n38134) );
  HS65_LH_IVX2 U22409 ( .A(n38134), .Z(n38135) );
  HS65_LH_IVX2 U22410 ( .A(n38146), .Z(n38136) );
  HS65_LH_IVX2 U22411 ( .A(n38136), .Z(n38137) );
  HS65_LH_IVX2 U22412 ( .A(n38143), .Z(n38138) );
  HS65_LH_IVX2 U22413 ( .A(n38138), .Z(n38139) );
  HS65_LH_IVX2 U22414 ( .A(n38145), .Z(n38140) );
  HS65_LH_IVX2 U22415 ( .A(n38140), .Z(n38141) );
  HS65_LH_IVX2 U22416 ( .A(n38148), .Z(n38142) );
  HS65_LH_IVX2 U22417 ( .A(n38142), .Z(n38143) );
  HS65_LH_IVX2 U22418 ( .A(n38150), .Z(n38144) );
  HS65_LH_IVX2 U22419 ( .A(n38144), .Z(n38145) );
  HS65_LH_BFX2 U22420 ( .A(n38151), .Z(n38146) );
  HS65_LH_IVX2 U22421 ( .A(n38153), .Z(n38147) );
  HS65_LH_IVX2 U22422 ( .A(n38147), .Z(n38148) );
  HS65_LH_IVX2 U22423 ( .A(n38155), .Z(n38149) );
  HS65_LH_IVX2 U22424 ( .A(n38149), .Z(n38150) );
  HS65_LH_BFX2 U22425 ( .A(n38156), .Z(n38151) );
  HS65_LH_IVX2 U22426 ( .A(n38158), .Z(n38152) );
  HS65_LH_IVX2 U22427 ( .A(n38152), .Z(n38153) );
  HS65_LH_IVX2 U22428 ( .A(n38160), .Z(n38154) );
  HS65_LH_IVX2 U22429 ( .A(n38154), .Z(n38155) );
  HS65_LH_BFX2 U22430 ( .A(n38161), .Z(n38156) );
  HS65_LH_IVX2 U22431 ( .A(n38163), .Z(n38157) );
  HS65_LH_IVX2 U22432 ( .A(n38157), .Z(n38158) );
  HS65_LH_IVX2 U22433 ( .A(n38165), .Z(n38159) );
  HS65_LH_IVX2 U22434 ( .A(n38159), .Z(n38160) );
  HS65_LH_BFX2 U22435 ( .A(n38166), .Z(n38161) );
  HS65_LH_IVX2 U22436 ( .A(n38170), .Z(n38162) );
  HS65_LH_IVX2 U22437 ( .A(n38162), .Z(n38163) );
  HS65_LH_IVX2 U22438 ( .A(n38168), .Z(n38164) );
  HS65_LH_IVX2 U22439 ( .A(n38164), .Z(n38165) );
  HS65_LH_BFX2 U22440 ( .A(n38169), .Z(n38166) );
  HS65_LH_IVX2 U22441 ( .A(n38172), .Z(n38167) );
  HS65_LH_IVX2 U22442 ( .A(n38167), .Z(n38168) );
  HS65_LH_BFX2 U22443 ( .A(n38173), .Z(n38169) );
  HS65_LH_BFX2 U22444 ( .A(n38174), .Z(n38170) );
  HS65_LH_IVX2 U22445 ( .A(n1404), .Z(n38171) );
  HS65_LH_IVX2 U22446 ( .A(n38171), .Z(n38172) );
  HS65_LH_BFX2 U22447 ( .A(n38175), .Z(n38173) );
  HS65_LH_BFX2 U22448 ( .A(n38176), .Z(n38174) );
  HS65_LH_BFX2 U22449 ( .A(n38177), .Z(n38175) );
  HS65_LH_BFX2 U22450 ( .A(n1403), .Z(n38176) );
  HS65_LH_BFX2 U22451 ( .A(n38178), .Z(n38177) );
  HS65_LH_BFX2 U22452 ( .A(n38179), .Z(n38178) );
  HS65_LH_BFX2 U22453 ( .A(n38180), .Z(n38179) );
  HS65_LH_BFX2 U22454 ( .A(n17895), .Z(n38180) );
  HS65_LH_NAND4ABX3 U22455 ( .A(n17032), .B(n17031), .C(n17030), .D(n17029), 
        .Z(n1266) );
  HS65_LH_BFX2 U22456 ( .A(n38183), .Z(n38181) );
  HS65_LH_IVX2 U22457 ( .A(n38188), .Z(n38182) );
  HS65_LH_IVX2 U22458 ( .A(n38182), .Z(n38183) );
  HS65_LH_BFX2 U22459 ( .A(n1265), .Z(n38184) );
  HS65_LH_BFX2 U22460 ( .A(n38187), .Z(n38185) );
  HS65_LH_BFX2 U22461 ( .A(n38184), .Z(n38186) );
  HS65_LH_BFX2 U22462 ( .A(n38190), .Z(n38187) );
  HS65_LH_BFX2 U22463 ( .A(n38191), .Z(n38188) );
  HS65_LH_BFX2 U22464 ( .A(n38186), .Z(n38189) );
  HS65_LH_BFX2 U22465 ( .A(n38193), .Z(n38190) );
  HS65_LH_BFX2 U22466 ( .A(n38194), .Z(n38191) );
  HS65_LH_BFX2 U22467 ( .A(n38189), .Z(n38192) );
  HS65_LH_BFX2 U22468 ( .A(n38196), .Z(n38193) );
  HS65_LH_BFX2 U22469 ( .A(n38197), .Z(n38194) );
  HS65_LH_BFX2 U22470 ( .A(n38192), .Z(n38195) );
  HS65_LH_BFX2 U22471 ( .A(n38199), .Z(n38196) );
  HS65_LH_BFX2 U22472 ( .A(n38200), .Z(n38197) );
  HS65_LH_BFX2 U22473 ( .A(n38195), .Z(n38198) );
  HS65_LH_BFX2 U22474 ( .A(n38202), .Z(n38199) );
  HS65_LH_BFX2 U22475 ( .A(n38203), .Z(n38200) );
  HS65_LH_BFX2 U22476 ( .A(n38198), .Z(n38201) );
  HS65_LH_BFX2 U22477 ( .A(n38205), .Z(n38202) );
  HS65_LH_BFX2 U22478 ( .A(n38206), .Z(n38203) );
  HS65_LH_BFX2 U22479 ( .A(n38201), .Z(n38204) );
  HS65_LH_BFX2 U22480 ( .A(n38208), .Z(n38205) );
  HS65_LH_BFX2 U22481 ( .A(n38209), .Z(n38206) );
  HS65_LH_BFX2 U22482 ( .A(n38204), .Z(n38207) );
  HS65_LH_BFX2 U22483 ( .A(n38211), .Z(n38208) );
  HS65_LH_BFX2 U22484 ( .A(n38212), .Z(n38209) );
  HS65_LH_BFX2 U22485 ( .A(n38207), .Z(n38210) );
  HS65_LH_BFX2 U22486 ( .A(n38214), .Z(n38211) );
  HS65_LH_BFX2 U22487 ( .A(n38215), .Z(n38212) );
  HS65_LH_BFX2 U22488 ( .A(n38210), .Z(n38213) );
  HS65_LH_BFX2 U22489 ( .A(n38217), .Z(n38214) );
  HS65_LH_BFX2 U22490 ( .A(n38218), .Z(n38215) );
  HS65_LH_BFX2 U22491 ( .A(n38213), .Z(n38216) );
  HS65_LH_BFX2 U22492 ( .A(n38220), .Z(n38217) );
  HS65_LH_BFX2 U22493 ( .A(n38221), .Z(n38218) );
  HS65_LH_BFX2 U22494 ( .A(n38216), .Z(n38219) );
  HS65_LH_BFX2 U22495 ( .A(n38223), .Z(n38220) );
  HS65_LH_BFX2 U22496 ( .A(n38224), .Z(n38221) );
  HS65_LH_BFX2 U22497 ( .A(n38219), .Z(n38222) );
  HS65_LH_BFX2 U22498 ( .A(n38226), .Z(n38223) );
  HS65_LH_BFX2 U22499 ( .A(n38227), .Z(n38224) );
  HS65_LH_BFX2 U22500 ( .A(n38222), .Z(n38225) );
  HS65_LH_BFX2 U22501 ( .A(n38231), .Z(n38226) );
  HS65_LH_BFX2 U22502 ( .A(n38230), .Z(n38227) );
  HS65_LH_BFX2 U22503 ( .A(n17019), .Z(n38228) );
  HS65_LH_IVX2 U22504 ( .A(n1266), .Z(n38229) );
  HS65_LH_IVX2 U22505 ( .A(n38229), .Z(n38230) );
  HS65_LH_BFX2 U22506 ( .A(n38234), .Z(n38231) );
  HS65_LH_IVX2 U22507 ( .A(n38225), .Z(n38232) );
  HS65_LH_IVX2 U22508 ( .A(n38232), .Z(n38233) );
  HS65_LH_BFX2 U22509 ( .A(n38235), .Z(n38234) );
  HS65_LH_BFX2 U22510 ( .A(n38236), .Z(n38235) );
  HS65_LH_BFX2 U22511 ( .A(n38237), .Z(n38236) );
  HS65_LH_BFX2 U22512 ( .A(n17965), .Z(n38237) );
  HS65_LH_BFX2 U22513 ( .A(n38241), .Z(n38238) );
  HS65_LH_BFX2 U22514 ( .A(n38244), .Z(n38239) );
  HS65_LH_IVX2 U22515 ( .A(n38248), .Z(n38240) );
  HS65_LH_IVX2 U22516 ( .A(n38240), .Z(n38241) );
  HS65_LH_BFX2 U22517 ( .A(n38246), .Z(n38242) );
  HS65_LH_IVX2 U22518 ( .A(n38250), .Z(n38243) );
  HS65_LH_IVX2 U22519 ( .A(n38243), .Z(n38244) );
  HS65_LH_IVX2 U22520 ( .A(n38252), .Z(n38245) );
  HS65_LH_IVX2 U22521 ( .A(n38245), .Z(n38246) );
  HS65_LH_IVX2 U22522 ( .A(n38254), .Z(n38247) );
  HS65_LH_IVX2 U22523 ( .A(n38247), .Z(n38248) );
  HS65_LH_IVX2 U22524 ( .A(n38256), .Z(n38249) );
  HS65_LH_IVX2 U22525 ( .A(n38249), .Z(n38250) );
  HS65_LH_IVX2 U22526 ( .A(n38258), .Z(n38251) );
  HS65_LH_IVX2 U22527 ( .A(n38251), .Z(n38252) );
  HS65_LH_IVX2 U22528 ( .A(n38260), .Z(n38253) );
  HS65_LH_IVX2 U22529 ( .A(n38253), .Z(n38254) );
  HS65_LH_IVX2 U22530 ( .A(n38262), .Z(n38255) );
  HS65_LH_IVX2 U22531 ( .A(n38255), .Z(n38256) );
  HS65_LH_IVX2 U22532 ( .A(n38264), .Z(n38257) );
  HS65_LH_IVX2 U22533 ( .A(n38257), .Z(n38258) );
  HS65_LH_IVX2 U22534 ( .A(n38266), .Z(n38259) );
  HS65_LH_IVX2 U22535 ( .A(n38259), .Z(n38260) );
  HS65_LH_IVX2 U22536 ( .A(n38268), .Z(n38261) );
  HS65_LH_IVX2 U22537 ( .A(n38261), .Z(n38262) );
  HS65_LH_IVX2 U22538 ( .A(n38270), .Z(n38263) );
  HS65_LH_IVX2 U22539 ( .A(n38263), .Z(n38264) );
  HS65_LH_IVX2 U22540 ( .A(n38272), .Z(n38265) );
  HS65_LH_IVX2 U22541 ( .A(n38265), .Z(n38266) );
  HS65_LH_IVX2 U22542 ( .A(n38274), .Z(n38267) );
  HS65_LH_IVX2 U22543 ( .A(n38267), .Z(n38268) );
  HS65_LH_IVX2 U22544 ( .A(n38276), .Z(n38269) );
  HS65_LH_IVX2 U22545 ( .A(n38269), .Z(n38270) );
  HS65_LH_IVX2 U22546 ( .A(n38278), .Z(n38271) );
  HS65_LH_IVX2 U22547 ( .A(n38271), .Z(n38272) );
  HS65_LH_IVX2 U22548 ( .A(n38280), .Z(n38273) );
  HS65_LH_IVX2 U22549 ( .A(n38273), .Z(n38274) );
  HS65_LH_IVX2 U22550 ( .A(n38282), .Z(n38275) );
  HS65_LH_IVX2 U22551 ( .A(n38275), .Z(n38276) );
  HS65_LH_IVX2 U22552 ( .A(n38284), .Z(n38277) );
  HS65_LH_IVX2 U22553 ( .A(n38277), .Z(n38278) );
  HS65_LH_IVX2 U22554 ( .A(n38286), .Z(n38279) );
  HS65_LH_IVX2 U22555 ( .A(n38279), .Z(n38280) );
  HS65_LH_IVX2 U22556 ( .A(n38288), .Z(n38281) );
  HS65_LH_IVX2 U22557 ( .A(n38281), .Z(n38282) );
  HS65_LH_IVX2 U22558 ( .A(n38290), .Z(n38283) );
  HS65_LH_IVX2 U22559 ( .A(n38283), .Z(n38284) );
  HS65_LH_IVX2 U22560 ( .A(n38292), .Z(n38285) );
  HS65_LH_IVX2 U22561 ( .A(n38285), .Z(n38286) );
  HS65_LH_IVX2 U22562 ( .A(n38294), .Z(n38287) );
  HS65_LH_IVX2 U22563 ( .A(n38287), .Z(n38288) );
  HS65_LH_IVX2 U22565 ( .A(n38296), .Z(n38289) );
  HS65_LH_IVX2 U22566 ( .A(n38289), .Z(n38290) );
  HS65_LH_IVX2 U22567 ( .A(n38298), .Z(n38291) );
  HS65_LH_IVX2 U22568 ( .A(n38291), .Z(n38292) );
  HS65_LH_IVX2 U22569 ( .A(n38300), .Z(n38293) );
  HS65_LH_IVX2 U22570 ( .A(n38293), .Z(n38294) );
  HS65_LH_IVX2 U22571 ( .A(n38302), .Z(n38295) );
  HS65_LH_IVX2 U22572 ( .A(n38295), .Z(n38296) );
  HS65_LH_IVX2 U22573 ( .A(n38304), .Z(n38297) );
  HS65_LH_IVX2 U22574 ( .A(n38297), .Z(n38298) );
  HS65_LH_IVX2 U22575 ( .A(n38306), .Z(n38299) );
  HS65_LH_IVX2 U22576 ( .A(n38299), .Z(n38300) );
  HS65_LH_IVX2 U22577 ( .A(n38311), .Z(n38301) );
  HS65_LH_IVX2 U22578 ( .A(n38301), .Z(n38302) );
  HS65_LH_IVX2 U22579 ( .A(n38308), .Z(n38303) );
  HS65_LH_IVX2 U22580 ( .A(n38303), .Z(n38304) );
  HS65_LH_IVX2 U22581 ( .A(n38310), .Z(n38305) );
  HS65_LH_IVX2 U22582 ( .A(n38305), .Z(n38306) );
  HS65_LH_IVX2 U22583 ( .A(n38313), .Z(n38307) );
  HS65_LH_IVX2 U22584 ( .A(n38307), .Z(n38308) );
  HS65_LH_IVX2 U22585 ( .A(n38315), .Z(n38309) );
  HS65_LH_IVX2 U22586 ( .A(n38309), .Z(n38310) );
  HS65_LH_BFX2 U22587 ( .A(n38316), .Z(n38311) );
  HS65_LH_IVX2 U22588 ( .A(n38318), .Z(n38312) );
  HS65_LH_IVX2 U22589 ( .A(n38312), .Z(n38313) );
  HS65_LH_IVX2 U22590 ( .A(n38320), .Z(n38314) );
  HS65_LH_IVX2 U22591 ( .A(n38314), .Z(n38315) );
  HS65_LH_BFX2 U22592 ( .A(n38321), .Z(n38316) );
  HS65_LH_IVX2 U22593 ( .A(n1173), .Z(n38317) );
  HS65_LH_IVX2 U22594 ( .A(n38317), .Z(n38318) );
  HS65_LH_IVX2 U22595 ( .A(n1174), .Z(n38319) );
  HS65_LH_IVX2 U22596 ( .A(n38319), .Z(n38320) );
  HS65_LH_BFX2 U22597 ( .A(n38322), .Z(n38321) );
  HS65_LH_BFX2 U22598 ( .A(n38323), .Z(n38322) );
  HS65_LH_BFX2 U22599 ( .A(n38324), .Z(n38323) );
  HS65_LH_BFX2 U22600 ( .A(n38325), .Z(n38324) );
  HS65_LH_BFX2 U22601 ( .A(n17955), .Z(n38325) );
  HS65_LH_NAND4ABX3 U22602 ( .A(n17109), .B(n17108), .C(n17107), .D(n17106), 
        .Z(n1197) );
  HS65_LH_IVX2 U22603 ( .A(n38332), .Z(n38326) );
  HS65_LH_IVX2 U22604 ( .A(n38326), .Z(n38327) );
  HS65_LH_NAND4ABX3 U22605 ( .A(n17096), .B(n17095), .C(n17094), .D(n17093), 
        .Z(n1196) );
  HS65_LH_BFX2 U22606 ( .A(n1196), .Z(n38328) );
  HS65_LH_BFX2 U22607 ( .A(n38331), .Z(n38329) );
  HS65_LH_BFX2 U22608 ( .A(n38328), .Z(n38330) );
  HS65_LH_BFX2 U22609 ( .A(n38334), .Z(n38331) );
  HS65_LH_BFX2 U22610 ( .A(n38335), .Z(n38332) );
  HS65_LH_BFX2 U22611 ( .A(n38330), .Z(n38333) );
  HS65_LH_BFX2 U22612 ( .A(n38337), .Z(n38334) );
  HS65_LH_BFX2 U22613 ( .A(n38338), .Z(n38335) );
  HS65_LH_BFX2 U22614 ( .A(n38333), .Z(n38336) );
  HS65_LH_BFX2 U22615 ( .A(n38340), .Z(n38337) );
  HS65_LH_BFX2 U22616 ( .A(n38341), .Z(n38338) );
  HS65_LH_BFX2 U22617 ( .A(n38336), .Z(n38339) );
  HS65_LH_BFX2 U22618 ( .A(n38343), .Z(n38340) );
  HS65_LH_BFX2 U22619 ( .A(n38344), .Z(n38341) );
  HS65_LH_BFX2 U22620 ( .A(n38339), .Z(n38342) );
  HS65_LH_BFX2 U22621 ( .A(n38346), .Z(n38343) );
  HS65_LH_BFX2 U22622 ( .A(n38347), .Z(n38344) );
  HS65_LH_BFX2 U22623 ( .A(n38342), .Z(n38345) );
  HS65_LH_BFX2 U22624 ( .A(n38349), .Z(n38346) );
  HS65_LH_BFX2 U22625 ( .A(n38350), .Z(n38347) );
  HS65_LH_BFX2 U22626 ( .A(n38345), .Z(n38348) );
  HS65_LH_BFX2 U22627 ( .A(n38352), .Z(n38349) );
  HS65_LH_BFX2 U22628 ( .A(n38353), .Z(n38350) );
  HS65_LH_BFX2 U22629 ( .A(n38348), .Z(n38351) );
  HS65_LH_BFX2 U22630 ( .A(n38355), .Z(n38352) );
  HS65_LH_BFX2 U22631 ( .A(n38356), .Z(n38353) );
  HS65_LH_BFX2 U22632 ( .A(n38351), .Z(n38354) );
  HS65_LH_BFX2 U22633 ( .A(n38358), .Z(n38355) );
  HS65_LH_BFX2 U22634 ( .A(n38359), .Z(n38356) );
  HS65_LH_BFX2 U22635 ( .A(n38354), .Z(n38357) );
  HS65_LH_BFX2 U22636 ( .A(n38361), .Z(n38358) );
  HS65_LH_BFX2 U22637 ( .A(n38362), .Z(n38359) );
  HS65_LH_BFX2 U22638 ( .A(n38357), .Z(n38360) );
  HS65_LH_BFX2 U22639 ( .A(n38364), .Z(n38361) );
  HS65_LH_BFX2 U22640 ( .A(n38365), .Z(n38362) );
  HS65_LH_BFX2 U22641 ( .A(n38360), .Z(n38363) );
  HS65_LH_BFX2 U22642 ( .A(n38367), .Z(n38364) );
  HS65_LH_BFX2 U22643 ( .A(n38368), .Z(n38365) );
  HS65_LH_BFX2 U22644 ( .A(n38363), .Z(n38366) );
  HS65_LH_BFX2 U22645 ( .A(n38370), .Z(n38367) );
  HS65_LH_BFX2 U22646 ( .A(n38371), .Z(n38368) );
  HS65_LH_BFX2 U22647 ( .A(n38366), .Z(n38369) );
  HS65_LH_BFX2 U22648 ( .A(n38377), .Z(n38370) );
  HS65_LH_BFX2 U22649 ( .A(n38374), .Z(n38371) );
  HS65_LH_BFX2 U22650 ( .A(n38369), .Z(n38372) );
  HS65_LH_IVX2 U22651 ( .A(n1197), .Z(n38373) );
  HS65_LH_IVX2 U22652 ( .A(n38373), .Z(n38374) );
  HS65_LH_IVX2 U22653 ( .A(n38372), .Z(n38375) );
  HS65_LH_IVX2 U22654 ( .A(n38375), .Z(n38376) );
  HS65_LH_BFX2 U22655 ( .A(n38378), .Z(n38377) );
  HS65_LH_BFX2 U22656 ( .A(n38379), .Z(n38378) );
  HS65_LH_BFX2 U22657 ( .A(n38380), .Z(n38379) );
  HS65_LH_BFX2 U22658 ( .A(n38381), .Z(n38380) );
  HS65_LH_BFX2 U22659 ( .A(n17941), .Z(n38381) );
  HS65_LH_IVX2 U22660 ( .A(n38388), .Z(n38382) );
  HS65_LH_IVX2 U22661 ( .A(n38382), .Z(n38383) );
  HS65_LH_BFX2 U22662 ( .A(n1817), .Z(n38384) );
  HS65_LH_BFX2 U22663 ( .A(n38387), .Z(n38385) );
  HS65_LH_BFX2 U22664 ( .A(n38384), .Z(n38386) );
  HS65_LH_BFX2 U22665 ( .A(n38390), .Z(n38387) );
  HS65_LH_BFX2 U22666 ( .A(n38391), .Z(n38388) );
  HS65_LH_BFX2 U22667 ( .A(n38386), .Z(n38389) );
  HS65_LH_BFX2 U22668 ( .A(n38393), .Z(n38390) );
  HS65_LH_BFX2 U22669 ( .A(n38394), .Z(n38391) );
  HS65_LH_BFX2 U22670 ( .A(n38389), .Z(n38392) );
  HS65_LH_BFX2 U22671 ( .A(n38396), .Z(n38393) );
  HS65_LH_BFX2 U22672 ( .A(n38397), .Z(n38394) );
  HS65_LH_BFX2 U22673 ( .A(n38392), .Z(n38395) );
  HS65_LH_BFX2 U22674 ( .A(n38399), .Z(n38396) );
  HS65_LH_BFX2 U22675 ( .A(n38400), .Z(n38397) );
  HS65_LH_BFX2 U22676 ( .A(n38395), .Z(n38398) );
  HS65_LH_BFX2 U22677 ( .A(n38402), .Z(n38399) );
  HS65_LH_BFX2 U22678 ( .A(n38403), .Z(n38400) );
  HS65_LH_BFX2 U22679 ( .A(n38398), .Z(n38401) );
  HS65_LH_BFX2 U22680 ( .A(n38405), .Z(n38402) );
  HS65_LH_BFX2 U22681 ( .A(n38406), .Z(n38403) );
  HS65_LH_BFX2 U22682 ( .A(n38401), .Z(n38404) );
  HS65_LH_BFX2 U22683 ( .A(n38408), .Z(n38405) );
  HS65_LH_BFX2 U22684 ( .A(n38409), .Z(n38406) );
  HS65_LH_BFX2 U22685 ( .A(n38404), .Z(n38407) );
  HS65_LH_BFX2 U22686 ( .A(n38411), .Z(n38408) );
  HS65_LH_BFX2 U22687 ( .A(n38412), .Z(n38409) );
  HS65_LH_BFX2 U22688 ( .A(n38407), .Z(n38410) );
  HS65_LH_BFX2 U22689 ( .A(n38414), .Z(n38411) );
  HS65_LH_BFX2 U22690 ( .A(n38415), .Z(n38412) );
  HS65_LH_BFX2 U22691 ( .A(n38410), .Z(n38413) );
  HS65_LH_BFX2 U22692 ( .A(n38417), .Z(n38414) );
  HS65_LH_BFX2 U22693 ( .A(n38418), .Z(n38415) );
  HS65_LH_BFX2 U22694 ( .A(n38413), .Z(n38416) );
  HS65_LH_BFX2 U22695 ( .A(n38420), .Z(n38417) );
  HS65_LH_BFX2 U22696 ( .A(n38421), .Z(n38418) );
  HS65_LH_BFX2 U22697 ( .A(n38416), .Z(n38419) );
  HS65_LH_BFX2 U22698 ( .A(n38423), .Z(n38420) );
  HS65_LH_BFX2 U22699 ( .A(n38424), .Z(n38421) );
  HS65_LH_BFX2 U22700 ( .A(n38419), .Z(n38422) );
  HS65_LH_BFX2 U22701 ( .A(n38426), .Z(n38423) );
  HS65_LH_BFX2 U22702 ( .A(n38427), .Z(n38424) );
  HS65_LH_BFX2 U22703 ( .A(n38422), .Z(n38425) );
  HS65_LH_BFX2 U22704 ( .A(n38431), .Z(n38426) );
  HS65_LH_BFX2 U22705 ( .A(n38432), .Z(n38427) );
  HS65_LH_BFX2 U22706 ( .A(n16539), .Z(n38428) );
  HS65_LH_IVX2 U22707 ( .A(n38425), .Z(n38429) );
  HS65_LH_IVX2 U22708 ( .A(n38429), .Z(n38430) );
  HS65_LH_BFX2 U22709 ( .A(n38433), .Z(n38431) );
  HS65_LH_BFX2 U22710 ( .A(n1818), .Z(n38432) );
  HS65_LH_BFX2 U22711 ( .A(n38434), .Z(n38433) );
  HS65_LH_BFX2 U22712 ( .A(n38435), .Z(n38434) );
  HS65_LH_BFX2 U22713 ( .A(n38436), .Z(n38435) );
  HS65_LH_BFX2 U22714 ( .A(n17880), .Z(n38436) );
  HS65_LH_BFX2 U22715 ( .A(n38439), .Z(n38437) );
  HS65_LH_IVX2 U22716 ( .A(n38444), .Z(n38438) );
  HS65_LH_IVX2 U22717 ( .A(n38438), .Z(n38439) );
  HS65_LH_NAND2X2 U22718 ( .A(n16554), .B(n16553), .Z(n16562) );
  HS65_LH_BFX2 U22719 ( .A(n16562), .Z(n38440) );
  HS65_LH_BFX2 U22720 ( .A(n38442), .Z(n38441) );
  HS65_LH_BFX2 U22721 ( .A(n38445), .Z(n38442) );
  HS65_LH_BFX2 U22722 ( .A(n38446), .Z(n38443) );
  HS65_LH_BFX2 U22723 ( .A(n38447), .Z(n38444) );
  HS65_LH_BFX2 U22724 ( .A(n38448), .Z(n38445) );
  HS65_LH_BFX2 U22725 ( .A(n38449), .Z(n38446) );
  HS65_LH_BFX2 U22726 ( .A(n38450), .Z(n38447) );
  HS65_LH_BFX2 U22727 ( .A(n38451), .Z(n38448) );
  HS65_LH_BFX2 U22728 ( .A(n38452), .Z(n38449) );
  HS65_LH_BFX2 U22729 ( .A(n38453), .Z(n38450) );
  HS65_LH_BFX2 U22730 ( .A(n38454), .Z(n38451) );
  HS65_LH_BFX2 U22731 ( .A(n38455), .Z(n38452) );
  HS65_LH_BFX2 U22732 ( .A(n38456), .Z(n38453) );
  HS65_LH_BFX2 U22733 ( .A(n38457), .Z(n38454) );
  HS65_LH_BFX2 U22734 ( .A(n38458), .Z(n38455) );
  HS65_LH_BFX2 U22735 ( .A(n38459), .Z(n38456) );
  HS65_LH_BFX2 U22736 ( .A(n38460), .Z(n38457) );
  HS65_LH_BFX2 U22737 ( .A(n38461), .Z(n38458) );
  HS65_LH_BFX2 U22738 ( .A(n38462), .Z(n38459) );
  HS65_LH_BFX2 U22739 ( .A(n38463), .Z(n38460) );
  HS65_LH_BFX2 U22740 ( .A(n38464), .Z(n38461) );
  HS65_LH_BFX2 U22741 ( .A(n38465), .Z(n38462) );
  HS65_LH_BFX2 U22742 ( .A(n38466), .Z(n38463) );
  HS65_LH_BFX2 U22743 ( .A(n38467), .Z(n38464) );
  HS65_LH_BFX2 U22744 ( .A(n38468), .Z(n38465) );
  HS65_LH_BFX2 U22745 ( .A(n38469), .Z(n38466) );
  HS65_LH_BFX2 U22746 ( .A(n38470), .Z(n38467) );
  HS65_LH_BFX2 U22747 ( .A(n38471), .Z(n38468) );
  HS65_LH_BFX2 U22748 ( .A(n38472), .Z(n38469) );
  HS65_LH_BFX2 U22749 ( .A(n38473), .Z(n38470) );
  HS65_LH_BFX2 U22750 ( .A(n38474), .Z(n38471) );
  HS65_LH_BFX2 U22751 ( .A(n38475), .Z(n38472) );
  HS65_LH_BFX2 U22752 ( .A(n38476), .Z(n38473) );
  HS65_LH_BFX2 U22753 ( .A(n38477), .Z(n38474) );
  HS65_LH_BFX2 U22754 ( .A(n38478), .Z(n38475) );
  HS65_LH_BFX2 U22755 ( .A(n38479), .Z(n38476) );
  HS65_LH_BFX2 U22756 ( .A(n38480), .Z(n38477) );
  HS65_LH_BFX2 U22757 ( .A(n38481), .Z(n38478) );
  HS65_LH_BFX2 U22758 ( .A(n38482), .Z(n38479) );
  HS65_LH_BFX2 U22759 ( .A(n38483), .Z(n38480) );
  HS65_LH_BFX2 U22760 ( .A(n38484), .Z(n38481) );
  HS65_LH_BFX2 U22761 ( .A(n38485), .Z(n38482) );
  HS65_LH_BFX2 U22762 ( .A(n38486), .Z(n38483) );
  HS65_LH_BFX2 U22763 ( .A(n1795), .Z(n38484) );
  HS65_LH_BFX2 U22764 ( .A(n38487), .Z(n38485) );
  HS65_LH_BFX2 U22765 ( .A(n38488), .Z(n38486) );
  HS65_LH_BFX2 U22766 ( .A(n38489), .Z(n38487) );
  HS65_LH_BFX2 U22767 ( .A(n38490), .Z(n38488) );
  HS65_LH_BFX2 U22768 ( .A(n1794), .Z(n38489) );
  HS65_LH_BFX2 U22769 ( .A(n38491), .Z(n38490) );
  HS65_LH_BFX2 U22770 ( .A(n38492), .Z(n38491) );
  HS65_LH_BFX2 U22771 ( .A(n17973), .Z(n38492) );
  HS65_LH_BFX2 U22772 ( .A(n38495), .Z(n38493) );
  HS65_LH_IVX2 U22773 ( .A(n38506), .Z(n38494) );
  HS65_LH_IVX2 U22774 ( .A(n38494), .Z(n38495) );
  HS65_LH_BFX2 U22775 ( .A(n38499), .Z(n38496) );
  HS65_LH_BFX2 U22776 ( .A(n38501), .Z(n38497) );
  HS65_LH_IVX2 U22777 ( .A(n39511), .Z(n38498) );
  HS65_LH_IVX2 U22778 ( .A(n38498), .Z(n38499) );
  HS65_LH_IVX2 U22779 ( .A(n38507), .Z(n38500) );
  HS65_LH_IVX2 U22780 ( .A(n38500), .Z(n38501) );
  HS65_LH_BFX2 U22781 ( .A(n17783), .Z(n38502) );
  HS65_LH_BFX2 U22782 ( .A(n17782), .Z(n38503) );
  HS65_LH_BFX2 U22783 ( .A(n17781), .Z(n38504) );
  HS65_LH_BFX2 U22784 ( .A(n38502), .Z(n38505) );
  HS65_LH_BFX2 U22785 ( .A(n38509), .Z(n38506) );
  HS65_LH_BFX2 U22786 ( .A(n38510), .Z(n38507) );
  HS65_LH_BFX2 U22787 ( .A(n38505), .Z(n38508) );
  HS65_LH_BFX2 U22788 ( .A(n38512), .Z(n38509) );
  HS65_LH_BFX2 U22789 ( .A(n38513), .Z(n38510) );
  HS65_LH_BFX2 U22790 ( .A(n38508), .Z(n38511) );
  HS65_LH_BFX2 U22791 ( .A(n38515), .Z(n38512) );
  HS65_LH_BFX2 U22792 ( .A(n38516), .Z(n38513) );
  HS65_LH_BFX2 U22793 ( .A(n38511), .Z(n38514) );
  HS65_LH_BFX2 U22794 ( .A(n38518), .Z(n38515) );
  HS65_LH_BFX2 U22795 ( .A(n38519), .Z(n38516) );
  HS65_LH_BFX2 U22796 ( .A(n38514), .Z(n38517) );
  HS65_LH_BFX2 U22797 ( .A(n38521), .Z(n38518) );
  HS65_LH_BFX2 U22798 ( .A(n38522), .Z(n38519) );
  HS65_LH_BFX2 U22799 ( .A(n38517), .Z(n38520) );
  HS65_LH_BFX2 U22800 ( .A(n38524), .Z(n38521) );
  HS65_LH_BFX2 U22801 ( .A(n38525), .Z(n38522) );
  HS65_LH_BFX2 U22802 ( .A(n38520), .Z(n38523) );
  HS65_LH_BFX2 U22803 ( .A(n38527), .Z(n38524) );
  HS65_LH_BFX2 U22804 ( .A(n38528), .Z(n38525) );
  HS65_LH_BFX2 U22805 ( .A(n38523), .Z(n38526) );
  HS65_LH_BFX2 U22806 ( .A(n38530), .Z(n38527) );
  HS65_LH_BFX2 U22807 ( .A(n38531), .Z(n38528) );
  HS65_LH_BFX2 U22808 ( .A(n38526), .Z(n38529) );
  HS65_LH_BFX2 U22809 ( .A(n38533), .Z(n38530) );
  HS65_LH_BFX2 U22810 ( .A(n38534), .Z(n38531) );
  HS65_LH_BFX2 U22811 ( .A(n38529), .Z(n38532) );
  HS65_LH_BFX2 U22812 ( .A(n38536), .Z(n38533) );
  HS65_LH_BFX2 U22813 ( .A(n38537), .Z(n38534) );
  HS65_LH_BFX2 U22814 ( .A(n38532), .Z(n38535) );
  HS65_LH_BFX2 U22815 ( .A(n38539), .Z(n38536) );
  HS65_LH_BFX2 U22816 ( .A(n38540), .Z(n38537) );
  HS65_LH_BFX2 U22817 ( .A(n38535), .Z(n38538) );
  HS65_LH_BFX2 U22818 ( .A(n38542), .Z(n38539) );
  HS65_LH_BFX2 U22819 ( .A(n38543), .Z(n38540) );
  HS65_LH_BFX2 U22820 ( .A(n38538), .Z(n38541) );
  HS65_LH_BFX2 U22822 ( .A(n38545), .Z(n38542) );
  HS65_LH_BFX2 U22823 ( .A(n38546), .Z(n38543) );
  HS65_LH_BFX2 U22824 ( .A(n38541), .Z(n38544) );
  HS65_LH_BFX2 U22825 ( .A(n38548), .Z(n38545) );
  HS65_LH_BFX2 U22826 ( .A(n38549), .Z(n38546) );
  HS65_LH_BFX2 U22827 ( .A(n38544), .Z(n38547) );
  HS65_LH_BFX2 U22828 ( .A(n38551), .Z(n38548) );
  HS65_LH_BFX2 U22829 ( .A(n38552), .Z(n38549) );
  HS65_LH_BFX2 U22830 ( .A(n38547), .Z(n38550) );
  HS65_LH_BFX2 U22831 ( .A(n38554), .Z(n38551) );
  HS65_LH_BFX2 U22832 ( .A(n38555), .Z(n38552) );
  HS65_LH_BFX2 U22833 ( .A(n38550), .Z(n38553) );
  HS65_LH_BFX2 U22834 ( .A(n38557), .Z(n38554) );
  HS65_LH_BFX2 U22835 ( .A(n38558), .Z(n38555) );
  HS65_LH_BFX2 U22836 ( .A(n38553), .Z(n38556) );
  HS65_LH_BFX2 U22837 ( .A(n38564), .Z(n38557) );
  HS65_LH_BFX2 U22838 ( .A(n38561), .Z(n38558) );
  HS65_LH_BFX2 U22839 ( .A(n38556), .Z(n38559) );
  HS65_LH_IVX2 U22840 ( .A(n17784), .Z(n38560) );
  HS65_LH_IVX2 U22841 ( .A(n38560), .Z(n38561) );
  HS65_LH_IVX2 U22842 ( .A(n38559), .Z(n38562) );
  HS65_LH_IVX2 U22843 ( .A(n38562), .Z(n38563) );
  HS65_LH_BFX2 U22844 ( .A(n17687), .Z(n38564) );
  HS65_LH_BFX2 U22845 ( .A(n15724), .Z(n38565) );
  HS65_LH_BFX2 U22846 ( .A(n38567), .Z(n38566) );
  HS65_LH_BFX2 U22847 ( .A(n38568), .Z(n38567) );
  HS65_LH_BFX2 U22848 ( .A(n38569), .Z(n38568) );
  HS65_LH_BFX2 U22849 ( .A(n38570), .Z(n38569) );
  HS65_LH_BFX2 U22850 ( .A(n38571), .Z(n38570) );
  HS65_LH_BFX2 U22851 ( .A(n38572), .Z(n38571) );
  HS65_LH_BFX2 U22852 ( .A(n38573), .Z(n38572) );
  HS65_LH_BFX2 U22853 ( .A(n38574), .Z(n38573) );
  HS65_LH_BFX2 U22854 ( .A(n38575), .Z(n38574) );
  HS65_LH_BFX2 U22855 ( .A(n38577), .Z(n38575) );
  HS65_LH_IVX2 U22856 ( .A(n15427), .Z(n38576) );
  HS65_LH_IVX2 U22857 ( .A(n38576), .Z(n38577) );
  HS65_LH_BFX2 U22858 ( .A(n38580), .Z(n38578) );
  HS65_LH_BFX2 U22859 ( .A(n38582), .Z(n38579) );
  HS65_LH_BFX2 U22860 ( .A(n38581), .Z(n38580) );
  HS65_LH_BFX2 U22861 ( .A(n32337), .Z(n38581) );
  HS65_LH_BFX2 U22862 ( .A(n29559), .Z(n38582) );
  HS65_LH_BFX2 U22863 ( .A(n38584), .Z(n38583) );
  HS65_LH_BFX2 U22864 ( .A(n38585), .Z(n38584) );
  HS65_LH_BFX2 U22865 ( .A(n38586), .Z(n38585) );
  HS65_LH_BFX2 U22866 ( .A(n38587), .Z(n38586) );
  HS65_LH_BFX2 U22867 ( .A(n38588), .Z(n38587) );
  HS65_LH_BFX2 U22869 ( .A(n38589), .Z(n38588) );
  HS65_LH_BFX2 U22870 ( .A(n38590), .Z(n38589) );
  HS65_LH_BFX2 U22871 ( .A(n38591), .Z(n38590) );
  HS65_LH_BFX2 U22872 ( .A(n38592), .Z(n38591) );
  HS65_LH_BFX2 U22873 ( .A(n38593), .Z(n38592) );
  HS65_LH_BFX2 U22874 ( .A(n38594), .Z(n38593) );
  HS65_LH_BFX2 U22875 ( .A(n38595), .Z(n38594) );
  HS65_LH_BFX2 U22876 ( .A(n38596), .Z(n38595) );
  HS65_LH_BFX2 U22877 ( .A(n38597), .Z(n38596) );
  HS65_LH_BFX2 U22878 ( .A(n38598), .Z(n38597) );
  HS65_LH_BFX2 U22879 ( .A(n38599), .Z(n38598) );
  HS65_LH_BFX2 U22880 ( .A(n38600), .Z(n38599) );
  HS65_LH_BFX2 U22881 ( .A(n38601), .Z(n38600) );
  HS65_LH_BFX2 U22882 ( .A(n38602), .Z(n38601) );
  HS65_LH_BFX2 U22883 ( .A(n38603), .Z(n38602) );
  HS65_LH_BFX2 U22884 ( .A(n17572), .Z(n38603) );
  HS65_LH_BFX2 U22885 ( .A(n38605), .Z(n38604) );
  HS65_LH_BFX2 U22886 ( .A(n38606), .Z(n38605) );
  HS65_LH_BFX2 U22887 ( .A(n38607), .Z(n38606) );
  HS65_LH_BFX2 U22888 ( .A(n38608), .Z(n38607) );
  HS65_LH_BFX2 U22889 ( .A(n38609), .Z(n38608) );
  HS65_LH_BFX2 U22890 ( .A(n38610), .Z(n38609) );
  HS65_LH_BFX2 U22891 ( .A(n38611), .Z(n38610) );
  HS65_LH_BFX2 U22892 ( .A(n38612), .Z(n38611) );
  HS65_LH_BFX2 U22893 ( .A(n38613), .Z(n38612) );
  HS65_LH_BFX2 U22894 ( .A(n38614), .Z(n38613) );
  HS65_LH_BFX2 U22895 ( .A(n38615), .Z(n38614) );
  HS65_LH_BFX2 U22896 ( .A(n38616), .Z(n38615) );
  HS65_LH_BFX2 U22897 ( .A(n38617), .Z(n38616) );
  HS65_LH_BFX2 U22898 ( .A(n38618), .Z(n38617) );
  HS65_LH_BFX2 U22899 ( .A(n38619), .Z(n38618) );
  HS65_LH_BFX2 U22900 ( .A(n38620), .Z(n38619) );
  HS65_LH_BFX2 U22901 ( .A(n38621), .Z(n38620) );
  HS65_LH_BFX2 U22903 ( .A(n38622), .Z(n38621) );
  HS65_LH_BFX2 U22904 ( .A(n38623), .Z(n38622) );
  HS65_LH_BFX2 U22905 ( .A(n38624), .Z(n38623) );
  HS65_LH_BFX2 U22906 ( .A(n17579), .Z(n38624) );
  HS65_LH_IVX2 U22907 ( .A(n38627), .Z(n38625) );
  HS65_LH_IVX2 U22908 ( .A(n38625), .Z(n38626) );
  HS65_LH_BFX2 U22909 ( .A(n38628), .Z(n38627) );
  HS65_LH_BFX2 U22910 ( .A(n38629), .Z(n38628) );
  HS65_LH_BFX2 U22911 ( .A(n38630), .Z(n38629) );
  HS65_LH_BFX2 U22912 ( .A(n38631), .Z(n38630) );
  HS65_LH_BFX2 U22913 ( .A(n38632), .Z(n38631) );
  HS65_LH_BFX2 U22914 ( .A(n38633), .Z(n38632) );
  HS65_LH_BFX2 U22915 ( .A(n38634), .Z(n38633) );
  HS65_LH_BFX2 U22916 ( .A(n38635), .Z(n38634) );
  HS65_LH_BFX2 U22917 ( .A(n38636), .Z(n38635) );
  HS65_LH_BFX2 U22918 ( .A(n38637), .Z(n38636) );
  HS65_LH_BFX2 U22919 ( .A(n38638), .Z(n38637) );
  HS65_LH_BFX2 U22920 ( .A(n38639), .Z(n38638) );
  HS65_LH_BFX2 U22921 ( .A(n38640), .Z(n38639) );
  HS65_LH_BFX2 U22922 ( .A(n38641), .Z(n38640) );
  HS65_LH_BFX2 U22923 ( .A(n38642), .Z(n38641) );
  HS65_LH_BFX2 U22924 ( .A(n38643), .Z(n38642) );
  HS65_LH_BFX2 U22925 ( .A(n38644), .Z(n38643) );
  HS65_LH_BFX2 U22926 ( .A(n38645), .Z(n38644) );
  HS65_LH_BFX2 U22927 ( .A(n38646), .Z(n38645) );
  HS65_LH_BFX2 U22928 ( .A(n38647), .Z(n38646) );
  HS65_LH_BFX2 U22929 ( .A(n17633), .Z(n38647) );
  HS65_LH_BFX2 U22930 ( .A(n38649), .Z(n38648) );
  HS65_LH_BFX2 U22931 ( .A(n38650), .Z(n38649) );
  HS65_LH_BFX2 U22932 ( .A(n38651), .Z(n38650) );
  HS65_LH_BFX2 U22933 ( .A(n38652), .Z(n38651) );
  HS65_LH_BFX2 U22934 ( .A(n38653), .Z(n38652) );
  HS65_LH_BFX2 U22935 ( .A(n38654), .Z(n38653) );
  HS65_LH_BFX2 U22936 ( .A(n38655), .Z(n38654) );
  HS65_LH_BFX2 U22937 ( .A(n38656), .Z(n38655) );
  HS65_LH_BFX2 U22938 ( .A(n38657), .Z(n38656) );
  HS65_LH_BFX2 U22939 ( .A(n38658), .Z(n38657) );
  HS65_LH_BFX2 U22940 ( .A(n38659), .Z(n38658) );
  HS65_LH_BFX2 U22941 ( .A(n38660), .Z(n38659) );
  HS65_LH_BFX2 U22942 ( .A(n38661), .Z(n38660) );
  HS65_LH_BFX2 U22943 ( .A(n38662), .Z(n38661) );
  HS65_LH_BFX2 U22944 ( .A(n38663), .Z(n38662) );
  HS65_LH_BFX2 U22945 ( .A(n38664), .Z(n38663) );
  HS65_LH_BFX2 U22946 ( .A(n38665), .Z(n38664) );
  HS65_LH_BFX2 U22947 ( .A(n38666), .Z(n38665) );
  HS65_LH_BFX2 U22948 ( .A(n38667), .Z(n38666) );
  HS65_LH_BFX2 U22949 ( .A(n38668), .Z(n38667) );
  HS65_LH_BFX2 U22950 ( .A(n38669), .Z(n38668) );
  HS65_LH_BFX2 U22951 ( .A(n17732), .Z(n38669) );
  HS65_LH_BFX2 U22952 ( .A(n38671), .Z(n38670) );
  HS65_LH_BFX2 U22953 ( .A(n38672), .Z(n38671) );
  HS65_LH_BFX2 U22954 ( .A(n38673), .Z(n38672) );
  HS65_LH_BFX2 U22955 ( .A(n38674), .Z(n38673) );
  HS65_LH_BFX2 U22956 ( .A(n38675), .Z(n38674) );
  HS65_LH_BFX2 U22957 ( .A(n40602), .Z(n38675) );
  HS65_LH_BFX2 U22958 ( .A(n38677), .Z(n38676) );
  HS65_LH_BFX2 U22959 ( .A(n38678), .Z(n38677) );
  HS65_LH_BFX2 U22960 ( .A(n38679), .Z(n38678) );
  HS65_LH_BFX2 U22961 ( .A(n38680), .Z(n38679) );
  HS65_LH_BFX2 U22962 ( .A(n38681), .Z(n38680) );
  HS65_LH_BFX2 U22963 ( .A(n38682), .Z(n38681) );
  HS65_LH_BFX2 U22964 ( .A(n38683), .Z(n38682) );
  HS65_LH_BFX2 U22965 ( .A(n38684), .Z(n38683) );
  HS65_LH_BFX2 U22966 ( .A(n38685), .Z(n38684) );
  HS65_LH_BFX2 U22967 ( .A(n38686), .Z(n38685) );
  HS65_LH_BFX2 U22968 ( .A(n38687), .Z(n38686) );
  HS65_LH_BFX2 U22969 ( .A(n38688), .Z(n38687) );
  HS65_LH_BFX2 U22970 ( .A(n38689), .Z(n38688) );
  HS65_LH_BFX2 U22971 ( .A(n38690), .Z(n38689) );
  HS65_LH_BFX2 U22972 ( .A(n38691), .Z(n38690) );
  HS65_LH_BFX2 U22973 ( .A(n38692), .Z(n38691) );
  HS65_LH_BFX2 U22974 ( .A(n38693), .Z(n38692) );
  HS65_LH_BFX2 U22975 ( .A(n38694), .Z(n38693) );
  HS65_LH_BFX2 U22976 ( .A(n38695), .Z(n38694) );
  HS65_LH_BFX2 U22977 ( .A(n38696), .Z(n38695) );
  HS65_LH_BFX2 U22978 ( .A(n14482), .Z(n38696) );
  HS65_LH_BFX2 U22979 ( .A(n18081), .Z(n38697) );
  HS65_LH_BFX2 U22980 ( .A(n17724), .Z(n38698) );
  HS65_LH_BFX2 U22981 ( .A(n17703), .Z(n38699) );
  HS65_LH_BFX2 U22982 ( .A(n17727), .Z(n38700) );
  HS65_LH_BFX2 U22983 ( .A(n17774), .Z(n38701) );
  HS65_LH_BFX2 U22984 ( .A(n17695), .Z(n38702) );
  HS65_LH_BFX2 U22985 ( .A(n38704), .Z(n38703) );
  HS65_LH_BFX2 U22986 ( .A(n17708), .Z(n38704) );
  HS65_LH_IVX2 U22987 ( .A(n40162), .Z(n38705) );
  HS65_LH_IVX2 U22988 ( .A(n38705), .Z(n38706) );
  HS65_LH_BFX2 U22989 ( .A(n38709), .Z(n38707) );
  HS65_LH_IVX2 U22990 ( .A(n38710), .Z(n38708) );
  HS65_LH_IVX2 U22991 ( .A(n38708), .Z(n38709) );
  HS65_LH_BFX2 U22992 ( .A(n17729), .Z(n38710) );
  HS65_LH_BFX2 U22993 ( .A(n38712), .Z(n38711) );
  HS65_LH_BFX2 U22994 ( .A(n38713), .Z(n38712) );
  HS65_LH_BFX2 U22995 ( .A(n17700), .Z(n38713) );
  HS65_LH_BFX2 U22996 ( .A(n38715), .Z(n38714) );
  HS65_LH_BFX2 U22997 ( .A(n38716), .Z(n38715) );
  HS65_LH_BFX2 U22998 ( .A(n17699), .Z(n38716) );
  HS65_LH_BFX2 U22999 ( .A(n38718), .Z(n38717) );
  HS65_LH_BFX2 U23000 ( .A(n38719), .Z(n38718) );
  HS65_LH_BFX2 U23001 ( .A(n17697), .Z(n38719) );
  HS65_LH_BFX2 U23002 ( .A(n38722), .Z(n38720) );
  HS65_LH_IVX2 U23003 ( .A(n38723), .Z(n38721) );
  HS65_LH_IVX2 U23004 ( .A(n38721), .Z(n38722) );
  HS65_LH_BFX2 U23005 ( .A(n38724), .Z(n38723) );
  HS65_LH_BFX2 U23006 ( .A(n38725), .Z(n38724) );
  HS65_LH_BFX2 U23007 ( .A(n38726), .Z(n38725) );
  HS65_LH_BFX2 U23008 ( .A(n38727), .Z(n38726) );
  HS65_LH_BFX2 U23009 ( .A(n38728), .Z(n38727) );
  HS65_LH_BFX2 U23010 ( .A(n38729), .Z(n38728) );
  HS65_LH_BFX2 U23011 ( .A(n38730), .Z(n38729) );
  HS65_LH_BFX2 U23012 ( .A(n38731), .Z(n38730) );
  HS65_LH_BFX2 U23013 ( .A(n38732), .Z(n38731) );
  HS65_LH_BFX2 U23014 ( .A(n38733), .Z(n38732) );
  HS65_LH_BFX2 U23015 ( .A(n17706), .Z(n38733) );
  HS65_LH_IVX2 U23016 ( .A(n38780), .Z(n38734) );
  HS65_LH_IVX2 U23017 ( .A(n38734), .Z(n38735) );
  HS65_LH_BFX2 U23018 ( .A(n30321), .Z(n38736) );
  HS65_LH_IVX2 U23019 ( .A(n38784), .Z(n38737) );
  HS65_LH_IVX2 U23020 ( .A(n38737), .Z(n38738) );
  HS65_LH_BFX2 U23021 ( .A(n29897), .Z(n38739) );
  HS65_LH_BFX2 U23022 ( .A(n38785), .Z(n38740) );
  HS65_LH_IVX2 U23023 ( .A(n38790), .Z(n38741) );
  HS65_LH_IVX2 U23024 ( .A(n38741), .Z(n38742) );
  HS65_LH_BFX2 U23025 ( .A(n38786), .Z(n38743) );
  HS65_LH_IVX2 U23026 ( .A(n38793), .Z(n38744) );
  HS65_LH_IVX2 U23027 ( .A(n38744), .Z(n38745) );
  HS65_LH_BFX2 U23028 ( .A(n30234), .Z(n38746) );
  HS65_LH_BFX2 U23029 ( .A(n38788), .Z(n38747) );
  HS65_LH_BFX2 U23030 ( .A(n38791), .Z(n38748) );
  HS65_LH_BFX2 U23031 ( .A(n38796), .Z(n38749) );
  HS65_LH_BFX2 U23032 ( .A(n38795), .Z(n38750) );
  HS65_LH_BFX2 U23033 ( .A(n29931), .Z(n38751) );
  HS65_LH_BFX2 U23034 ( .A(n30368), .Z(n38752) );
  HS65_LH_BFX2 U23035 ( .A(n38803), .Z(n38753) );
  HS65_LH_BFX2 U23036 ( .A(n38804), .Z(n38754) );
  HS65_LH_BFX2 U23037 ( .A(n39293), .Z(n38755) );
  HS65_LH_BFX2 U23038 ( .A(n38805), .Z(n38756) );
  HS65_LH_IVX2 U23039 ( .A(n38811), .Z(n38757) );
  HS65_LH_IVX2 U23040 ( .A(n38757), .Z(n38758) );
  HS65_LH_IVX2 U23041 ( .A(n38814), .Z(n38759) );
  HS65_LH_IVX2 U23042 ( .A(n38759), .Z(n38760) );
  HS65_LH_BFX2 U23043 ( .A(n29950), .Z(n38761) );
  HS65_LH_BFX2 U23044 ( .A(n30198), .Z(n38762) );
  HS65_LH_BFX2 U23045 ( .A(n30122), .Z(n38763) );
  HS65_LH_IVX2 U23046 ( .A(n38764), .Z(n38765) );
  HS65_LH_BFX2 U23047 ( .A(n29875), .Z(n38766) );
  HS65_LH_BFX2 U23048 ( .A(n38817), .Z(n38767) );
  HS65_LH_BFX2 U23049 ( .A(n30002), .Z(n38768) );
  HS65_LH_BFX2 U23050 ( .A(n30518), .Z(n38769) );
  HS65_LH_BFX2 U23051 ( .A(n38819), .Z(n38770) );
  HS65_LH_BFX2 U23052 ( .A(n38820), .Z(n38771) );
  HS65_LH_BFX2 U23053 ( .A(n38821), .Z(n38772) );
  HS65_LH_BFX2 U23054 ( .A(n38822), .Z(n38773) );
  HS65_LH_BFX2 U23055 ( .A(n38736), .Z(n38774) );
  HS65_LH_BFX2 U23056 ( .A(n38823), .Z(n38775) );
  HS65_LH_IVX2 U23057 ( .A(n38769), .Z(n38776) );
  HS65_LH_IVX2 U23058 ( .A(n38776), .Z(n38777) );
  HS65_LH_BFX2 U23059 ( .A(n38739), .Z(n38778) );
  HS65_LH_IVX2 U23060 ( .A(n38828), .Z(n38779) );
  HS65_LH_IVX2 U23061 ( .A(n38779), .Z(n38780) );
  HS65_LH_IVX2 U23062 ( .A(n38774), .Z(n38781) );
  HS65_LH_IVX2 U23063 ( .A(n38781), .Z(n38782) );
  HS65_LH_IVX2 U23064 ( .A(n38830), .Z(n38783) );
  HS65_LH_IVX2 U23065 ( .A(n38783), .Z(n38784) );
  HS65_LH_BFX2 U23066 ( .A(n38825), .Z(n38785) );
  HS65_LH_BFX2 U23067 ( .A(n38826), .Z(n38786) );
  HS65_LH_BFX2 U23068 ( .A(n38746), .Z(n38787) );
  HS65_LH_BFX2 U23069 ( .A(n38832), .Z(n38788) );
  HS65_LH_IVX2 U23070 ( .A(n38871), .Z(n38789) );
  HS65_LH_IVX2 U23071 ( .A(n38789), .Z(n38790) );
  HS65_LH_BFX2 U23072 ( .A(n38833), .Z(n38791) );
  HS65_LH_IVX2 U23073 ( .A(n38838), .Z(n38792) );
  HS65_LH_IVX2 U23074 ( .A(n38792), .Z(n38793) );
  HS65_LH_BFX2 U23075 ( .A(n30022), .Z(n38794) );
  HS65_LH_BFX2 U23076 ( .A(n17670), .Z(n38795) );
  HS65_LH_BFX2 U23077 ( .A(n38835), .Z(n38796) );
  HS65_LH_BFX2 U23078 ( .A(n30087), .Z(n38797) );
  HS65_LH_BFX2 U23079 ( .A(n38839), .Z(n38798) );
  HS65_LH_BFX2 U23080 ( .A(n38840), .Z(n38799) );
  HS65_LH_BFX2 U23081 ( .A(n38841), .Z(n38800) );
  HS65_LH_BFX2 U23082 ( .A(n38751), .Z(n38801) );
  HS65_LH_BFX2 U23083 ( .A(n38752), .Z(n38802) );
  HS65_LH_BFX2 U23084 ( .A(n38844), .Z(n38803) );
  HS65_LH_BFX2 U23085 ( .A(n38845), .Z(n38804) );
  HS65_LH_BFX2 U23086 ( .A(n38846), .Z(n38805) );
  HS65_LH_BFX2 U23087 ( .A(n38847), .Z(n38806) );
  HS65_LH_BFX2 U23088 ( .A(n38761), .Z(n38807) );
  HS65_LH_BFX2 U23089 ( .A(n38849), .Z(n38808) );
  HS65_LH_BFX2 U23090 ( .A(n38762), .Z(n38809) );
  HS65_LH_IVX2 U23091 ( .A(n38853), .Z(n38810) );
  HS65_LH_IVX2 U23092 ( .A(n38810), .Z(n38811) );
  HS65_LH_BFX2 U23093 ( .A(n18070), .Z(n38812) );
  HS65_LH_IVX2 U23094 ( .A(n38856), .Z(n38813) );
  HS65_LH_IVX2 U23095 ( .A(n38813), .Z(n38814) );
  HS65_LH_BFX2 U23096 ( .A(n38763), .Z(n38815) );
  HS65_LH_BFX2 U23097 ( .A(n38766), .Z(n38816) );
  HS65_LH_BFX2 U23098 ( .A(n38857), .Z(n38817) );
  HS65_LH_BFX2 U23099 ( .A(n38768), .Z(n38818) );
  HS65_LH_BFX2 U23100 ( .A(n38859), .Z(n38819) );
  HS65_LH_BFX2 U23101 ( .A(n38860), .Z(n38820) );
  HS65_LH_BFX2 U23102 ( .A(n38861), .Z(n38821) );
  HS65_LH_BFX2 U23103 ( .A(n38862), .Z(n38822) );
  HS65_LH_BFX2 U23104 ( .A(n38863), .Z(n38823) );
  HS65_LH_BFX2 U23105 ( .A(n38778), .Z(n38824) );
  HS65_LH_BFX2 U23106 ( .A(n38865), .Z(n38825) );
  HS65_LH_BFX2 U23107 ( .A(n38866), .Z(n38826) );
  HS65_LH_IVX2 U23108 ( .A(n38875), .Z(n38827) );
  HS65_LH_IVX2 U23109 ( .A(n38827), .Z(n38828) );
  HS65_LH_IVX2 U23110 ( .A(n38878), .Z(n38829) );
  HS65_LH_IVX2 U23111 ( .A(n38829), .Z(n38830) );
  HS65_LH_BFX2 U23112 ( .A(n38787), .Z(n38831) );
  HS65_LH_BFX2 U23113 ( .A(n38870), .Z(n38832) );
  HS65_LH_BFX2 U23114 ( .A(n38872), .Z(n38833) );
  HS65_LH_BFX2 U23115 ( .A(n38794), .Z(n38834) );
  HS65_LH_BFX2 U23116 ( .A(n38876), .Z(n38835) );
  HS65_LH_BFX2 U23117 ( .A(n38797), .Z(n38836) );
  HS65_LH_IVX2 U23118 ( .A(n38883), .Z(n38837) );
  HS65_LH_IVX2 U23119 ( .A(n38837), .Z(n38838) );
  HS65_LH_BFX2 U23120 ( .A(n38880), .Z(n38839) );
  HS65_LH_BFX2 U23121 ( .A(n38881), .Z(n38840) );
  HS65_LH_BFX2 U23122 ( .A(n38884), .Z(n38841) );
  HS65_LH_BFX2 U23123 ( .A(n38801), .Z(n38842) );
  HS65_LH_BFX2 U23124 ( .A(n38802), .Z(n38843) );
  HS65_LH_BFX2 U23125 ( .A(n38887), .Z(n38844) );
  HS65_LH_BFX2 U23126 ( .A(n38888), .Z(n38845) );
  HS65_LH_BFX2 U23127 ( .A(n38889), .Z(n38846) );
  HS65_LH_BFX2 U23128 ( .A(n38890), .Z(n38847) );
  HS65_LH_BFX2 U23129 ( .A(n38807), .Z(n38848) );
  HS65_LH_BFX2 U23130 ( .A(n38893), .Z(n38849) );
  HS65_LH_BFX2 U23131 ( .A(n38809), .Z(n38850) );
  HS65_LH_BFX2 U23132 ( .A(n38815), .Z(n38851) );
  HS65_LH_IVX2 U23133 ( .A(n38905), .Z(n38852) );
  HS65_LH_IVX2 U23134 ( .A(n38852), .Z(n38853) );
  HS65_LH_BFX2 U23135 ( .A(n38816), .Z(n38854) );
  HS65_LH_IVX2 U23136 ( .A(n38907), .Z(n38855) );
  HS65_LH_IVX2 U23137 ( .A(n38855), .Z(n38856) );
  HS65_LH_BFX2 U23138 ( .A(n38902), .Z(n38857) );
  HS65_LH_BFX2 U23139 ( .A(n38818), .Z(n38858) );
  HS65_LH_BFX2 U23140 ( .A(n38909), .Z(n38859) );
  HS65_LH_BFX2 U23141 ( .A(n38908), .Z(n38860) );
  HS65_LH_BFX2 U23142 ( .A(n38910), .Z(n38861) );
  HS65_LH_BFX2 U23143 ( .A(n38911), .Z(n38862) );
  HS65_LH_BFX2 U23144 ( .A(n38912), .Z(n38863) );
  HS65_LH_BFX2 U23145 ( .A(n38824), .Z(n38864) );
  HS65_LH_BFX2 U23146 ( .A(n38913), .Z(n38865) );
  HS65_LH_BFX2 U23147 ( .A(n38914), .Z(n38866) );
  HS65_LH_IVX2 U23148 ( .A(n39026), .Z(n38867) );
  HS65_LH_IVX2 U23149 ( .A(n38867), .Z(n38868) );
  HS65_LH_BFX2 U23150 ( .A(n38831), .Z(n38869) );
  HS65_LH_BFX2 U23151 ( .A(n38916), .Z(n38870) );
  HS65_LH_BFX2 U23152 ( .A(n38917), .Z(n38871) );
  HS65_LH_BFX2 U23153 ( .A(n38918), .Z(n38872) );
  HS65_LH_BFX2 U23154 ( .A(n38834), .Z(n38873) );
  HS65_LH_IVX2 U23155 ( .A(n38923), .Z(n38874) );
  HS65_LH_IVX2 U23156 ( .A(n38874), .Z(n38875) );
  HS65_LH_BFX2 U23157 ( .A(n38920), .Z(n38876) );
  HS65_LH_IVX2 U23158 ( .A(n38927), .Z(n38877) );
  HS65_LH_IVX2 U23159 ( .A(n38877), .Z(n38878) );
  HS65_LH_BFX2 U23160 ( .A(n38836), .Z(n38879) );
  HS65_LH_BFX2 U23161 ( .A(n38924), .Z(n38880) );
  HS65_LH_BFX2 U23162 ( .A(n38925), .Z(n38881) );
  HS65_LH_IVX2 U23163 ( .A(n38882), .Z(n38883) );
  HS65_LH_BFX2 U23164 ( .A(n38928), .Z(n38884) );
  HS65_LH_BFX2 U23165 ( .A(n38842), .Z(n38885) );
  HS65_LH_BFX2 U23166 ( .A(n38843), .Z(n38886) );
  HS65_LH_BFX2 U23167 ( .A(n38930), .Z(n38887) );
  HS65_LH_BFX2 U23168 ( .A(n38931), .Z(n38888) );
  HS65_LH_BFX2 U23169 ( .A(n38932), .Z(n38889) );
  HS65_LH_BFX2 U23170 ( .A(n38933), .Z(n38890) );
  HS65_LH_BFX2 U23171 ( .A(n38850), .Z(n38891) );
  HS65_LH_BFX2 U23172 ( .A(n38848), .Z(n38892) );
  HS65_LH_BFX2 U23173 ( .A(n38934), .Z(n38893) );
  HS65_LH_IVX2 U23174 ( .A(n38886), .Z(n38894) );
  HS65_LH_IVX2 U23175 ( .A(n38894), .Z(n38895) );
  HS65_LH_IVX2 U23176 ( .A(n38974), .Z(n38896) );
  HS65_LH_IVX2 U23177 ( .A(n38896), .Z(n38897) );
  HS65_LH_IVX2 U23178 ( .A(n38891), .Z(n38898) );
  HS65_LH_IVX2 U23179 ( .A(n38898), .Z(n38899) );
  HS65_LH_BFX2 U23180 ( .A(n38851), .Z(n38900) );
  HS65_LH_BFX2 U23181 ( .A(n38854), .Z(n38901) );
  HS65_LH_BFX2 U23182 ( .A(n38937), .Z(n38902) );
  HS65_LH_BFX2 U23183 ( .A(n38858), .Z(n38903) );
  HS65_LH_IVX2 U23184 ( .A(n38977), .Z(n38904) );
  HS65_LH_IVX2 U23185 ( .A(n38904), .Z(n38905) );
  HS65_LH_IVX2 U23186 ( .A(n38942), .Z(n38906) );
  HS65_LH_IVX2 U23187 ( .A(n38906), .Z(n38907) );
  HS65_LH_BFX2 U23188 ( .A(n17666), .Z(n38908) );
  HS65_LH_BFX2 U23189 ( .A(n38939), .Z(n38909) );
  HS65_LH_BFX2 U23190 ( .A(n38940), .Z(n38910) );
  HS65_LH_BFX2 U23191 ( .A(n38943), .Z(n38911) );
  HS65_LH_BFX2 U23192 ( .A(n38944), .Z(n38912) );
  HS65_LH_BFX2 U23193 ( .A(n38945), .Z(n38913) );
  HS65_LH_BFX2 U23194 ( .A(n38946), .Z(n38914) );
  HS65_LH_BFX2 U23195 ( .A(n38869), .Z(n38915) );
  HS65_LH_BFX2 U23196 ( .A(n38949), .Z(n38916) );
  HS65_LH_BFX2 U23197 ( .A(n18067), .Z(n38917) );
  HS65_LH_BFX2 U23198 ( .A(n38950), .Z(n38918) );
  HS65_LH_BFX2 U23199 ( .A(n38873), .Z(n38919) );
  HS65_LH_BFX2 U23200 ( .A(n38952), .Z(n38920) );
  HS65_LH_BFX2 U23201 ( .A(n38879), .Z(n38921) );
  HS65_LH_IVX2 U23202 ( .A(n38958), .Z(n38922) );
  HS65_LH_IVX2 U23203 ( .A(n38922), .Z(n38923) );
  HS65_LH_BFX2 U23204 ( .A(n18065), .Z(n38924) );
  HS65_LH_BFX2 U23205 ( .A(n38956), .Z(n38925) );
  HS65_LH_IVX2 U23206 ( .A(n38960), .Z(n38926) );
  HS65_LH_IVX2 U23207 ( .A(n38926), .Z(n38927) );
  HS65_LH_BFX2 U23208 ( .A(n38961), .Z(n38928) );
  HS65_LH_BFX2 U23209 ( .A(n38885), .Z(n38929) );
  HS65_LH_BFX2 U23210 ( .A(n38963), .Z(n38930) );
  HS65_LH_BFX2 U23211 ( .A(n38964), .Z(n38931) );
  HS65_LH_BFX2 U23212 ( .A(n38965), .Z(n38932) );
  HS65_LH_BFX2 U23213 ( .A(n38968), .Z(n38933) );
  HS65_LH_BFX2 U23214 ( .A(n38969), .Z(n38934) );
  HS65_LH_BFX2 U23215 ( .A(n38900), .Z(n38935) );
  HS65_LH_BFX2 U23216 ( .A(n38901), .Z(n38936) );
  HS65_LH_BFX2 U23217 ( .A(n38975), .Z(n38937) );
  HS65_LH_BFX2 U23218 ( .A(n38903), .Z(n38938) );
  HS65_LH_BFX2 U23219 ( .A(n38978), .Z(n38939) );
  HS65_LH_BFX2 U23220 ( .A(n38979), .Z(n38940) );
  HS65_LH_IVX2 U23221 ( .A(n38983), .Z(n38941) );
  HS65_LH_IVX2 U23222 ( .A(n38941), .Z(n38942) );
  HS65_LH_BFX2 U23223 ( .A(n38980), .Z(n38943) );
  HS65_LH_BFX2 U23224 ( .A(n38981), .Z(n38944) );
  HS65_LH_BFX2 U23225 ( .A(n38984), .Z(n38945) );
  HS65_LH_BFX2 U23226 ( .A(n38985), .Z(n38946) );
  HS65_LH_BFX2 U23227 ( .A(n38864), .Z(n38947) );
  HS65_LH_BFX2 U23228 ( .A(n38915), .Z(n38948) );
  HS65_LH_BFX2 U23229 ( .A(n38990), .Z(n38949) );
  HS65_LH_BFX2 U23231 ( .A(n38991), .Z(n38950) );
  HS65_LH_BFX2 U23232 ( .A(n38919), .Z(n38951) );
  HS65_LH_BFX2 U23233 ( .A(n38992), .Z(n38952) );
  HS65_LH_BFX2 U23234 ( .A(n38921), .Z(n38953) );
  HS65_LH_IVX2 U23235 ( .A(n39057), .Z(n38954) );
  HS65_LH_IVX2 U23236 ( .A(n38954), .Z(n38955) );
  HS65_LH_BFX2 U23237 ( .A(n38996), .Z(n38956) );
  HS65_LH_IVX2 U23238 ( .A(n39001), .Z(n38957) );
  HS65_LH_IVX2 U23239 ( .A(n38957), .Z(n38958) );
  HS65_LH_IVX2 U23240 ( .A(n39003), .Z(n38959) );
  HS65_LH_IVX2 U23241 ( .A(n38959), .Z(n38960) );
  HS65_LH_BFX2 U23242 ( .A(n38999), .Z(n38961) );
  HS65_LH_BFX2 U23243 ( .A(n38929), .Z(n38962) );
  HS65_LH_BFX2 U23245 ( .A(n39004), .Z(n38963) );
  HS65_LH_BFX2 U23246 ( .A(n39005), .Z(n38964) );
  HS65_LH_BFX2 U23247 ( .A(n39006), .Z(n38965) );
  HS65_LH_IVX2 U23248 ( .A(n39136), .Z(n38966) );
  HS65_LH_IVX2 U23249 ( .A(n38966), .Z(n38967) );
  HS65_LH_BFX2 U23250 ( .A(n39007), .Z(n38968) );
  HS65_LH_BFX2 U23251 ( .A(n39008), .Z(n38969) );
  HS65_LH_BFX2 U23252 ( .A(n38892), .Z(n38970) );
  HS65_LH_BFX2 U23253 ( .A(n38935), .Z(n38971) );
  HS65_LH_BFX2 U23254 ( .A(n38936), .Z(n38972) );
  HS65_LH_IVX2 U23255 ( .A(n39014), .Z(n38973) );
  HS65_LH_IVX2 U23256 ( .A(n38973), .Z(n38974) );
  HS65_LH_BFX2 U23257 ( .A(n39011), .Z(n38975) );
  HS65_LH_BFX2 U23258 ( .A(n38938), .Z(n38976) );
  HS65_LH_BFX2 U23259 ( .A(n39292), .Z(n38977) );
  HS65_LH_BFX2 U23260 ( .A(n39015), .Z(n38978) );
  HS65_LH_BFX2 U23261 ( .A(n39016), .Z(n38979) );
  HS65_LH_BFX2 U23262 ( .A(n39019), .Z(n38980) );
  HS65_LH_BFX2 U23263 ( .A(n39020), .Z(n38981) );
  HS65_LH_IVX2 U23265 ( .A(n38982), .Z(n38983) );
  HS65_LH_BFX2 U23266 ( .A(n38989), .Z(n38984) );
  HS65_LH_BFX2 U23267 ( .A(n39021), .Z(n38985) );
  HS65_LH_BFX2 U23268 ( .A(n38947), .Z(n38986) );
  HS65_LH_BFX2 U23269 ( .A(n38948), .Z(n38987) );
  HS65_LH_IVX2 U23270 ( .A(n39029), .Z(n38988) );
  HS65_LH_IVX2 U23271 ( .A(n38988), .Z(n38989) );
  HS65_LH_BFX2 U23272 ( .A(n39023), .Z(n38990) );
  HS65_LH_BFX2 U23273 ( .A(n39024), .Z(n38991) );
  HS65_LH_BFX2 U23274 ( .A(n39027), .Z(n38992) );
  HS65_LH_BFX2 U23275 ( .A(n38953), .Z(n38993) );
  HS65_LH_IVX2 U23276 ( .A(n38987), .Z(n38994) );
  HS65_LH_IVX2 U23277 ( .A(n38994), .Z(n38995) );
  HS65_LH_BFX2 U23278 ( .A(n39031), .Z(n38996) );
  HS65_LH_IVX2 U23279 ( .A(n38993), .Z(n38997) );
  HS65_LH_IVX2 U23280 ( .A(n38997), .Z(n38998) );
  HS65_LH_BFX2 U23281 ( .A(n39032), .Z(n38999) );
  HS65_LH_IVX2 U23282 ( .A(n39059), .Z(n39000) );
  HS65_LH_IVX2 U23284 ( .A(n39000), .Z(n39001) );
  HS65_LH_IVX2 U23285 ( .A(n39037), .Z(n39002) );
  HS65_LH_IVX2 U23286 ( .A(n39002), .Z(n39003) );
  HS65_LH_BFX2 U23287 ( .A(n17662), .Z(n39004) );
  HS65_LH_BFX2 U23288 ( .A(n39033), .Z(n39005) );
  HS65_LH_BFX2 U23289 ( .A(n39034), .Z(n39006) );
  HS65_LH_BFX2 U23290 ( .A(n39038), .Z(n39007) );
  HS65_LH_BFX2 U23291 ( .A(n39039), .Z(n39008) );
  HS65_LH_BFX2 U23292 ( .A(n38971), .Z(n39009) );
  HS65_LH_BFX2 U23293 ( .A(n38972), .Z(n39010) );
  HS65_LH_BFX2 U23294 ( .A(n39044), .Z(n39011) );
  HS65_LH_BFX2 U23295 ( .A(n38976), .Z(n39012) );
  HS65_LH_IVX2 U23296 ( .A(n39120), .Z(n39013) );
  HS65_LH_IVX2 U23297 ( .A(n39013), .Z(n39014) );
  HS65_LH_BFX2 U23298 ( .A(n39045), .Z(n39015) );
  HS65_LH_BFX2 U23299 ( .A(n39046), .Z(n39016) );
  HS65_LH_IVX2 U23301 ( .A(n39077), .Z(n39017) );
  HS65_LH_IVX2 U23302 ( .A(n39017), .Z(n39018) );
  HS65_LH_BFX2 U23303 ( .A(n18060), .Z(n39019) );
  HS65_LH_BFX2 U23304 ( .A(n39047), .Z(n39020) );
  HS65_LH_BFX2 U23305 ( .A(n39048), .Z(n39021) );
  HS65_LH_BFX2 U23306 ( .A(n38986), .Z(n39022) );
  HS65_LH_BFX2 U23307 ( .A(n39049), .Z(n39023) );
  HS65_LH_BFX2 U23308 ( .A(n39050), .Z(n39024) );
  HS65_LH_IVX2 U23309 ( .A(n39176), .Z(n39025) );
  HS65_LH_IVX2 U23310 ( .A(n39025), .Z(n39026) );
  HS65_LH_BFX2 U23311 ( .A(n39051), .Z(n39027) );
  HS65_LH_IVX2 U23312 ( .A(n39055), .Z(n39028) );
  HS65_LH_IVX2 U23313 ( .A(n39028), .Z(n39029) );
  HS65_LH_BFX2 U23314 ( .A(n38951), .Z(n39030) );
  HS65_LH_BFX2 U23315 ( .A(n39053), .Z(n39031) );
  HS65_LH_BFX2 U23316 ( .A(n39058), .Z(n39032) );
  HS65_LH_BFX2 U23317 ( .A(n39060), .Z(n39033) );
  HS65_LH_BFX2 U23319 ( .A(n39061), .Z(n39034) );
  HS65_LH_BFX2 U23320 ( .A(n38962), .Z(n39035) );
  HS65_LH_IVX2 U23321 ( .A(n39066), .Z(n39036) );
  HS65_LH_IVX2 U23322 ( .A(n39036), .Z(n39037) );
  HS65_LH_BFX2 U23323 ( .A(n39063), .Z(n39038) );
  HS65_LH_BFX2 U23324 ( .A(n39064), .Z(n39039) );
  HS65_LH_BFX2 U23325 ( .A(n39009), .Z(n39040) );
  HS65_LH_BFX2 U23326 ( .A(n39010), .Z(n39041) );
  HS65_LH_IVX2 U23327 ( .A(n39074), .Z(n39042) );
  HS65_LH_IVX2 U23328 ( .A(n39042), .Z(n39043) );
  HS65_LH_BFX2 U23329 ( .A(n39068), .Z(n39044) );
  HS65_LH_BFX2 U23330 ( .A(n39070), .Z(n39045) );
  HS65_LH_BFX2 U23331 ( .A(n39072), .Z(n39046) );
  HS65_LH_BFX2 U23332 ( .A(n39075), .Z(n39047) );
  HS65_LH_BFX2 U23333 ( .A(n39078), .Z(n39048) );
  HS65_LH_BFX2 U23334 ( .A(n39079), .Z(n39049) );
  HS65_LH_BFX2 U23335 ( .A(n39080), .Z(n39050) );
  HS65_LH_BFX2 U23337 ( .A(n39082), .Z(n39051) );
  HS65_LH_BFX2 U23338 ( .A(n39030), .Z(n39052) );
  HS65_LH_BFX2 U23339 ( .A(n39083), .Z(n39053) );
  HS65_LH_IVX2 U23340 ( .A(n39085), .Z(n39054) );
  HS65_LH_IVX2 U23341 ( .A(n39054), .Z(n39055) );
  HS65_LH_IVX2 U23342 ( .A(n39087), .Z(n39056) );
  HS65_LH_IVX2 U23343 ( .A(n39056), .Z(n39057) );
  HS65_LH_BFX2 U23344 ( .A(n39088), .Z(n39058) );
  HS65_LH_BFX2 U23345 ( .A(n39291), .Z(n39059) );
  HS65_LH_BFX2 U23346 ( .A(n39089), .Z(n39060) );
  HS65_LH_BFX2 U23347 ( .A(n39090), .Z(n39061) );
  HS65_LH_BFX2 U23348 ( .A(n39035), .Z(n39062) );
  HS65_LH_BFX2 U23349 ( .A(n39092), .Z(n39063) );
  HS65_LH_BFX2 U23350 ( .A(n39093), .Z(n39064) );
  HS65_LH_IVX2 U23351 ( .A(n39065), .Z(n39066) );
  HS65_LH_BFX2 U23352 ( .A(n39041), .Z(n39067) );
  HS65_LH_BFX2 U23353 ( .A(n39095), .Z(n39068) );
  HS65_LH_BFX2 U23354 ( .A(n38970), .Z(n39069) );
  HS65_LH_BFX2 U23355 ( .A(n39097), .Z(n39070) );
  HS65_LH_BFX2 U23356 ( .A(n39012), .Z(n39071) );
  HS65_LH_BFX2 U23358 ( .A(n39098), .Z(n39072) );
  HS65_LH_IVX2 U23359 ( .A(n39040), .Z(n39073) );
  HS65_LH_IVX2 U23360 ( .A(n39073), .Z(n39074) );
  HS65_LH_BFX2 U23361 ( .A(n39099), .Z(n39075) );
  HS65_LH_IVX2 U23362 ( .A(n39071), .Z(n39076) );
  HS65_LH_IVX2 U23363 ( .A(n39076), .Z(n39077) );
  HS65_LH_BFX2 U23364 ( .A(n39100), .Z(n39078) );
  HS65_LH_BFX2 U23365 ( .A(n17658), .Z(n39079) );
  HS65_LH_BFX2 U23366 ( .A(n39101), .Z(n39080) );
  HS65_LH_BFX2 U23367 ( .A(n39022), .Z(n39081) );
  HS65_LH_BFX2 U23368 ( .A(n39103), .Z(n39082) );
  HS65_LH_BFX2 U23369 ( .A(n39104), .Z(n39083) );
  HS65_LH_IVX2 U23370 ( .A(n39107), .Z(n39084) );
  HS65_LH_IVX2 U23371 ( .A(n39084), .Z(n39085) );
  HS65_LH_IVX2 U23372 ( .A(n39133), .Z(n39086) );
  HS65_LH_IVX2 U23373 ( .A(n39086), .Z(n39087) );
  HS65_LH_BFX2 U23374 ( .A(n39105), .Z(n39088) );
  HS65_LH_BFX2 U23376 ( .A(n39108), .Z(n39089) );
  HS65_LH_BFX2 U23377 ( .A(n39109), .Z(n39090) );
  HS65_LH_BFX2 U23378 ( .A(n39062), .Z(n39091) );
  HS65_LH_BFX2 U23379 ( .A(n18055), .Z(n39092) );
  HS65_LH_BFX2 U23380 ( .A(n39111), .Z(n39093) );
  HS65_LH_BFX2 U23381 ( .A(n39067), .Z(n39094) );
  HS65_LH_BFX2 U23382 ( .A(n39113), .Z(n39095) );
  HS65_LH_BFX2 U23383 ( .A(n39069), .Z(n39096) );
  HS65_LH_BFX2 U23384 ( .A(n39117), .Z(n39097) );
  HS65_LH_BFX2 U23385 ( .A(n39118), .Z(n39098) );
  HS65_LH_BFX2 U23386 ( .A(n39121), .Z(n39099) );
  HS65_LH_BFX2 U23387 ( .A(n39122), .Z(n39100) );
  HS65_LH_BFX2 U23388 ( .A(n39123), .Z(n39101) );
  HS65_LH_BFX2 U23389 ( .A(n39081), .Z(n39102) );
  HS65_LH_BFX2 U23390 ( .A(n39125), .Z(n39103) );
  HS65_LH_BFX2 U23391 ( .A(n39126), .Z(n39104) );
  HS65_LH_BFX2 U23392 ( .A(n39128), .Z(n39105) );
  HS65_LH_IVX2 U23394 ( .A(n39153), .Z(n39106) );
  HS65_LH_IVX2 U23395 ( .A(n39106), .Z(n39107) );
  HS65_LH_BFX2 U23396 ( .A(n39129), .Z(n39108) );
  HS65_LH_BFX2 U23397 ( .A(n39131), .Z(n39109) );
  HS65_LH_BFX2 U23398 ( .A(n39091), .Z(n39110) );
  HS65_LH_BFX2 U23399 ( .A(n39134), .Z(n39111) );
  HS65_LH_BFX2 U23400 ( .A(n39094), .Z(n39112) );
  HS65_LH_BFX2 U23401 ( .A(n39137), .Z(n39113) );
  HS65_LH_BFX2 U23402 ( .A(n39096), .Z(n39114) );
  HS65_LH_IVX2 U23403 ( .A(n39202), .Z(n39115) );
  HS65_LH_IVX2 U23404 ( .A(n39115), .Z(n39116) );
  HS65_LH_BFX2 U23405 ( .A(n39138), .Z(n39117) );
  HS65_LH_BFX2 U23406 ( .A(n39139), .Z(n39118) );
  HS65_LH_IVX2 U23407 ( .A(n39142), .Z(n39119) );
  HS65_LH_IVX2 U23408 ( .A(n39119), .Z(n39120) );
  HS65_LH_BFX2 U23409 ( .A(n39140), .Z(n39121) );
  HS65_LH_BFX2 U23410 ( .A(n39143), .Z(n39122) );
  HS65_LH_BFX2 U23412 ( .A(n39144), .Z(n39123) );
  HS65_LH_BFX2 U23413 ( .A(n39102), .Z(n39124) );
  HS65_LH_BFX2 U23414 ( .A(n39146), .Z(n39125) );
  HS65_LH_BFX2 U23415 ( .A(n39147), .Z(n39126) );
  HS65_LH_BFX2 U23416 ( .A(n39052), .Z(n39127) );
  HS65_LH_BFX2 U23417 ( .A(n39148), .Z(n39128) );
  HS65_LH_BFX2 U23418 ( .A(n39150), .Z(n39129) );
  HS65_LH_BFX2 U23419 ( .A(n39110), .Z(n39130) );
  HS65_LH_BFX2 U23420 ( .A(n39151), .Z(n39131) );
  HS65_LH_IVX2 U23421 ( .A(n39127), .Z(n39132) );
  HS65_LH_IVX2 U23422 ( .A(n39132), .Z(n39133) );
  HS65_LH_BFX2 U23423 ( .A(n39154), .Z(n39134) );
  HS65_LH_IVX2 U23424 ( .A(n39130), .Z(n39135) );
  HS65_LH_IVX2 U23425 ( .A(n39135), .Z(n39136) );
  HS65_LH_BFX2 U23426 ( .A(n17722), .Z(n39137) );
  HS65_LH_BFX2 U23427 ( .A(n39156), .Z(n39138) );
  HS65_LH_BFX2 U23429 ( .A(n17656), .Z(n39139) );
  HS65_LH_BFX2 U23430 ( .A(n39157), .Z(n39140) );
  HS65_LH_IVX2 U23431 ( .A(n39159), .Z(n39141) );
  HS65_LH_IVX2 U23432 ( .A(n39141), .Z(n39142) );
  HS65_LH_BFX2 U23433 ( .A(n39160), .Z(n39143) );
  HS65_LH_BFX2 U23434 ( .A(n39161), .Z(n39144) );
  HS65_LH_BFX2 U23435 ( .A(n39124), .Z(n39145) );
  HS65_LH_BFX2 U23436 ( .A(n18051), .Z(n39146) );
  HS65_LH_BFX2 U23437 ( .A(n18053), .Z(n39147) );
  HS65_LH_BFX2 U23438 ( .A(n39163), .Z(n39148) );
  HS65_LH_BFX2 U23439 ( .A(n18042), .Z(n39149) );
  HS65_LH_BFX2 U23440 ( .A(n39164), .Z(n39150) );
  HS65_LH_BFX2 U23442 ( .A(n39165), .Z(n39151) );
  HS65_LH_IVX2 U23443 ( .A(n39183), .Z(n39152) );
  HS65_LH_IVX2 U23444 ( .A(n39152), .Z(n39153) );
  HS65_LH_BFX2 U23445 ( .A(n39166), .Z(n39154) );
  HS65_LH_BFX2 U23446 ( .A(n39112), .Z(n39155) );
  HS65_LH_BFX2 U23447 ( .A(n39168), .Z(n39156) );
  HS65_LH_BFX2 U23448 ( .A(n39169), .Z(n39157) );
  HS65_LH_IVX2 U23449 ( .A(n39174), .Z(n39158) );
  HS65_LH_IVX2 U23450 ( .A(n39158), .Z(n39159) );
  HS65_LH_BFX2 U23451 ( .A(n39170), .Z(n39160) );
  HS65_LH_BFX2 U23452 ( .A(n39172), .Z(n39161) );
  HS65_LH_BFX2 U23453 ( .A(n39145), .Z(n39162) );
  HS65_LH_BFX2 U23455 ( .A(n39177), .Z(n39163) );
  HS65_LH_BFX2 U23456 ( .A(n39178), .Z(n39164) );
  HS65_LH_BFX2 U23457 ( .A(n39179), .Z(n39165) );
  HS65_LH_BFX2 U23458 ( .A(n39181), .Z(n39166) );
  HS65_LH_BFX2 U23459 ( .A(n39155), .Z(n39167) );
  HS65_LH_BFX2 U23460 ( .A(n39185), .Z(n39168) );
  HS65_LH_BFX2 U23461 ( .A(n39186), .Z(n39169) );
  HS65_LH_BFX2 U23462 ( .A(n39187), .Z(n39170) );
  HS65_LH_BFX2 U23463 ( .A(n39162), .Z(n39171) );
  HS65_LH_BFX2 U23464 ( .A(n39188), .Z(n39172) );
  HS65_LH_IVX2 U23465 ( .A(n39114), .Z(n39173) );
  HS65_LH_IVX2 U23466 ( .A(n39173), .Z(n39174) );
  HS65_LH_IVX2 U23468 ( .A(n39171), .Z(n39175) );
  HS65_LH_IVX2 U23469 ( .A(n39175), .Z(n39176) );
  HS65_LH_BFX2 U23470 ( .A(n17718), .Z(n39177) );
  HS65_LH_BFX2 U23471 ( .A(n39189), .Z(n39178) );
  HS65_LH_BFX2 U23472 ( .A(n17720), .Z(n39179) );
  HS65_LH_BFX2 U23473 ( .A(n39149), .Z(n39180) );
  HS65_LH_BFX2 U23474 ( .A(n39190), .Z(n39181) );
  HS65_LH_IVX2 U23475 ( .A(n39192), .Z(n39182) );
  HS65_LH_IVX2 U23476 ( .A(n39182), .Z(n39183) );
  HS65_LH_BFX2 U23477 ( .A(n39167), .Z(n39184) );
  HS65_LH_BFX2 U23478 ( .A(n18047), .Z(n39185) );
  HS65_LH_BFX2 U23479 ( .A(n18049), .Z(n39186) );
  HS65_LH_BFX2 U23480 ( .A(n39194), .Z(n39187) );
  HS65_LH_BFX2 U23481 ( .A(n39195), .Z(n39188) );
  HS65_LH_BFX2 U23482 ( .A(n39196), .Z(n39189) );
  HS65_LH_BFX2 U23483 ( .A(n39197), .Z(n39190) );
  HS65_LH_IVX2 U23484 ( .A(n39200), .Z(n39191) );
  HS65_LH_IVX2 U23485 ( .A(n39191), .Z(n39192) );
  HS65_LH_BFX2 U23486 ( .A(n39184), .Z(n39193) );
  HS65_LH_BFX2 U23487 ( .A(n39203), .Z(n39194) );
  HS65_LH_BFX2 U23488 ( .A(n39204), .Z(n39195) );
  HS65_LH_BFX2 U23489 ( .A(n39205), .Z(n39196) );
  HS65_LH_BFX2 U23490 ( .A(n39206), .Z(n39197) );
  HS65_LH_BFX2 U23491 ( .A(n39193), .Z(n39198) );
  HS65_LH_IVX2 U23492 ( .A(n39180), .Z(n39199) );
  HS65_LH_IVX2 U23493 ( .A(n39199), .Z(n39200) );
  HS65_LH_IVX2 U23494 ( .A(n39198), .Z(n39201) );
  HS65_LH_IVX2 U23495 ( .A(n39201), .Z(n39202) );
  HS65_LH_BFX2 U23496 ( .A(n17714), .Z(n39203) );
  HS65_LH_BFX2 U23497 ( .A(n17716), .Z(n39204) );
  HS65_LH_BFX2 U23498 ( .A(n18043), .Z(n39205) );
  HS65_LH_BFX2 U23499 ( .A(n18045), .Z(n39206) );
  HS65_LH_BFX2 U23500 ( .A(n39210), .Z(n39207) );
  HS65_LH_BFX2 U23501 ( .A(n18032), .Z(n39208) );
  HS65_LH_BFX2 U23502 ( .A(n39212), .Z(n39209) );
  HS65_LH_BFX2 U23503 ( .A(n39213), .Z(n39210) );
  HS65_LH_BFX2 U23504 ( .A(n39208), .Z(n39211) );
  HS65_LH_BFX2 U23505 ( .A(n39215), .Z(n39212) );
  HS65_LH_BFX2 U23506 ( .A(n39216), .Z(n39213) );
  HS65_LH_BFX2 U23507 ( .A(n39211), .Z(n39214) );
  HS65_LH_BFX2 U23508 ( .A(n39218), .Z(n39215) );
  HS65_LH_BFX2 U23509 ( .A(n39219), .Z(n39216) );
  HS65_LH_BFX2 U23510 ( .A(n39214), .Z(n39217) );
  HS65_LH_BFX2 U23511 ( .A(n39221), .Z(n39218) );
  HS65_LH_BFX2 U23512 ( .A(n39222), .Z(n39219) );
  HS65_LH_BFX2 U23513 ( .A(n39217), .Z(n39220) );
  HS65_LH_BFX2 U23514 ( .A(n39224), .Z(n39221) );
  HS65_LH_BFX2 U23515 ( .A(n39225), .Z(n39222) );
  HS65_LH_BFX2 U23516 ( .A(n39220), .Z(n39223) );
  HS65_LH_BFX2 U23517 ( .A(n39227), .Z(n39224) );
  HS65_LH_BFX2 U23518 ( .A(n39228), .Z(n39225) );
  HS65_LH_BFX2 U23519 ( .A(n39223), .Z(n39226) );
  HS65_LH_BFX2 U23520 ( .A(n39230), .Z(n39227) );
  HS65_LH_BFX2 U23521 ( .A(n39231), .Z(n39228) );
  HS65_LH_BFX2 U23522 ( .A(n39226), .Z(n39229) );
  HS65_LH_BFX2 U23523 ( .A(n39233), .Z(n39230) );
  HS65_LH_BFX2 U23524 ( .A(n39234), .Z(n39231) );
  HS65_LH_BFX2 U23525 ( .A(n39229), .Z(n39232) );
  HS65_LH_BFX2 U23526 ( .A(n39236), .Z(n39233) );
  HS65_LH_BFX2 U23527 ( .A(n39237), .Z(n39234) );
  HS65_LH_BFX2 U23528 ( .A(n39232), .Z(n39235) );
  HS65_LH_BFX2 U23529 ( .A(n39239), .Z(n39236) );
  HS65_LH_BFX2 U23530 ( .A(n39240), .Z(n39237) );
  HS65_LH_BFX2 U23531 ( .A(n39235), .Z(n39238) );
  HS65_LH_BFX2 U23532 ( .A(n39242), .Z(n39239) );
  HS65_LH_BFX2 U23533 ( .A(n39243), .Z(n39240) );
  HS65_LH_BFX2 U23534 ( .A(n39238), .Z(n39241) );
  HS65_LH_BFX2 U23535 ( .A(n39245), .Z(n39242) );
  HS65_LH_BFX2 U23536 ( .A(n39246), .Z(n39243) );
  HS65_LH_BFX2 U23537 ( .A(n39241), .Z(n39244) );
  HS65_LH_BFX2 U23538 ( .A(n39248), .Z(n39245) );
  HS65_LH_BFX2 U23539 ( .A(n39249), .Z(n39246) );
  HS65_LH_BFX2 U23540 ( .A(n39244), .Z(n39247) );
  HS65_LH_BFX2 U23541 ( .A(n39251), .Z(n39248) );
  HS65_LH_BFX2 U23542 ( .A(n39252), .Z(n39249) );
  HS65_LH_BFX2 U23543 ( .A(n39247), .Z(n39250) );
  HS65_LH_BFX2 U23544 ( .A(n39254), .Z(n39251) );
  HS65_LH_BFX2 U23545 ( .A(n39255), .Z(n39252) );
  HS65_LH_BFX2 U23546 ( .A(n39250), .Z(n39253) );
  HS65_LH_BFX2 U23547 ( .A(n39257), .Z(n39254) );
  HS65_LH_BFX2 U23548 ( .A(n39258), .Z(n39255) );
  HS65_LH_BFX2 U23549 ( .A(n39253), .Z(n39256) );
  HS65_LH_BFX2 U23550 ( .A(n39260), .Z(n39257) );
  HS65_LH_BFX2 U23551 ( .A(n39261), .Z(n39258) );
  HS65_LH_BFX2 U23552 ( .A(n39256), .Z(n39259) );
  HS65_LH_BFX2 U23553 ( .A(n15466), .Z(n39260) );
  HS65_LH_BFX2 U23554 ( .A(n39264), .Z(n39261) );
  HS65_LH_BFX2 U23555 ( .A(n39259), .Z(n39262) );
  HS65_LH_IVX2 U23556 ( .A(n18033), .Z(n39263) );
  HS65_LH_IVX2 U23557 ( .A(n39263), .Z(n39264) );
  HS65_LH_IVX2 U23558 ( .A(n39262), .Z(n39265) );
  HS65_LH_IVX2 U23559 ( .A(n39265), .Z(n39266) );
  HS65_LH_BFX2 U23560 ( .A(n39297), .Z(n39267) );
  HS65_LH_BFX2 U23561 ( .A(n18027), .Z(n39268) );
  HS65_LH_BFX2 U23562 ( .A(n39299), .Z(n39269) );
  HS65_LH_BFX2 U23563 ( .A(n39271), .Z(n39270) );
  HS65_LH_BFX2 U23564 ( .A(n39272), .Z(n39271) );
  HS65_LH_BFX2 U23565 ( .A(n39273), .Z(n39272) );
  HS65_LH_BFX2 U23566 ( .A(n39274), .Z(n39273) );
  HS65_LH_BFX2 U23567 ( .A(n39275), .Z(n39274) );
  HS65_LH_BFX2 U23568 ( .A(n39276), .Z(n39275) );
  HS65_LH_BFX2 U23569 ( .A(n39277), .Z(n39276) );
  HS65_LH_BFX2 U23570 ( .A(n39278), .Z(n39277) );
  HS65_LH_BFX2 U23571 ( .A(n39279), .Z(n39278) );
  HS65_LH_BFX2 U23572 ( .A(n39280), .Z(n39279) );
  HS65_LH_BFX2 U23573 ( .A(n39281), .Z(n39280) );
  HS65_LH_BFX2 U23574 ( .A(n39282), .Z(n39281) );
  HS65_LH_BFX2 U23575 ( .A(n39283), .Z(n39282) );
  HS65_LH_BFX2 U23576 ( .A(n39284), .Z(n39283) );
  HS65_LH_BFX2 U23577 ( .A(n39285), .Z(n39284) );
  HS65_LH_BFX2 U23578 ( .A(n39286), .Z(n39285) );
  HS65_LH_BFX2 U23579 ( .A(n39287), .Z(n39286) );
  HS65_LH_BFX2 U23580 ( .A(n39288), .Z(n39287) );
  HS65_LH_BFX2 U23581 ( .A(n39289), .Z(n39288) );
  HS65_LH_BFX2 U23582 ( .A(n39290), .Z(n39289) );
  HS65_LH_BFX2 U23583 ( .A(n17738), .Z(n39290) );
  HS65_LH_BFX2 U23584 ( .A(n18056), .Z(n39291) );
  HS65_LH_BFX2 U23585 ( .A(n18062), .Z(n39292) );
  HS65_LH_BFX2 U23586 ( .A(n18072), .Z(n39293) );
  HS65_LH_BFX2 U23587 ( .A(n18077), .Z(n39294) );
  HS65_LH_BFX2 U23588 ( .A(n18086), .Z(n39295) );
  HS65_LH_BFX2 U23590 ( .A(n18085), .Z(n39296) );
  HS65_LH_BFX2 U23591 ( .A(n39300), .Z(n39297) );
  HS65_LH_BFX2 U23593 ( .A(n39268), .Z(n39298) );
  HS65_LH_BFX2 U23594 ( .A(n39302), .Z(n39299) );
  HS65_LH_BFX2 U23595 ( .A(n39303), .Z(n39300) );
  HS65_LH_BFX2 U23596 ( .A(n39298), .Z(n39301) );
  HS65_LH_BFX2 U23597 ( .A(n39305), .Z(n39302) );
  HS65_LH_BFX2 U23598 ( .A(n39306), .Z(n39303) );
  HS65_LH_BFX2 U23599 ( .A(n39301), .Z(n39304) );
  HS65_LH_BFX2 U23600 ( .A(n39308), .Z(n39305) );
  HS65_LH_BFX2 U23601 ( .A(n39309), .Z(n39306) );
  HS65_LH_BFX2 U23602 ( .A(n39304), .Z(n39307) );
  HS65_LH_BFX2 U23603 ( .A(n39311), .Z(n39308) );
  HS65_LH_BFX2 U23604 ( .A(n39312), .Z(n39309) );
  HS65_LH_BFX2 U23605 ( .A(n39307), .Z(n39310) );
  HS65_LH_BFX2 U23606 ( .A(n39314), .Z(n39311) );
  HS65_LH_BFX2 U23607 ( .A(n39315), .Z(n39312) );
  HS65_LH_BFX2 U23608 ( .A(n39310), .Z(n39313) );
  HS65_LH_BFX2 U23609 ( .A(n39317), .Z(n39314) );
  HS65_LH_BFX2 U23610 ( .A(n39318), .Z(n39315) );
  HS65_LH_BFX2 U23611 ( .A(n39313), .Z(n39316) );
  HS65_LH_BFX2 U23612 ( .A(n39320), .Z(n39317) );
  HS65_LH_BFX2 U23613 ( .A(n39321), .Z(n39318) );
  HS65_LH_BFX2 U23614 ( .A(n39316), .Z(n39319) );
  HS65_LH_BFX2 U23615 ( .A(n39323), .Z(n39320) );
  HS65_LH_BFX2 U23616 ( .A(n39324), .Z(n39321) );
  HS65_LH_BFX2 U23617 ( .A(n39319), .Z(n39322) );
  HS65_LH_BFX2 U23618 ( .A(n39326), .Z(n39323) );
  HS65_LH_BFX2 U23619 ( .A(n39327), .Z(n39324) );
  HS65_LH_BFX2 U23620 ( .A(n39322), .Z(n39325) );
  HS65_LH_BFX2 U23621 ( .A(n39329), .Z(n39326) );
  HS65_LH_BFX2 U23622 ( .A(n39330), .Z(n39327) );
  HS65_LH_BFX2 U23623 ( .A(n39325), .Z(n39328) );
  HS65_LH_BFX2 U23624 ( .A(n39332), .Z(n39329) );
  HS65_LH_BFX2 U23625 ( .A(n39333), .Z(n39330) );
  HS65_LH_BFX2 U23626 ( .A(n39328), .Z(n39331) );
  HS65_LH_BFX2 U23627 ( .A(n39335), .Z(n39332) );
  HS65_LH_BFX2 U23628 ( .A(n39336), .Z(n39333) );
  HS65_LH_BFX2 U23629 ( .A(n39331), .Z(n39334) );
  HS65_LH_BFX2 U23630 ( .A(n39338), .Z(n39335) );
  HS65_LH_BFX2 U23631 ( .A(n39339), .Z(n39336) );
  HS65_LH_BFX2 U23632 ( .A(n39334), .Z(n39337) );
  HS65_LH_BFX2 U23633 ( .A(n39341), .Z(n39338) );
  HS65_LH_BFX2 U23634 ( .A(n39342), .Z(n39339) );
  HS65_LH_BFX2 U23635 ( .A(n39337), .Z(n39340) );
  HS65_LH_BFX2 U23636 ( .A(n39344), .Z(n39341) );
  HS65_LH_BFX2 U23637 ( .A(n39345), .Z(n39342) );
  HS65_LH_BFX2 U23638 ( .A(n39340), .Z(n39343) );
  HS65_LH_BFX2 U23639 ( .A(n39347), .Z(n39344) );
  HS65_LH_BFX2 U23640 ( .A(n39348), .Z(n39345) );
  HS65_LH_BFX2 U23641 ( .A(n39343), .Z(n39346) );
  HS65_LH_BFX2 U23642 ( .A(n39354), .Z(n39347) );
  HS65_LH_BFX2 U23643 ( .A(n39351), .Z(n39348) );
  HS65_LH_BFX2 U23644 ( .A(n39346), .Z(n39349) );
  HS65_LH_IVX2 U23645 ( .A(n18028), .Z(n39350) );
  HS65_LH_IVX2 U23646 ( .A(n39350), .Z(n39351) );
  HS65_LH_IVX2 U23647 ( .A(n39349), .Z(n39352) );
  HS65_LH_IVX2 U23648 ( .A(n39352), .Z(n39353) );
  HS65_LH_BFX2 U23649 ( .A(n15469), .Z(n39354) );
  HS65_LH_BFX2 U23650 ( .A(n40503), .Z(n39355) );
  HS65_LH_BFX2 U23651 ( .A(n39357), .Z(n39356) );
  HS65_LH_BFX2 U23652 ( .A(n39358), .Z(n39357) );
  HS65_LH_BFX2 U23653 ( .A(n39359), .Z(n39358) );
  HS65_LH_BFX2 U23654 ( .A(n39360), .Z(n39359) );
  HS65_LH_BFX2 U23655 ( .A(n39361), .Z(n39360) );
  HS65_LH_BFX2 U23656 ( .A(n39362), .Z(n39361) );
  HS65_LH_BFX2 U23657 ( .A(n39363), .Z(n39362) );
  HS65_LH_BFX2 U23658 ( .A(n39364), .Z(n39363) );
  HS65_LH_BFX2 U23659 ( .A(n39365), .Z(n39364) );
  HS65_LH_BFX2 U23660 ( .A(n39366), .Z(n39365) );
  HS65_LH_BFX2 U23661 ( .A(n39367), .Z(n39366) );
  HS65_LH_BFX2 U23662 ( .A(n39368), .Z(n39367) );
  HS65_LH_BFX2 U23663 ( .A(n39369), .Z(n39368) );
  HS65_LH_BFX2 U23664 ( .A(n39370), .Z(n39369) );
  HS65_LH_BFX2 U23665 ( .A(n39371), .Z(n39370) );
  HS65_LH_BFX2 U23666 ( .A(n39372), .Z(n39371) );
  HS65_LH_BFX2 U23667 ( .A(n39373), .Z(n39372) );
  HS65_LH_BFX2 U23668 ( .A(n39374), .Z(n39373) );
  HS65_LH_BFX2 U23669 ( .A(n39375), .Z(n39374) );
  HS65_LH_BFX2 U23670 ( .A(n39376), .Z(n39375) );
  HS65_LH_BFX2 U23671 ( .A(n39377), .Z(n39376) );
  HS65_LH_BFX2 U23672 ( .A(n17795), .Z(n39377) );
  HS65_LH_BFX2 U23673 ( .A(n39379), .Z(n39378) );
  HS65_LH_BFX2 U23674 ( .A(n39380), .Z(n39379) );
  HS65_LH_BFX2 U23675 ( .A(n39381), .Z(n39380) );
  HS65_LH_BFX2 U23676 ( .A(n39382), .Z(n39381) );
  HS65_LH_BFX2 U23677 ( .A(n39383), .Z(n39382) );
  HS65_LH_BFX2 U23678 ( .A(n39384), .Z(n39383) );
  HS65_LH_BFX2 U23679 ( .A(n39385), .Z(n39384) );
  HS65_LH_BFX2 U23680 ( .A(n39386), .Z(n39385) );
  HS65_LH_BFX2 U23681 ( .A(n39387), .Z(n39386) );
  HS65_LH_BFX2 U23682 ( .A(n39388), .Z(n39387) );
  HS65_LH_BFX2 U23683 ( .A(n39389), .Z(n39388) );
  HS65_LH_BFX2 U23684 ( .A(n39390), .Z(n39389) );
  HS65_LH_BFX2 U23685 ( .A(n39391), .Z(n39390) );
  HS65_LH_BFX2 U23686 ( .A(n39392), .Z(n39391) );
  HS65_LH_BFX2 U23687 ( .A(n39393), .Z(n39392) );
  HS65_LH_BFX2 U23688 ( .A(n39394), .Z(n39393) );
  HS65_LH_BFX2 U23689 ( .A(n39395), .Z(n39394) );
  HS65_LH_BFX2 U23690 ( .A(n39396), .Z(n39395) );
  HS65_LH_BFX2 U23691 ( .A(n39397), .Z(n39396) );
  HS65_LH_BFX2 U23692 ( .A(n39398), .Z(n39397) );
  HS65_LH_BFX2 U23693 ( .A(n39399), .Z(n39398) );
  HS65_LH_BFX2 U23694 ( .A(n17794), .Z(n39399) );
  HS65_LH_BFX2 U23695 ( .A(n39401), .Z(n39400) );
  HS65_LH_BFX2 U23696 ( .A(n39402), .Z(n39401) );
  HS65_LH_BFX2 U23697 ( .A(n39403), .Z(n39402) );
  HS65_LH_BFX2 U23698 ( .A(n39404), .Z(n39403) );
  HS65_LH_BFX2 U23699 ( .A(n39405), .Z(n39404) );
  HS65_LH_BFX2 U23700 ( .A(n39406), .Z(n39405) );
  HS65_LH_BFX2 U23701 ( .A(n39407), .Z(n39406) );
  HS65_LH_BFX2 U23702 ( .A(n39408), .Z(n39407) );
  HS65_LH_BFX2 U23703 ( .A(n39409), .Z(n39408) );
  HS65_LH_BFX2 U23704 ( .A(n39410), .Z(n39409) );
  HS65_LH_BFX2 U23705 ( .A(n39411), .Z(n39410) );
  HS65_LH_BFX2 U23706 ( .A(n39412), .Z(n39411) );
  HS65_LH_BFX2 U23707 ( .A(n39413), .Z(n39412) );
  HS65_LH_BFX2 U23708 ( .A(n39414), .Z(n39413) );
  HS65_LH_BFX2 U23709 ( .A(n39415), .Z(n39414) );
  HS65_LH_BFX2 U23710 ( .A(n39416), .Z(n39415) );
  HS65_LH_BFX2 U23711 ( .A(n39417), .Z(n39416) );
  HS65_LH_BFX2 U23712 ( .A(n39418), .Z(n39417) );
  HS65_LH_BFX2 U23713 ( .A(n39419), .Z(n39418) );
  HS65_LH_BFX2 U23714 ( .A(n39420), .Z(n39419) );
  HS65_LH_BFX2 U23715 ( .A(n39421), .Z(n39420) );
  HS65_LH_BFX2 U23716 ( .A(n17801), .Z(n39421) );
  HS65_LH_BFX2 U23717 ( .A(n39423), .Z(n39422) );
  HS65_LH_BFX2 U23718 ( .A(n39424), .Z(n39423) );
  HS65_LH_BFX2 U23719 ( .A(n39425), .Z(n39424) );
  HS65_LH_BFX2 U23720 ( .A(n39426), .Z(n39425) );
  HS65_LH_BFX2 U23721 ( .A(n39427), .Z(n39426) );
  HS65_LH_BFX2 U23722 ( .A(n39428), .Z(n39427) );
  HS65_LH_BFX2 U23723 ( .A(n39429), .Z(n39428) );
  HS65_LH_BFX2 U23724 ( .A(n39430), .Z(n39429) );
  HS65_LH_BFX2 U23725 ( .A(n39431), .Z(n39430) );
  HS65_LH_BFX2 U23726 ( .A(n39432), .Z(n39431) );
  HS65_LH_BFX2 U23727 ( .A(n39433), .Z(n39432) );
  HS65_LH_BFX2 U23728 ( .A(n39434), .Z(n39433) );
  HS65_LH_BFX2 U23729 ( .A(n39435), .Z(n39434) );
  HS65_LH_BFX2 U23730 ( .A(n39436), .Z(n39435) );
  HS65_LH_BFX2 U23731 ( .A(n39437), .Z(n39436) );
  HS65_LH_BFX2 U23732 ( .A(n39438), .Z(n39437) );
  HS65_LH_BFX2 U23733 ( .A(n39439), .Z(n39438) );
  HS65_LH_BFX2 U23734 ( .A(n39440), .Z(n39439) );
  HS65_LH_BFX2 U23735 ( .A(n39441), .Z(n39440) );
  HS65_LH_BFX2 U23736 ( .A(n39442), .Z(n39441) );
  HS65_LH_BFX2 U23737 ( .A(n39443), .Z(n39442) );
  HS65_LH_BFX2 U23738 ( .A(n17773), .Z(n39443) );
  HS65_LH_BFX2 U23739 ( .A(n39447), .Z(n39444) );
  HS65_LH_BFX2 U23740 ( .A(n39459), .Z(n39445) );
  HS65_LH_BFX2 U23741 ( .A(n39463), .Z(n39446) );
  HS65_LH_BFX2 U23742 ( .A(n39450), .Z(n39447) );
  HS65_LH_BFX2 U23743 ( .A(n17741), .Z(n39448) );
  HS65_LH_IVX2 U23744 ( .A(n39455), .Z(n39449) );
  HS65_LH_IVX2 U23745 ( .A(n39449), .Z(n39450) );
  HS65_LH_BFX2 U23746 ( .A(n137), .Z(n39451) );
  HS65_LH_BFX2 U23747 ( .A(n39448), .Z(n39452) );
  HS65_LH_BFX2 U23748 ( .A(n39451), .Z(n39453) );
  HS65_LH_IVX2 U23749 ( .A(n39461), .Z(n39454) );
  HS65_LH_IVX2 U23750 ( .A(n39454), .Z(n39455) );
  HS65_LH_BFX2 U23751 ( .A(n39452), .Z(n39456) );
  HS65_LH_BFX2 U23752 ( .A(n39453), .Z(n39457) );
  HS65_LH_IVX2 U23753 ( .A(n39465), .Z(n39458) );
  HS65_LH_IVX2 U23754 ( .A(n39458), .Z(n39459) );
  HS65_LH_IVX2 U23755 ( .A(n39467), .Z(n39460) );
  HS65_LH_IVX2 U23756 ( .A(n39460), .Z(n39461) );
  HS65_LH_IVX2 U23757 ( .A(n39469), .Z(n39462) );
  HS65_LH_IVX2 U23758 ( .A(n39462), .Z(n39463) );
  HS65_LH_IVX2 U23759 ( .A(n39471), .Z(n39464) );
  HS65_LH_IVX2 U23760 ( .A(n39464), .Z(n39465) );
  HS65_LH_IVX2 U23761 ( .A(n39475), .Z(n39466) );
  HS65_LH_IVX2 U23762 ( .A(n39466), .Z(n39467) );
  HS65_LH_IVX2 U23763 ( .A(n39473), .Z(n39468) );
  HS65_LH_IVX2 U23764 ( .A(n39468), .Z(n39469) );
  HS65_LH_IVX2 U23765 ( .A(n39483), .Z(n39470) );
  HS65_LH_IVX2 U23766 ( .A(n39470), .Z(n39471) );
  HS65_LH_IVX2 U23767 ( .A(n39457), .Z(n39472) );
  HS65_LH_IVX2 U23768 ( .A(n39472), .Z(n39473) );
  HS65_LH_IVX2 U23769 ( .A(n39485), .Z(n39474) );
  HS65_LH_IVX2 U23770 ( .A(n39474), .Z(n39475) );
  HS65_LH_BFX2 U23771 ( .A(n15490), .Z(n39476) );
  HS65_LH_BFX2 U23772 ( .A(n39481), .Z(n39477) );
  HS65_LH_IVX2 U23773 ( .A(n17742), .Z(n39478) );
  HS65_LH_IVX2 U23774 ( .A(n39478), .Z(n39479) );
  HS65_LH_IVX2 U23775 ( .A(n17636), .Z(n39480) );
  HS65_LH_IVX2 U23776 ( .A(n39480), .Z(n39481) );
  HS65_LH_IVX2 U23777 ( .A(n39487), .Z(n39482) );
  HS65_LH_IVX2 U23778 ( .A(n39482), .Z(n39483) );
  HS65_LH_IVX2 U23779 ( .A(n39490), .Z(n39484) );
  HS65_LH_IVX2 U23780 ( .A(n39484), .Z(n39485) );
  HS65_LH_IVX2 U23781 ( .A(n39492), .Z(n39486) );
  HS65_LH_IVX2 U23782 ( .A(n39486), .Z(n39487) );
  HS65_LH_BFX2 U23783 ( .A(n17646), .Z(n39488) );
  HS65_LH_IVX2 U23784 ( .A(n39493), .Z(n39489) );
  HS65_LH_IVX2 U23785 ( .A(n39489), .Z(n39490) );
  HS65_LH_IVX2 U23786 ( .A(n39456), .Z(n39491) );
  HS65_LH_IVX2 U23787 ( .A(n39491), .Z(n39492) );
  HS65_LH_BFX2 U23788 ( .A(n39494), .Z(n39493) );
  HS65_LH_BFX2 U23789 ( .A(n39495), .Z(n39494) );
  HS65_LH_BFX2 U23790 ( .A(n27787), .Z(n39495) );
  HS65_LH_BFX2 U23791 ( .A(n15476), .Z(n39496) );
  HS65_LH_BFX2 U23792 ( .A(n18037), .Z(n39497) );
  HS65_LH_BFX2 U23793 ( .A(n39501), .Z(n39498) );
  HS65_LH_BFX2 U23794 ( .A(n39503), .Z(n39499) );
  HS65_LH_IVX2 U23795 ( .A(n39513), .Z(n39500) );
  HS65_LH_IVX2 U23796 ( .A(n39500), .Z(n39501) );
  HS65_LH_IVX2 U23797 ( .A(n39509), .Z(n39502) );
  HS65_LH_IVX2 U23798 ( .A(n39502), .Z(n39503) );
  HS65_LH_BFX2 U23799 ( .A(n38503), .Z(n39504) );
  HS65_LH_BFX2 U23800 ( .A(n38504), .Z(n39505) );
  HS65_LH_BFX2 U23801 ( .A(n39497), .Z(n39506) );
  HS65_LH_BFX2 U23802 ( .A(n39504), .Z(n39507) );
  HS65_LH_IVX2 U23803 ( .A(n39516), .Z(n39508) );
  HS65_LH_IVX2 U23804 ( .A(n39508), .Z(n39509) );
  HS65_LH_BFX2 U23805 ( .A(n39505), .Z(n39510) );
  HS65_LH_BFX2 U23806 ( .A(n39518), .Z(n39511) );
  HS65_LH_BFX2 U23807 ( .A(n39506), .Z(n39512) );
  HS65_LH_BFX2 U23808 ( .A(n39520), .Z(n39513) );
  HS65_LH_BFX2 U23809 ( .A(n39507), .Z(n39514) );
  HS65_LH_IVX2 U23810 ( .A(n39524), .Z(n39515) );
  HS65_LH_IVX2 U23811 ( .A(n39515), .Z(n39516) );
  HS65_LH_BFX2 U23812 ( .A(n39510), .Z(n39517) );
  HS65_LH_BFX2 U23813 ( .A(n39527), .Z(n39518) );
  HS65_LH_BFX2 U23814 ( .A(n39512), .Z(n39519) );
  HS65_LH_BFX2 U23815 ( .A(n39529), .Z(n39520) );
  HS65_LH_BFX2 U23816 ( .A(n39514), .Z(n39521) );
  HS65_LH_BFX2 U23817 ( .A(n39517), .Z(n39522) );
  HS65_LH_IVX2 U23818 ( .A(n39532), .Z(n39523) );
  HS65_LH_IVX2 U23819 ( .A(n39523), .Z(n39524) );
  HS65_LH_IVX2 U23820 ( .A(n39534), .Z(n39525) );
  HS65_LH_IVX2 U23821 ( .A(n39525), .Z(n39526) );
  HS65_LH_BFX2 U23822 ( .A(n39535), .Z(n39527) );
  HS65_LH_BFX2 U23823 ( .A(n39519), .Z(n39528) );
  HS65_LH_BFX2 U23824 ( .A(n39537), .Z(n39529) );
  HS65_LH_BFX2 U23825 ( .A(n39521), .Z(n39530) );
  HS65_LH_IVX2 U23826 ( .A(n39542), .Z(n39531) );
  HS65_LH_IVX2 U23827 ( .A(n39531), .Z(n39532) );
  HS65_LH_IVX2 U23828 ( .A(n39544), .Z(n39533) );
  HS65_LH_IVX2 U23829 ( .A(n39533), .Z(n39534) );
  HS65_LH_BFX2 U23830 ( .A(n39545), .Z(n39535) );
  HS65_LH_BFX2 U23831 ( .A(n39528), .Z(n39536) );
  HS65_LH_BFX2 U23832 ( .A(n39540), .Z(n39537) );
  HS65_LH_BFX2 U23833 ( .A(n39530), .Z(n39538) );
  HS65_LH_IVX2 U23834 ( .A(n39549), .Z(n39539) );
  HS65_LH_IVX2 U23835 ( .A(n39539), .Z(n39540) );
  HS65_LH_IVX2 U23836 ( .A(n39551), .Z(n39541) );
  HS65_LH_IVX2 U23837 ( .A(n39541), .Z(n39542) );
  HS65_LH_IVX2 U23838 ( .A(n39553), .Z(n39543) );
  HS65_LH_IVX2 U23839 ( .A(n39543), .Z(n39544) );
  HS65_LH_BFX2 U23840 ( .A(n39554), .Z(n39545) );
  HS65_LH_BFX2 U23841 ( .A(n39536), .Z(n39546) );
  HS65_LH_BFX2 U23842 ( .A(n39538), .Z(n39547) );
  HS65_LH_IVX2 U23843 ( .A(n39560), .Z(n39548) );
  HS65_LH_IVX2 U23844 ( .A(n39548), .Z(n39549) );
  HS65_LH_IVX2 U23845 ( .A(n39562), .Z(n39550) );
  HS65_LH_IVX2 U23846 ( .A(n39550), .Z(n39551) );
  HS65_LH_IVX2 U23847 ( .A(n39564), .Z(n39552) );
  HS65_LH_IVX2 U23848 ( .A(n39552), .Z(n39553) );
  HS65_LH_BFX2 U23849 ( .A(n25851), .Z(n39554) );
  HS65_LH_BFX2 U23850 ( .A(n39546), .Z(n39555) );
  HS65_LH_BFX2 U23851 ( .A(n39547), .Z(n39556) );
  HS65_LH_IVX2 U23852 ( .A(n39567), .Z(n39557) );
  HS65_LH_IVX2 U23853 ( .A(n39557), .Z(n39558) );
  HS65_LH_IVX2 U23854 ( .A(n39569), .Z(n39559) );
  HS65_LH_IVX2 U23855 ( .A(n39559), .Z(n39560) );
  HS65_LH_IVX2 U23856 ( .A(n39571), .Z(n39561) );
  HS65_LH_IVX2 U23857 ( .A(n39561), .Z(n39562) );
  HS65_LH_IVX2 U23858 ( .A(n39573), .Z(n39563) );
  HS65_LH_IVX2 U23859 ( .A(n39563), .Z(n39564) );
  HS65_LH_BFX2 U23860 ( .A(n39555), .Z(n39565) );
  HS65_LH_IVX2 U23861 ( .A(n39576), .Z(n39566) );
  HS65_LH_IVX2 U23862 ( .A(n39566), .Z(n39567) );
  HS65_LH_IVX2 U23863 ( .A(n39578), .Z(n39568) );
  HS65_LH_IVX2 U23864 ( .A(n39568), .Z(n39569) );
  HS65_LH_IVX2 U23865 ( .A(n39581), .Z(n39570) );
  HS65_LH_IVX2 U23866 ( .A(n39570), .Z(n39571) );
  HS65_LH_IVX2 U23867 ( .A(n39583), .Z(n39572) );
  HS65_LH_IVX2 U23868 ( .A(n39572), .Z(n39573) );
  HS65_LH_BFX2 U23869 ( .A(n39565), .Z(n39574) );
  HS65_LH_IVX2 U23870 ( .A(n39585), .Z(n39575) );
  HS65_LH_IVX2 U23871 ( .A(n39575), .Z(n39576) );
  HS65_LH_IVX2 U23872 ( .A(n39587), .Z(n39577) );
  HS65_LH_IVX2 U23873 ( .A(n39577), .Z(n39578) );
  HS65_LH_BFX2 U23874 ( .A(n39574), .Z(n39579) );
  HS65_LH_IVX2 U23875 ( .A(n39590), .Z(n39580) );
  HS65_LH_IVX2 U23876 ( .A(n39580), .Z(n39581) );
  HS65_LH_IVX2 U23877 ( .A(n39592), .Z(n39582) );
  HS65_LH_IVX2 U23878 ( .A(n39582), .Z(n39583) );
  HS65_LH_IVX2 U23879 ( .A(n39594), .Z(n39584) );
  HS65_LH_IVX2 U23880 ( .A(n39584), .Z(n39585) );
  HS65_LH_IVX2 U23881 ( .A(n39596), .Z(n39586) );
  HS65_LH_IVX2 U23882 ( .A(n39586), .Z(n39587) );
  HS65_LH_BFX2 U23883 ( .A(n39579), .Z(n39588) );
  HS65_LH_IVX2 U23884 ( .A(n39599), .Z(n39589) );
  HS65_LH_IVX2 U23885 ( .A(n39589), .Z(n39590) );
  HS65_LH_IVX2 U23886 ( .A(n39601), .Z(n39591) );
  HS65_LH_IVX2 U23887 ( .A(n39591), .Z(n39592) );
  HS65_LH_IVX2 U23888 ( .A(n39603), .Z(n39593) );
  HS65_LH_IVX2 U23889 ( .A(n39593), .Z(n39594) );
  HS65_LH_IVX2 U23890 ( .A(n39605), .Z(n39595) );
  HS65_LH_IVX2 U23891 ( .A(n39595), .Z(n39596) );
  HS65_LH_BFX2 U23892 ( .A(n39588), .Z(n39597) );
  HS65_LH_IVX2 U23893 ( .A(n39608), .Z(n39598) );
  HS65_LH_IVX2 U23894 ( .A(n39598), .Z(n39599) );
  HS65_LH_IVX2 U23895 ( .A(n39610), .Z(n39600) );
  HS65_LH_IVX2 U23896 ( .A(n39600), .Z(n39601) );
  HS65_LH_IVX2 U23897 ( .A(n39556), .Z(n39602) );
  HS65_LH_IVX2 U23898 ( .A(n39602), .Z(n39603) );
  HS65_LH_IVX2 U23899 ( .A(n39612), .Z(n39604) );
  HS65_LH_IVX2 U23900 ( .A(n39604), .Z(n39605) );
  HS65_LH_BFX2 U23901 ( .A(n39597), .Z(n39606) );
  HS65_LH_IVX2 U23902 ( .A(n39614), .Z(n39607) );
  HS65_LH_IVX2 U23903 ( .A(n39607), .Z(n39608) );
  HS65_LH_IVX2 U23904 ( .A(n26241), .Z(n39609) );
  HS65_LH_IVX2 U23905 ( .A(n39609), .Z(n39610) );
  HS65_LH_BFX2 U23906 ( .A(n39606), .Z(n39611) );
  HS65_LH_BFX2 U23907 ( .A(n39615), .Z(n39612) );
  HS65_LH_BFX2 U23908 ( .A(n39611), .Z(n39613) );
  HS65_LH_BFX2 U23909 ( .A(n39617), .Z(n39614) );
  HS65_LH_BFX2 U23910 ( .A(n39618), .Z(n39615) );
  HS65_LH_BFX2 U23911 ( .A(n39613), .Z(n39616) );
  HS65_LH_BFX2 U23912 ( .A(n39620), .Z(n39617) );
  HS65_LH_BFX2 U23913 ( .A(n39621), .Z(n39618) );
  HS65_LH_BFX2 U23914 ( .A(n39616), .Z(n39619) );
  HS65_LH_BFX2 U23915 ( .A(n39627), .Z(n39620) );
  HS65_LH_BFX2 U23916 ( .A(n39624), .Z(n39621) );
  HS65_LH_BFX2 U23917 ( .A(n39619), .Z(n39622) );
  HS65_LH_IVX2 U23918 ( .A(n18038), .Z(n39623) );
  HS65_LH_IVX2 U23919 ( .A(n39623), .Z(n39624) );
  HS65_LH_IVX2 U23920 ( .A(n39622), .Z(n39625) );
  HS65_LH_IVX2 U23921 ( .A(n39625), .Z(n39626) );
  HS65_LH_BFX2 U23922 ( .A(n15463), .Z(n39627) );
  HS65_LH_BFX2 U23923 ( .A(n40191), .Z(n39628) );
  HS65_LH_BFX2 U23924 ( .A(n40255), .Z(n39629) );
  HS65_LH_BFX2 U23925 ( .A(n39631), .Z(n39630) );
  HS65_LH_BFX2 U23926 ( .A(n39632), .Z(n39631) );
  HS65_LH_BFX2 U23927 ( .A(n39633), .Z(n39632) );
  HS65_LH_BFX2 U23928 ( .A(n39634), .Z(n39633) );
  HS65_LH_BFX2 U23929 ( .A(n39635), .Z(n39634) );
  HS65_LH_BFX2 U23930 ( .A(n39636), .Z(n39635) );
  HS65_LH_BFX2 U23931 ( .A(n39637), .Z(n39636) );
  HS65_LH_BFX2 U23932 ( .A(n39638), .Z(n39637) );
  HS65_LH_BFX2 U23933 ( .A(n39639), .Z(n39638) );
  HS65_LH_BFX2 U23934 ( .A(n39640), .Z(n39639) );
  HS65_LH_BFX2 U23935 ( .A(n39641), .Z(n39640) );
  HS65_LH_BFX2 U23936 ( .A(n39642), .Z(n39641) );
  HS65_LH_BFX2 U23937 ( .A(n39643), .Z(n39642) );
  HS65_LH_BFX2 U23938 ( .A(n39644), .Z(n39643) );
  HS65_LH_BFX2 U23939 ( .A(n39645), .Z(n39644) );
  HS65_LH_BFX2 U23940 ( .A(n39646), .Z(n39645) );
  HS65_LH_BFX2 U23941 ( .A(n39647), .Z(n39646) );
  HS65_LH_BFX2 U23942 ( .A(n39648), .Z(n39647) );
  HS65_LH_BFX2 U23943 ( .A(n39649), .Z(n39648) );
  HS65_LH_BFX2 U23944 ( .A(n39650), .Z(n39649) );
  HS65_LH_BFX2 U23945 ( .A(n17736), .Z(n39650) );
  HS65_LH_BFX2 U23946 ( .A(n39652), .Z(n39651) );
  HS65_LH_BFX2 U23947 ( .A(n39653), .Z(n39652) );
  HS65_LH_BFX2 U23948 ( .A(n39654), .Z(n39653) );
  HS65_LH_BFX2 U23949 ( .A(n39655), .Z(n39654) );
  HS65_LH_BFX2 U23950 ( .A(n39656), .Z(n39655) );
  HS65_LH_BFX2 U23951 ( .A(n39657), .Z(n39656) );
  HS65_LH_BFX2 U23952 ( .A(n39658), .Z(n39657) );
  HS65_LH_BFX2 U23953 ( .A(n39659), .Z(n39658) );
  HS65_LH_BFX2 U23954 ( .A(n39660), .Z(n39659) );
  HS65_LH_BFX2 U23955 ( .A(n39661), .Z(n39660) );
  HS65_LH_BFX2 U23956 ( .A(n39662), .Z(n39661) );
  HS65_LH_BFX2 U23957 ( .A(n39663), .Z(n39662) );
  HS65_LH_BFX2 U23958 ( .A(n39664), .Z(n39663) );
  HS65_LH_BFX2 U23959 ( .A(n39665), .Z(n39664) );
  HS65_LH_BFX2 U23960 ( .A(n39666), .Z(n39665) );
  HS65_LH_BFX2 U23961 ( .A(n39667), .Z(n39666) );
  HS65_LH_BFX2 U23962 ( .A(n39668), .Z(n39667) );
  HS65_LH_BFX2 U23963 ( .A(n39669), .Z(n39668) );
  HS65_LH_BFX2 U23964 ( .A(n39670), .Z(n39669) );
  HS65_LH_BFX2 U23965 ( .A(n39671), .Z(n39670) );
  HS65_LH_BFX2 U23966 ( .A(n17737), .Z(n39671) );
  HS65_LH_BFX2 U23967 ( .A(n39674), .Z(n39672) );
  HS65_LH_IVX2 U23968 ( .A(n39675), .Z(n39673) );
  HS65_LH_IVX2 U23969 ( .A(n39673), .Z(n39674) );
  HS65_LH_BFX2 U23970 ( .A(n39676), .Z(n39675) );
  HS65_LH_BFX2 U23971 ( .A(n39677), .Z(n39676) );
  HS65_LH_BFX2 U23972 ( .A(n39678), .Z(n39677) );
  HS65_LH_BFX2 U23973 ( .A(n39679), .Z(n39678) );
  HS65_LH_BFX2 U23974 ( .A(n39680), .Z(n39679) );
  HS65_LH_BFX2 U23975 ( .A(n39681), .Z(n39680) );
  HS65_LH_BFX2 U23976 ( .A(n39682), .Z(n39681) );
  HS65_LH_BFX2 U23977 ( .A(n39683), .Z(n39682) );
  HS65_LH_BFX2 U23978 ( .A(n39684), .Z(n39683) );
  HS65_LH_BFX2 U23979 ( .A(n39685), .Z(n39684) );
  HS65_LH_BFX2 U23980 ( .A(n39686), .Z(n39685) );
  HS65_LH_BFX2 U23981 ( .A(n39687), .Z(n39686) );
  HS65_LH_BFX2 U23982 ( .A(n39688), .Z(n39687) );
  HS65_LH_BFX2 U23983 ( .A(n39689), .Z(n39688) );
  HS65_LH_BFX2 U23984 ( .A(n39690), .Z(n39689) );
  HS65_LH_BFX2 U23985 ( .A(n39691), .Z(n39690) );
  HS65_LH_BFX2 U23986 ( .A(n39692), .Z(n39691) );
  HS65_LH_BFX2 U23987 ( .A(n39693), .Z(n39692) );
  HS65_LH_BFX2 U23988 ( .A(n39694), .Z(n39693) );
  HS65_LH_BFX2 U23989 ( .A(n17726), .Z(n39694) );
  HS65_LH_BFX2 U23990 ( .A(n39696), .Z(n39695) );
  HS65_LH_BFX2 U23991 ( .A(n39697), .Z(n39696) );
  HS65_LH_BFX2 U23992 ( .A(n39698), .Z(n39697) );
  HS65_LH_BFX2 U23993 ( .A(n39699), .Z(n39698) );
  HS65_LH_BFX2 U23994 ( .A(n39700), .Z(n39699) );
  HS65_LH_BFX2 U23995 ( .A(n39701), .Z(n39700) );
  HS65_LH_BFX2 U23996 ( .A(n39702), .Z(n39701) );
  HS65_LH_BFX2 U23997 ( .A(n39703), .Z(n39702) );
  HS65_LH_BFX2 U23998 ( .A(n39704), .Z(n39703) );
  HS65_LH_BFX2 U23999 ( .A(n39705), .Z(n39704) );
  HS65_LH_BFX2 U24000 ( .A(n39706), .Z(n39705) );
  HS65_LH_BFX2 U24001 ( .A(n39707), .Z(n39706) );
  HS65_LH_BFX2 U24002 ( .A(n39708), .Z(n39707) );
  HS65_LH_BFX2 U24003 ( .A(n39709), .Z(n39708) );
  HS65_LH_BFX2 U24004 ( .A(n39710), .Z(n39709) );
  HS65_LH_BFX2 U24005 ( .A(n39711), .Z(n39710) );
  HS65_LH_BFX2 U24006 ( .A(n39712), .Z(n39711) );
  HS65_LH_BFX2 U24007 ( .A(n39713), .Z(n39712) );
  HS65_LH_BFX2 U24008 ( .A(n39714), .Z(n39713) );
  HS65_LH_BFX2 U24009 ( .A(n39715), .Z(n39714) );
  HS65_LH_BFX2 U24010 ( .A(n17735), .Z(n39715) );
  HS65_LH_BFX2 U24011 ( .A(n40440), .Z(n39716) );
  HS65_LH_BFX2 U24012 ( .A(n39718), .Z(n39717) );
  HS65_LH_BFX2 U24013 ( .A(n39719), .Z(n39718) );
  HS65_LH_BFX2 U24014 ( .A(n39720), .Z(n39719) );
  HS65_LH_BFX2 U24015 ( .A(n39721), .Z(n39720) );
  HS65_LH_BFX2 U24016 ( .A(n39722), .Z(n39721) );
  HS65_LH_BFX2 U24017 ( .A(n39723), .Z(n39722) );
  HS65_LH_BFX2 U24018 ( .A(n39724), .Z(n39723) );
  HS65_LH_BFX2 U24019 ( .A(n39725), .Z(n39724) );
  HS65_LH_BFX2 U24020 ( .A(n39726), .Z(n39725) );
  HS65_LH_BFX2 U24021 ( .A(n39727), .Z(n39726) );
  HS65_LH_BFX2 U24022 ( .A(n39728), .Z(n39727) );
  HS65_LH_BFX2 U24023 ( .A(n39729), .Z(n39728) );
  HS65_LH_BFX2 U24024 ( .A(n39730), .Z(n39729) );
  HS65_LH_BFX2 U24025 ( .A(n39731), .Z(n39730) );
  HS65_LH_BFX2 U24026 ( .A(n39732), .Z(n39731) );
  HS65_LH_BFX2 U24027 ( .A(n39733), .Z(n39732) );
  HS65_LH_BFX2 U24028 ( .A(n39734), .Z(n39733) );
  HS65_LH_BFX2 U24029 ( .A(n39735), .Z(n39734) );
  HS65_LH_BFX2 U24030 ( .A(n39736), .Z(n39735) );
  HS65_LH_BFX2 U24031 ( .A(n39737), .Z(n39736) );
  HS65_LH_BFX2 U24032 ( .A(n39738), .Z(n39737) );
  HS65_LH_BFX2 U24033 ( .A(n17814), .Z(n39738) );
  HS65_LH_BFX2 U24034 ( .A(n39740), .Z(n39739) );
  HS65_LH_BFX2 U24035 ( .A(n39741), .Z(n39740) );
  HS65_LH_BFX2 U24036 ( .A(n39742), .Z(n39741) );
  HS65_LH_BFX2 U24037 ( .A(n39743), .Z(n39742) );
  HS65_LH_BFX2 U24038 ( .A(n39744), .Z(n39743) );
  HS65_LH_BFX2 U24039 ( .A(n39745), .Z(n39744) );
  HS65_LH_BFX2 U24040 ( .A(n39746), .Z(n39745) );
  HS65_LH_BFX2 U24041 ( .A(n39747), .Z(n39746) );
  HS65_LH_BFX2 U24042 ( .A(n39748), .Z(n39747) );
  HS65_LH_BFX2 U24043 ( .A(n39749), .Z(n39748) );
  HS65_LH_BFX2 U24044 ( .A(n39750), .Z(n39749) );
  HS65_LH_BFX2 U24045 ( .A(n39751), .Z(n39750) );
  HS65_LH_BFX2 U24046 ( .A(n39752), .Z(n39751) );
  HS65_LH_BFX2 U24047 ( .A(n39753), .Z(n39752) );
  HS65_LH_BFX2 U24048 ( .A(n39754), .Z(n39753) );
  HS65_LH_BFX2 U24049 ( .A(n39755), .Z(n39754) );
  HS65_LH_BFX2 U24050 ( .A(n39756), .Z(n39755) );
  HS65_LH_BFX2 U24051 ( .A(n39757), .Z(n39756) );
  HS65_LH_BFX2 U24052 ( .A(n39758), .Z(n39757) );
  HS65_LH_BFX2 U24053 ( .A(n39759), .Z(n39758) );
  HS65_LH_BFX2 U24054 ( .A(n39760), .Z(n39759) );
  HS65_LH_BFX2 U24055 ( .A(n17730), .Z(n39760) );
  HS65_LH_BFX2 U24056 ( .A(n39762), .Z(n39761) );
  HS65_LH_BFX2 U24057 ( .A(n39763), .Z(n39762) );
  HS65_LH_BFX2 U24058 ( .A(n39764), .Z(n39763) );
  HS65_LH_BFX2 U24059 ( .A(n39765), .Z(n39764) );
  HS65_LH_BFX2 U24060 ( .A(n39766), .Z(n39765) );
  HS65_LH_BFX2 U24061 ( .A(n39767), .Z(n39766) );
  HS65_LH_BFX2 U24062 ( .A(n39768), .Z(n39767) );
  HS65_LH_BFX2 U24063 ( .A(n39769), .Z(n39768) );
  HS65_LH_BFX2 U24064 ( .A(n39770), .Z(n39769) );
  HS65_LH_BFX2 U24065 ( .A(n39771), .Z(n39770) );
  HS65_LH_BFX2 U24066 ( .A(n39772), .Z(n39771) );
  HS65_LH_BFX2 U24067 ( .A(n39773), .Z(n39772) );
  HS65_LH_BFX2 U24068 ( .A(n39774), .Z(n39773) );
  HS65_LH_BFX2 U24069 ( .A(n39775), .Z(n39774) );
  HS65_LH_BFX2 U24070 ( .A(n39776), .Z(n39775) );
  HS65_LH_BFX2 U24071 ( .A(n39777), .Z(n39776) );
  HS65_LH_BFX2 U24072 ( .A(n39778), .Z(n39777) );
  HS65_LH_BFX2 U24073 ( .A(n39779), .Z(n39778) );
  HS65_LH_BFX2 U24074 ( .A(n39780), .Z(n39779) );
  HS65_LH_BFX2 U24075 ( .A(n39781), .Z(n39780) );
  HS65_LH_BFX2 U24076 ( .A(n39782), .Z(n39781) );
  HS65_LH_BFX2 U24077 ( .A(n17731), .Z(n39782) );
  HS65_LH_BFX2 U24078 ( .A(n39784), .Z(n39783) );
  HS65_LH_BFX2 U24079 ( .A(n39785), .Z(n39784) );
  HS65_LH_BFX2 U24080 ( .A(n39786), .Z(n39785) );
  HS65_LH_BFX2 U24081 ( .A(n39787), .Z(n39786) );
  HS65_LH_BFX2 U24082 ( .A(n39788), .Z(n39787) );
  HS65_LH_BFX2 U24083 ( .A(n39789), .Z(n39788) );
  HS65_LH_BFX2 U24084 ( .A(n39790), .Z(n39789) );
  HS65_LH_BFX2 U24085 ( .A(n39791), .Z(n39790) );
  HS65_LH_BFX2 U24086 ( .A(n39792), .Z(n39791) );
  HS65_LH_BFX2 U24087 ( .A(n39793), .Z(n39792) );
  HS65_LH_BFX2 U24088 ( .A(n39794), .Z(n39793) );
  HS65_LH_BFX2 U24089 ( .A(n39795), .Z(n39794) );
  HS65_LH_BFX2 U24090 ( .A(n39796), .Z(n39795) );
  HS65_LH_BFX2 U24091 ( .A(n39797), .Z(n39796) );
  HS65_LH_BFX2 U24092 ( .A(n39798), .Z(n39797) );
  HS65_LH_BFX2 U24093 ( .A(n39799), .Z(n39798) );
  HS65_LH_BFX2 U24094 ( .A(n39800), .Z(n39799) );
  HS65_LH_BFX2 U24095 ( .A(n39801), .Z(n39800) );
  HS65_LH_BFX2 U24096 ( .A(n39802), .Z(n39801) );
  HS65_LH_BFX2 U24097 ( .A(n39803), .Z(n39802) );
  HS65_LH_BFX2 U24098 ( .A(n39804), .Z(n39803) );
  HS65_LH_BFX2 U24099 ( .A(n17809), .Z(n39804) );
  HS65_LH_BFX2 U24100 ( .A(n39806), .Z(n39805) );
  HS65_LH_BFX2 U24101 ( .A(n39807), .Z(n39806) );
  HS65_LH_BFX2 U24102 ( .A(n39808), .Z(n39807) );
  HS65_LH_BFX2 U24103 ( .A(n39809), .Z(n39808) );
  HS65_LH_BFX2 U24104 ( .A(n39810), .Z(n39809) );
  HS65_LH_BFX2 U24105 ( .A(n39811), .Z(n39810) );
  HS65_LH_BFX2 U24106 ( .A(n39812), .Z(n39811) );
  HS65_LH_BFX2 U24107 ( .A(n39813), .Z(n39812) );
  HS65_LH_BFX2 U24108 ( .A(n39814), .Z(n39813) );
  HS65_LH_BFX2 U24109 ( .A(n39815), .Z(n39814) );
  HS65_LH_BFX2 U24110 ( .A(n39816), .Z(n39815) );
  HS65_LH_BFX2 U24111 ( .A(n39817), .Z(n39816) );
  HS65_LH_BFX2 U24112 ( .A(n39818), .Z(n39817) );
  HS65_LH_BFX2 U24113 ( .A(n39819), .Z(n39818) );
  HS65_LH_BFX2 U24114 ( .A(n39820), .Z(n39819) );
  HS65_LH_BFX2 U24115 ( .A(n39821), .Z(n39820) );
  HS65_LH_BFX2 U24116 ( .A(n39822), .Z(n39821) );
  HS65_LH_BFX2 U24117 ( .A(n39823), .Z(n39822) );
  HS65_LH_BFX2 U24118 ( .A(n39824), .Z(n39823) );
  HS65_LH_BFX2 U24119 ( .A(n39825), .Z(n39824) );
  HS65_LH_BFX2 U24120 ( .A(n39826), .Z(n39825) );
  HS65_LH_BFX2 U24121 ( .A(n17813), .Z(n39826) );
  HS65_LH_BFX2 U24122 ( .A(n40482), .Z(n39827) );
  HS65_LH_BFX2 U24123 ( .A(n39829), .Z(n39828) );
  HS65_LH_BFX2 U24124 ( .A(n39830), .Z(n39829) );
  HS65_LH_BFX2 U24125 ( .A(n39831), .Z(n39830) );
  HS65_LH_BFX2 U24126 ( .A(n39832), .Z(n39831) );
  HS65_LH_BFX2 U24127 ( .A(n39833), .Z(n39832) );
  HS65_LH_BFX2 U24128 ( .A(n39834), .Z(n39833) );
  HS65_LH_BFX2 U24129 ( .A(n39835), .Z(n39834) );
  HS65_LH_BFX2 U24130 ( .A(n39836), .Z(n39835) );
  HS65_LH_BFX2 U24131 ( .A(n39837), .Z(n39836) );
  HS65_LH_BFX2 U24132 ( .A(n39838), .Z(n39837) );
  HS65_LH_BFX2 U24133 ( .A(n39839), .Z(n39838) );
  HS65_LH_BFX2 U24134 ( .A(n39840), .Z(n39839) );
  HS65_LH_BFX2 U24135 ( .A(n39841), .Z(n39840) );
  HS65_LH_BFX2 U24136 ( .A(n39842), .Z(n39841) );
  HS65_LH_BFX2 U24137 ( .A(n39843), .Z(n39842) );
  HS65_LH_BFX2 U24138 ( .A(n39844), .Z(n39843) );
  HS65_LH_BFX2 U24139 ( .A(n39845), .Z(n39844) );
  HS65_LH_BFX2 U24140 ( .A(n39846), .Z(n39845) );
  HS65_LH_BFX2 U24141 ( .A(n39847), .Z(n39846) );
  HS65_LH_BFX2 U24142 ( .A(n39848), .Z(n39847) );
  HS65_LH_BFX2 U24143 ( .A(n39849), .Z(n39848) );
  HS65_LH_BFX2 U24144 ( .A(n17734), .Z(n39849) );
  HS65_LH_BFX2 U24145 ( .A(n39851), .Z(n39850) );
  HS65_LH_BFX2 U24146 ( .A(n39852), .Z(n39851) );
  HS65_LH_BFX2 U24147 ( .A(n39853), .Z(n39852) );
  HS65_LH_BFX2 U24148 ( .A(n39854), .Z(n39853) );
  HS65_LH_BFX2 U24149 ( .A(n39855), .Z(n39854) );
  HS65_LH_BFX2 U24150 ( .A(n39856), .Z(n39855) );
  HS65_LH_BFX2 U24151 ( .A(n39857), .Z(n39856) );
  HS65_LH_BFX2 U24152 ( .A(n39858), .Z(n39857) );
  HS65_LH_BFX2 U24153 ( .A(n39859), .Z(n39858) );
  HS65_LH_BFX2 U24154 ( .A(n39860), .Z(n39859) );
  HS65_LH_BFX2 U24155 ( .A(n39861), .Z(n39860) );
  HS65_LH_BFX2 U24156 ( .A(n39862), .Z(n39861) );
  HS65_LH_BFX2 U24157 ( .A(n39863), .Z(n39862) );
  HS65_LH_BFX2 U24158 ( .A(n39864), .Z(n39863) );
  HS65_LH_BFX2 U24159 ( .A(n39865), .Z(n39864) );
  HS65_LH_BFX2 U24160 ( .A(n39866), .Z(n39865) );
  HS65_LH_BFX2 U24161 ( .A(n39867), .Z(n39866) );
  HS65_LH_BFX2 U24162 ( .A(n39868), .Z(n39867) );
  HS65_LH_BFX2 U24163 ( .A(n39869), .Z(n39868) );
  HS65_LH_BFX2 U24164 ( .A(n39870), .Z(n39869) );
  HS65_LH_BFX2 U24165 ( .A(n39871), .Z(n39870) );
  HS65_LH_BFX2 U24166 ( .A(n17796), .Z(n39871) );
  HS65_LH_BFX2 U24167 ( .A(n39873), .Z(n39872) );
  HS65_LH_BFX2 U24168 ( .A(n39874), .Z(n39873) );
  HS65_LH_BFX2 U24169 ( .A(n39875), .Z(n39874) );
  HS65_LH_BFX2 U24170 ( .A(n39876), .Z(n39875) );
  HS65_LH_BFX2 U24171 ( .A(n39877), .Z(n39876) );
  HS65_LH_BFX2 U24172 ( .A(n39878), .Z(n39877) );
  HS65_LH_BFX2 U24173 ( .A(n39879), .Z(n39878) );
  HS65_LH_BFX2 U24174 ( .A(n39880), .Z(n39879) );
  HS65_LH_BFX2 U24175 ( .A(n39881), .Z(n39880) );
  HS65_LH_BFX2 U24176 ( .A(n39882), .Z(n39881) );
  HS65_LH_BFX2 U24177 ( .A(n39883), .Z(n39882) );
  HS65_LH_BFX2 U24178 ( .A(n39884), .Z(n39883) );
  HS65_LH_BFX2 U24179 ( .A(n39885), .Z(n39884) );
  HS65_LH_BFX2 U24180 ( .A(n39886), .Z(n39885) );
  HS65_LH_BFX2 U24181 ( .A(n39887), .Z(n39886) );
  HS65_LH_BFX2 U24182 ( .A(n39888), .Z(n39887) );
  HS65_LH_BFX2 U24183 ( .A(n39889), .Z(n39888) );
  HS65_LH_BFX2 U24184 ( .A(n39890), .Z(n39889) );
  HS65_LH_BFX2 U24185 ( .A(n39891), .Z(n39890) );
  HS65_LH_BFX2 U24186 ( .A(n39892), .Z(n39891) );
  HS65_LH_BFX2 U24187 ( .A(n39893), .Z(n39892) );
  HS65_LH_BFX2 U24188 ( .A(n17797), .Z(n39893) );
  HS65_LH_BFX2 U24189 ( .A(n39895), .Z(n39894) );
  HS65_LH_BFX2 U24190 ( .A(n39896), .Z(n39895) );
  HS65_LH_BFX2 U24191 ( .A(n39897), .Z(n39896) );
  HS65_LH_BFX2 U24192 ( .A(n39898), .Z(n39897) );
  HS65_LH_BFX2 U24193 ( .A(n39899), .Z(n39898) );
  HS65_LH_BFX2 U24194 ( .A(n39900), .Z(n39899) );
  HS65_LH_BFX2 U24195 ( .A(n39901), .Z(n39900) );
  HS65_LH_BFX2 U24196 ( .A(n39902), .Z(n39901) );
  HS65_LH_BFX2 U24197 ( .A(n39903), .Z(n39902) );
  HS65_LH_BFX2 U24198 ( .A(n39904), .Z(n39903) );
  HS65_LH_BFX2 U24199 ( .A(n39905), .Z(n39904) );
  HS65_LH_BFX2 U24200 ( .A(n39906), .Z(n39905) );
  HS65_LH_BFX2 U24201 ( .A(n39907), .Z(n39906) );
  HS65_LH_BFX2 U24202 ( .A(n39908), .Z(n39907) );
  HS65_LH_BFX2 U24203 ( .A(n39909), .Z(n39908) );
  HS65_LH_BFX2 U24204 ( .A(n39910), .Z(n39909) );
  HS65_LH_BFX2 U24205 ( .A(n39911), .Z(n39910) );
  HS65_LH_BFX2 U24206 ( .A(n39912), .Z(n39911) );
  HS65_LH_BFX2 U24207 ( .A(n39913), .Z(n39912) );
  HS65_LH_BFX2 U24208 ( .A(n39914), .Z(n39913) );
  HS65_LH_BFX2 U24209 ( .A(n39915), .Z(n39914) );
  HS65_LH_BFX2 U24210 ( .A(n17798), .Z(n39915) );
  HS65_LH_BFX2 U24211 ( .A(n39917), .Z(n39916) );
  HS65_LH_BFX2 U24212 ( .A(n39918), .Z(n39917) );
  HS65_LH_BFX2 U24213 ( .A(n39919), .Z(n39918) );
  HS65_LH_BFX2 U24214 ( .A(n39920), .Z(n39919) );
  HS65_LH_BFX2 U24215 ( .A(n39921), .Z(n39920) );
  HS65_LH_BFX2 U24216 ( .A(n39922), .Z(n39921) );
  HS65_LH_BFX2 U24217 ( .A(n39923), .Z(n39922) );
  HS65_LH_BFX2 U24218 ( .A(n39924), .Z(n39923) );
  HS65_LH_BFX2 U24219 ( .A(n39925), .Z(n39924) );
  HS65_LH_BFX2 U24220 ( .A(n39926), .Z(n39925) );
  HS65_LH_BFX2 U24221 ( .A(n39927), .Z(n39926) );
  HS65_LH_BFX2 U24222 ( .A(n39928), .Z(n39927) );
  HS65_LH_BFX2 U24223 ( .A(n39929), .Z(n39928) );
  HS65_LH_BFX2 U24224 ( .A(n39930), .Z(n39929) );
  HS65_LH_BFX2 U24225 ( .A(n39931), .Z(n39930) );
  HS65_LH_BFX2 U24226 ( .A(n39932), .Z(n39931) );
  HS65_LH_BFX2 U24227 ( .A(n39933), .Z(n39932) );
  HS65_LH_BFX2 U24228 ( .A(n39934), .Z(n39933) );
  HS65_LH_BFX2 U24229 ( .A(n39935), .Z(n39934) );
  HS65_LH_BFX2 U24230 ( .A(n39936), .Z(n39935) );
  HS65_LH_BFX2 U24231 ( .A(n39937), .Z(n39936) );
  HS65_LH_BFX2 U24232 ( .A(n17799), .Z(n39937) );
  HS65_LH_BFX2 U24233 ( .A(n39939), .Z(n39938) );
  HS65_LH_BFX2 U24234 ( .A(n39940), .Z(n39939) );
  HS65_LH_BFX2 U24235 ( .A(n39941), .Z(n39940) );
  HS65_LH_BFX2 U24236 ( .A(n39942), .Z(n39941) );
  HS65_LH_BFX2 U24237 ( .A(n39943), .Z(n39942) );
  HS65_LH_BFX2 U24238 ( .A(n39944), .Z(n39943) );
  HS65_LH_BFX2 U24239 ( .A(n39945), .Z(n39944) );
  HS65_LH_BFX2 U24240 ( .A(n39946), .Z(n39945) );
  HS65_LH_BFX2 U24241 ( .A(n39947), .Z(n39946) );
  HS65_LH_BFX2 U24242 ( .A(n39948), .Z(n39947) );
  HS65_LH_BFX2 U24243 ( .A(n39949), .Z(n39948) );
  HS65_LH_BFX2 U24244 ( .A(n39950), .Z(n39949) );
  HS65_LH_BFX2 U24245 ( .A(n39951), .Z(n39950) );
  HS65_LH_BFX2 U24246 ( .A(n39952), .Z(n39951) );
  HS65_LH_BFX2 U24247 ( .A(n39953), .Z(n39952) );
  HS65_LH_BFX2 U24248 ( .A(n39954), .Z(n39953) );
  HS65_LH_BFX2 U24249 ( .A(n39955), .Z(n39954) );
  HS65_LH_BFX2 U24250 ( .A(n39956), .Z(n39955) );
  HS65_LH_BFX2 U24251 ( .A(n39957), .Z(n39956) );
  HS65_LH_BFX2 U24252 ( .A(n39958), .Z(n39957) );
  HS65_LH_BFX2 U24253 ( .A(n39959), .Z(n39958) );
  HS65_LH_BFX2 U24254 ( .A(n17800), .Z(n39959) );
  HS65_LH_BFX2 U24255 ( .A(n39961), .Z(n39960) );
  HS65_LH_BFX2 U24256 ( .A(n39962), .Z(n39961) );
  HS65_LH_BFX2 U24257 ( .A(n39963), .Z(n39962) );
  HS65_LH_BFX2 U24258 ( .A(n39964), .Z(n39963) );
  HS65_LH_BFX2 U24259 ( .A(n39965), .Z(n39964) );
  HS65_LH_BFX2 U24260 ( .A(n39966), .Z(n39965) );
  HS65_LH_BFX2 U24261 ( .A(n39967), .Z(n39966) );
  HS65_LH_BFX2 U24262 ( .A(n39968), .Z(n39967) );
  HS65_LH_BFX2 U24263 ( .A(n39969), .Z(n39968) );
  HS65_LH_BFX2 U24264 ( .A(n39970), .Z(n39969) );
  HS65_LH_BFX2 U24265 ( .A(n39971), .Z(n39970) );
  HS65_LH_BFX2 U24266 ( .A(n39972), .Z(n39971) );
  HS65_LH_BFX2 U24267 ( .A(n39973), .Z(n39972) );
  HS65_LH_BFX2 U24268 ( .A(n39974), .Z(n39973) );
  HS65_LH_BFX2 U24269 ( .A(n39975), .Z(n39974) );
  HS65_LH_BFX2 U24270 ( .A(n39976), .Z(n39975) );
  HS65_LH_BFX2 U24271 ( .A(n39977), .Z(n39976) );
  HS65_LH_BFX2 U24272 ( .A(n39978), .Z(n39977) );
  HS65_LH_BFX2 U24273 ( .A(n39979), .Z(n39978) );
  HS65_LH_BFX2 U24274 ( .A(n39980), .Z(n39979) );
  HS65_LH_BFX2 U24275 ( .A(n39981), .Z(n39980) );
  HS65_LH_BFX2 U24276 ( .A(n17802), .Z(n39981) );
  HS65_LH_BFX2 U24277 ( .A(n39983), .Z(n39982) );
  HS65_LH_BFX2 U24278 ( .A(n39984), .Z(n39983) );
  HS65_LH_BFX2 U24279 ( .A(n39985), .Z(n39984) );
  HS65_LH_BFX2 U24280 ( .A(n39986), .Z(n39985) );
  HS65_LH_BFX2 U24281 ( .A(n39987), .Z(n39986) );
  HS65_LH_BFX2 U24282 ( .A(n39988), .Z(n39987) );
  HS65_LH_BFX2 U24283 ( .A(n39989), .Z(n39988) );
  HS65_LH_BFX2 U24284 ( .A(n39990), .Z(n39989) );
  HS65_LH_BFX2 U24285 ( .A(n39991), .Z(n39990) );
  HS65_LH_BFX2 U24286 ( .A(n39992), .Z(n39991) );
  HS65_LH_BFX2 U24287 ( .A(n39993), .Z(n39992) );
  HS65_LH_BFX2 U24288 ( .A(n39994), .Z(n39993) );
  HS65_LH_BFX2 U24289 ( .A(n39995), .Z(n39994) );
  HS65_LH_BFX2 U24290 ( .A(n39996), .Z(n39995) );
  HS65_LH_BFX2 U24291 ( .A(n39997), .Z(n39996) );
  HS65_LH_BFX2 U24292 ( .A(n39998), .Z(n39997) );
  HS65_LH_BFX2 U24293 ( .A(n39999), .Z(n39998) );
  HS65_LH_BFX2 U24294 ( .A(n40000), .Z(n39999) );
  HS65_LH_BFX2 U24295 ( .A(n40001), .Z(n40000) );
  HS65_LH_BFX2 U24296 ( .A(n40002), .Z(n40001) );
  HS65_LH_BFX2 U24297 ( .A(n40003), .Z(n40002) );
  HS65_LH_BFX2 U24298 ( .A(n17803), .Z(n40003) );
  HS65_LH_BFX2 U24299 ( .A(n40005), .Z(n40004) );
  HS65_LH_BFX2 U24300 ( .A(n40006), .Z(n40005) );
  HS65_LH_BFX2 U24301 ( .A(n40007), .Z(n40006) );
  HS65_LH_BFX2 U24302 ( .A(n40008), .Z(n40007) );
  HS65_LH_BFX2 U24303 ( .A(n40009), .Z(n40008) );
  HS65_LH_BFX2 U24304 ( .A(n40010), .Z(n40009) );
  HS65_LH_BFX2 U24305 ( .A(n40011), .Z(n40010) );
  HS65_LH_BFX2 U24306 ( .A(n40012), .Z(n40011) );
  HS65_LH_BFX2 U24307 ( .A(n40013), .Z(n40012) );
  HS65_LH_BFX2 U24308 ( .A(n40014), .Z(n40013) );
  HS65_LH_BFX2 U24309 ( .A(n40015), .Z(n40014) );
  HS65_LH_BFX2 U24310 ( .A(n40016), .Z(n40015) );
  HS65_LH_BFX2 U24311 ( .A(n40017), .Z(n40016) );
  HS65_LH_BFX2 U24312 ( .A(n40018), .Z(n40017) );
  HS65_LH_BFX2 U24313 ( .A(n40019), .Z(n40018) );
  HS65_LH_BFX2 U24314 ( .A(n40020), .Z(n40019) );
  HS65_LH_BFX2 U24315 ( .A(n40021), .Z(n40020) );
  HS65_LH_BFX2 U24316 ( .A(n40022), .Z(n40021) );
  HS65_LH_BFX2 U24317 ( .A(n40023), .Z(n40022) );
  HS65_LH_BFX2 U24318 ( .A(n40024), .Z(n40023) );
  HS65_LH_BFX2 U24319 ( .A(n40025), .Z(n40024) );
  HS65_LH_BFX2 U24320 ( .A(n17804), .Z(n40025) );
  HS65_LH_BFX2 U24321 ( .A(n40027), .Z(n40026) );
  HS65_LH_BFX2 U24322 ( .A(n40028), .Z(n40027) );
  HS65_LH_BFX2 U24323 ( .A(n40029), .Z(n40028) );
  HS65_LH_BFX2 U24324 ( .A(n40030), .Z(n40029) );
  HS65_LH_BFX2 U24325 ( .A(n40031), .Z(n40030) );
  HS65_LH_BFX2 U24326 ( .A(n40032), .Z(n40031) );
  HS65_LH_BFX2 U24327 ( .A(n40033), .Z(n40032) );
  HS65_LH_BFX2 U24328 ( .A(n40034), .Z(n40033) );
  HS65_LH_BFX2 U24329 ( .A(n40035), .Z(n40034) );
  HS65_LH_BFX2 U24330 ( .A(n40036), .Z(n40035) );
  HS65_LH_BFX2 U24331 ( .A(n40037), .Z(n40036) );
  HS65_LH_BFX2 U24332 ( .A(n40038), .Z(n40037) );
  HS65_LH_BFX2 U24333 ( .A(n40039), .Z(n40038) );
  HS65_LH_BFX2 U24334 ( .A(n40040), .Z(n40039) );
  HS65_LH_BFX2 U24335 ( .A(n40041), .Z(n40040) );
  HS65_LH_BFX2 U24336 ( .A(n40042), .Z(n40041) );
  HS65_LH_BFX2 U24337 ( .A(n40043), .Z(n40042) );
  HS65_LH_BFX2 U24338 ( .A(n40044), .Z(n40043) );
  HS65_LH_BFX2 U24339 ( .A(n40045), .Z(n40044) );
  HS65_LH_BFX2 U24340 ( .A(n40046), .Z(n40045) );
  HS65_LH_BFX2 U24341 ( .A(n40047), .Z(n40046) );
  HS65_LH_BFX2 U24342 ( .A(n17805), .Z(n40047) );
  HS65_LH_BFX2 U24343 ( .A(n40049), .Z(n40048) );
  HS65_LH_BFX2 U24344 ( .A(n40050), .Z(n40049) );
  HS65_LH_BFX2 U24345 ( .A(n40051), .Z(n40050) );
  HS65_LH_BFX2 U24346 ( .A(n40052), .Z(n40051) );
  HS65_LH_BFX2 U24347 ( .A(n40053), .Z(n40052) );
  HS65_LH_BFX2 U24348 ( .A(n40054), .Z(n40053) );
  HS65_LH_BFX2 U24349 ( .A(n40055), .Z(n40054) );
  HS65_LH_BFX2 U24350 ( .A(n40056), .Z(n40055) );
  HS65_LH_BFX2 U24351 ( .A(n40057), .Z(n40056) );
  HS65_LH_BFX2 U24352 ( .A(n40058), .Z(n40057) );
  HS65_LH_BFX2 U24353 ( .A(n40059), .Z(n40058) );
  HS65_LH_BFX2 U24354 ( .A(n40060), .Z(n40059) );
  HS65_LH_BFX2 U24355 ( .A(n40061), .Z(n40060) );
  HS65_LH_BFX2 U24356 ( .A(n40062), .Z(n40061) );
  HS65_LH_BFX2 U24357 ( .A(n40063), .Z(n40062) );
  HS65_LH_BFX2 U24358 ( .A(n40064), .Z(n40063) );
  HS65_LH_BFX2 U24359 ( .A(n40065), .Z(n40064) );
  HS65_LH_BFX2 U24360 ( .A(n40066), .Z(n40065) );
  HS65_LH_BFX2 U24361 ( .A(n40067), .Z(n40066) );
  HS65_LH_BFX2 U24362 ( .A(n40068), .Z(n40067) );
  HS65_LH_BFX2 U24363 ( .A(n40069), .Z(n40068) );
  HS65_LH_BFX2 U24364 ( .A(n17806), .Z(n40069) );
  HS65_LH_BFX2 U24365 ( .A(n40071), .Z(n40070) );
  HS65_LH_BFX2 U24366 ( .A(n40072), .Z(n40071) );
  HS65_LH_BFX2 U24367 ( .A(n40073), .Z(n40072) );
  HS65_LH_BFX2 U24368 ( .A(n40074), .Z(n40073) );
  HS65_LH_BFX2 U24369 ( .A(n40075), .Z(n40074) );
  HS65_LH_BFX2 U24370 ( .A(n40076), .Z(n40075) );
  HS65_LH_BFX2 U24371 ( .A(n40077), .Z(n40076) );
  HS65_LH_BFX2 U24372 ( .A(n40078), .Z(n40077) );
  HS65_LH_BFX2 U24373 ( .A(n40079), .Z(n40078) );
  HS65_LH_BFX2 U24374 ( .A(n40080), .Z(n40079) );
  HS65_LH_BFX2 U24375 ( .A(n40081), .Z(n40080) );
  HS65_LH_BFX2 U24376 ( .A(n40082), .Z(n40081) );
  HS65_LH_BFX2 U24377 ( .A(n40083), .Z(n40082) );
  HS65_LH_BFX2 U24378 ( .A(n40084), .Z(n40083) );
  HS65_LH_BFX2 U24379 ( .A(n40085), .Z(n40084) );
  HS65_LH_BFX2 U24380 ( .A(n40086), .Z(n40085) );
  HS65_LH_BFX2 U24381 ( .A(n40087), .Z(n40086) );
  HS65_LH_BFX2 U24382 ( .A(n40088), .Z(n40087) );
  HS65_LH_BFX2 U24383 ( .A(n40089), .Z(n40088) );
  HS65_LH_BFX2 U24384 ( .A(n40090), .Z(n40089) );
  HS65_LH_BFX2 U24385 ( .A(n40091), .Z(n40090) );
  HS65_LH_BFX2 U24386 ( .A(n17807), .Z(n40091) );
  HS65_LH_BFX2 U24387 ( .A(n40093), .Z(n40092) );
  HS65_LH_BFX2 U24388 ( .A(n40094), .Z(n40093) );
  HS65_LH_BFX2 U24389 ( .A(n40095), .Z(n40094) );
  HS65_LH_BFX2 U24390 ( .A(n40096), .Z(n40095) );
  HS65_LH_BFX2 U24391 ( .A(n40097), .Z(n40096) );
  HS65_LH_BFX2 U24392 ( .A(n40098), .Z(n40097) );
  HS65_LH_BFX2 U24393 ( .A(n40099), .Z(n40098) );
  HS65_LH_BFX2 U24394 ( .A(n40100), .Z(n40099) );
  HS65_LH_BFX2 U24395 ( .A(n40101), .Z(n40100) );
  HS65_LH_BFX2 U24396 ( .A(n40102), .Z(n40101) );
  HS65_LH_BFX2 U24397 ( .A(n40103), .Z(n40102) );
  HS65_LH_BFX2 U24398 ( .A(n40104), .Z(n40103) );
  HS65_LH_BFX2 U24399 ( .A(n40105), .Z(n40104) );
  HS65_LH_BFX2 U24400 ( .A(n40106), .Z(n40105) );
  HS65_LH_BFX2 U24401 ( .A(n40107), .Z(n40106) );
  HS65_LH_BFX2 U24402 ( .A(n40108), .Z(n40107) );
  HS65_LH_BFX2 U24403 ( .A(n40109), .Z(n40108) );
  HS65_LH_BFX2 U24404 ( .A(n40110), .Z(n40109) );
  HS65_LH_BFX2 U24405 ( .A(n40111), .Z(n40110) );
  HS65_LH_BFX2 U24406 ( .A(n40112), .Z(n40111) );
  HS65_LH_BFX2 U24407 ( .A(n40113), .Z(n40112) );
  HS65_LH_BFX2 U24408 ( .A(n17808), .Z(n40113) );
  HS65_LH_BFX2 U24409 ( .A(n40115), .Z(n40114) );
  HS65_LH_BFX2 U24410 ( .A(n40116), .Z(n40115) );
  HS65_LH_BFX2 U24411 ( .A(n40117), .Z(n40116) );
  HS65_LH_BFX2 U24412 ( .A(n40118), .Z(n40117) );
  HS65_LH_BFX2 U24413 ( .A(n40119), .Z(n40118) );
  HS65_LH_BFX2 U24414 ( .A(n40120), .Z(n40119) );
  HS65_LH_BFX2 U24415 ( .A(n40121), .Z(n40120) );
  HS65_LH_BFX2 U24416 ( .A(n40122), .Z(n40121) );
  HS65_LH_BFX2 U24417 ( .A(n40123), .Z(n40122) );
  HS65_LH_BFX2 U24418 ( .A(n40124), .Z(n40123) );
  HS65_LH_BFX2 U24419 ( .A(n40125), .Z(n40124) );
  HS65_LH_BFX2 U24420 ( .A(n40126), .Z(n40125) );
  HS65_LH_BFX2 U24421 ( .A(n40127), .Z(n40126) );
  HS65_LH_BFX2 U24422 ( .A(n40128), .Z(n40127) );
  HS65_LH_BFX2 U24423 ( .A(n40129), .Z(n40128) );
  HS65_LH_BFX2 U24424 ( .A(n40130), .Z(n40129) );
  HS65_LH_BFX2 U24425 ( .A(n40131), .Z(n40130) );
  HS65_LH_BFX2 U24426 ( .A(n40132), .Z(n40131) );
  HS65_LH_BFX2 U24427 ( .A(n40133), .Z(n40132) );
  HS65_LH_BFX2 U24428 ( .A(n40134), .Z(n40133) );
  HS65_LH_BFX2 U24429 ( .A(n40135), .Z(n40134) );
  HS65_LH_BFX2 U24430 ( .A(n17810), .Z(n40135) );
  HS65_LH_BFX2 U24431 ( .A(n40137), .Z(n40136) );
  HS65_LH_BFX2 U24432 ( .A(n40138), .Z(n40137) );
  HS65_LH_BFX2 U24433 ( .A(n40139), .Z(n40138) );
  HS65_LH_BFX2 U24434 ( .A(n40140), .Z(n40139) );
  HS65_LH_BFX2 U24435 ( .A(n40141), .Z(n40140) );
  HS65_LH_BFX2 U24436 ( .A(n40142), .Z(n40141) );
  HS65_LH_BFX2 U24437 ( .A(n40143), .Z(n40142) );
  HS65_LH_BFX2 U24438 ( .A(n40144), .Z(n40143) );
  HS65_LH_BFX2 U24439 ( .A(n40145), .Z(n40144) );
  HS65_LH_BFX2 U24440 ( .A(n40146), .Z(n40145) );
  HS65_LH_BFX2 U24441 ( .A(n40147), .Z(n40146) );
  HS65_LH_BFX2 U24442 ( .A(n40148), .Z(n40147) );
  HS65_LH_BFX2 U24443 ( .A(n40149), .Z(n40148) );
  HS65_LH_BFX2 U24444 ( .A(n40150), .Z(n40149) );
  HS65_LH_BFX2 U24445 ( .A(n40151), .Z(n40150) );
  HS65_LH_BFX2 U24446 ( .A(n40152), .Z(n40151) );
  HS65_LH_BFX2 U24447 ( .A(n40153), .Z(n40152) );
  HS65_LH_BFX2 U24448 ( .A(n40154), .Z(n40153) );
  HS65_LH_BFX2 U24449 ( .A(n40155), .Z(n40154) );
  HS65_LH_BFX2 U24450 ( .A(n40156), .Z(n40155) );
  HS65_LH_BFX2 U24451 ( .A(n40157), .Z(n40156) );
  HS65_LH_BFX2 U24452 ( .A(n17812), .Z(n40157) );
  HS65_LH_IVX2 U24453 ( .A(n17645), .Z(n40158) );
  HS65_LH_IVX2 U24454 ( .A(n40158), .Z(n40159) );
  HS65_LH_BFX2 U24455 ( .A(n17693), .Z(n40160) );
  HS65_LH_BFX2 U24456 ( .A(n18082), .Z(n40161) );
  HS65_LH_BFX2 U24457 ( .A(n17710), .Z(n40162) );
  HS65_LH_BFX2 U24458 ( .A(n40170), .Z(n40163) );
  HS65_LH_BFX2 U24459 ( .A(n17575), .Z(n40164) );
  HS65_LH_BFX2 U24460 ( .A(n40164), .Z(n40165) );
  HS65_LH_BFX2 U24461 ( .A(n40165), .Z(n40166) );
  HS65_LH_BFX2 U24462 ( .A(n40166), .Z(n40167) );
  HS65_LH_BFX2 U24463 ( .A(n40167), .Z(n40168) );
  HS65_LH_BFX2 U24464 ( .A(n40168), .Z(n40169) );
  HS65_LH_BFX2 U24465 ( .A(n40171), .Z(n40170) );
  HS65_LH_BFX2 U24466 ( .A(n40172), .Z(n40171) );
  HS65_LH_BFX2 U24467 ( .A(n40173), .Z(n40172) );
  HS65_LH_BFX2 U24468 ( .A(n40174), .Z(n40173) );
  HS65_LH_BFX2 U24469 ( .A(n40175), .Z(n40174) );
  HS65_LH_BFX2 U24470 ( .A(n40176), .Z(n40175) );
  HS65_LH_BFX2 U24471 ( .A(n40177), .Z(n40176) );
  HS65_LH_BFX2 U24472 ( .A(n40178), .Z(n40177) );
  HS65_LH_BFX2 U24473 ( .A(n40179), .Z(n40178) );
  HS65_LH_BFX2 U24474 ( .A(n40180), .Z(n40179) );
  HS65_LH_BFX2 U24475 ( .A(n40181), .Z(n40180) );
  HS65_LH_BFX2 U24476 ( .A(n40182), .Z(n40181) );
  HS65_LH_BFX2 U24477 ( .A(n40183), .Z(n40182) );
  HS65_LH_BFX2 U24478 ( .A(n40169), .Z(n40183) );
  HS65_LH_BFX2 U24479 ( .A(n17581), .Z(n40184) );
  HS65_LH_BFX2 U24480 ( .A(n40184), .Z(n40185) );
  HS65_LH_BFX2 U24481 ( .A(n40185), .Z(n40186) );
  HS65_LH_BFX2 U24482 ( .A(n40186), .Z(n40187) );
  HS65_LH_BFX2 U24483 ( .A(n40187), .Z(n40188) );
  HS65_LH_BFX2 U24484 ( .A(n40188), .Z(n40189) );
  HS65_LH_BFX2 U24485 ( .A(n40189), .Z(n40190) );
  HS65_LH_BFX2 U24486 ( .A(n40192), .Z(n40191) );
  HS65_LH_BFX2 U24487 ( .A(n40193), .Z(n40192) );
  HS65_LH_BFX2 U24488 ( .A(n40194), .Z(n40193) );
  HS65_LH_BFX2 U24489 ( .A(n40195), .Z(n40194) );
  HS65_LH_BFX2 U24490 ( .A(n40196), .Z(n40195) );
  HS65_LH_BFX2 U24491 ( .A(n40197), .Z(n40196) );
  HS65_LH_BFX2 U24492 ( .A(n40198), .Z(n40197) );
  HS65_LH_BFX2 U24493 ( .A(n40199), .Z(n40198) );
  HS65_LH_BFX2 U24494 ( .A(n40200), .Z(n40199) );
  HS65_LH_BFX2 U24495 ( .A(n40201), .Z(n40200) );
  HS65_LH_BFX2 U24496 ( .A(n40202), .Z(n40201) );
  HS65_LH_BFX2 U24497 ( .A(n40203), .Z(n40202) );
  HS65_LH_BFX2 U24498 ( .A(n40204), .Z(n40203) );
  HS65_LH_BFX2 U24499 ( .A(n40190), .Z(n40204) );
  HS65_LH_BFX2 U24500 ( .A(n40206), .Z(n40205) );
  HS65_LH_BFX2 U24501 ( .A(n40207), .Z(n40206) );
  HS65_LH_BFX2 U24502 ( .A(n40208), .Z(n40207) );
  HS65_LH_BFX2 U24503 ( .A(n40209), .Z(n40208) );
  HS65_LH_BFX2 U24504 ( .A(n40210), .Z(n40209) );
  HS65_LH_BFX2 U24505 ( .A(n40211), .Z(n40210) );
  HS65_LH_BFX2 U24506 ( .A(n40212), .Z(n40211) );
  HS65_LH_BFX2 U24507 ( .A(n40213), .Z(n40212) );
  HS65_LH_BFX2 U24508 ( .A(n40214), .Z(n40213) );
  HS65_LH_BFX2 U24509 ( .A(n40215), .Z(n40214) );
  HS65_LH_BFX2 U24510 ( .A(n40216), .Z(n40215) );
  HS65_LH_BFX2 U24511 ( .A(n40217), .Z(n40216) );
  HS65_LH_BFX2 U24512 ( .A(n40218), .Z(n40217) );
  HS65_LH_BFX2 U24513 ( .A(n40219), .Z(n40218) );
  HS65_LH_BFX2 U24514 ( .A(n40220), .Z(n40219) );
  HS65_LH_BFX2 U24515 ( .A(n40221), .Z(n40220) );
  HS65_LH_BFX2 U24516 ( .A(n40222), .Z(n40221) );
  HS65_LH_BFX2 U24517 ( .A(n40223), .Z(n40222) );
  HS65_LH_BFX2 U24518 ( .A(n40224), .Z(n40223) );
  HS65_LH_BFX2 U24519 ( .A(n40225), .Z(n40224) );
  HS65_LH_BFX2 U24520 ( .A(n17740), .Z(n40225) );
  HS65_LH_BFX2 U24521 ( .A(n40227), .Z(n40226) );
  HS65_LH_BFX2 U24522 ( .A(n40718), .Z(n40227) );
  HS65_LH_BFX2 U24523 ( .A(n40236), .Z(n40228) );
  HS65_LH_BFX2 U24524 ( .A(n17586), .Z(n40229) );
  HS65_LH_BFX2 U24525 ( .A(n40229), .Z(n40230) );
  HS65_LH_BFX2 U24526 ( .A(n40230), .Z(n40231) );
  HS65_LH_BFX2 U24527 ( .A(n40231), .Z(n40232) );
  HS65_LH_BFX2 U24528 ( .A(n40232), .Z(n40233) );
  HS65_LH_BFX2 U24529 ( .A(n40233), .Z(n40234) );
  HS65_LH_BFX2 U24530 ( .A(n40234), .Z(n40235) );
  HS65_LH_BFX2 U24531 ( .A(n40237), .Z(n40236) );
  HS65_LH_BFX2 U24532 ( .A(n40238), .Z(n40237) );
  HS65_LH_BFX2 U24533 ( .A(n40239), .Z(n40238) );
  HS65_LH_BFX2 U24534 ( .A(n40240), .Z(n40239) );
  HS65_LH_BFX2 U24535 ( .A(n40241), .Z(n40240) );
  HS65_LH_BFX2 U24536 ( .A(n40242), .Z(n40241) );
  HS65_LH_BFX2 U24537 ( .A(n40243), .Z(n40242) );
  HS65_LH_BFX2 U24538 ( .A(n40244), .Z(n40243) );
  HS65_LH_BFX2 U24539 ( .A(n40245), .Z(n40244) );
  HS65_LH_BFX2 U24540 ( .A(n40246), .Z(n40245) );
  HS65_LH_BFX2 U24541 ( .A(n40247), .Z(n40246) );
  HS65_LH_BFX2 U24542 ( .A(n40248), .Z(n40247) );
  HS65_LH_BFX2 U24543 ( .A(n40235), .Z(n40248) );
  HS65_LH_BFX2 U24544 ( .A(n17626), .Z(n40249) );
  HS65_LH_BFX2 U24545 ( .A(n40249), .Z(n40250) );
  HS65_LH_BFX2 U24546 ( .A(n40250), .Z(n40251) );
  HS65_LH_BFX2 U24547 ( .A(n40251), .Z(n40252) );
  HS65_LH_BFX2 U24548 ( .A(n40252), .Z(n40253) );
  HS65_LH_BFX2 U24549 ( .A(n40253), .Z(n40254) );
  HS65_LH_BFX2 U24550 ( .A(n40256), .Z(n40255) );
  HS65_LH_BFX2 U24551 ( .A(n40257), .Z(n40256) );
  HS65_LH_BFX2 U24552 ( .A(n40258), .Z(n40257) );
  HS65_LH_BFX2 U24553 ( .A(n40259), .Z(n40258) );
  HS65_LH_BFX2 U24554 ( .A(n40260), .Z(n40259) );
  HS65_LH_BFX2 U24555 ( .A(n40261), .Z(n40260) );
  HS65_LH_BFX2 U24556 ( .A(n40262), .Z(n40261) );
  HS65_LH_BFX2 U24557 ( .A(n40263), .Z(n40262) );
  HS65_LH_BFX2 U24558 ( .A(n40264), .Z(n40263) );
  HS65_LH_BFX2 U24559 ( .A(n40265), .Z(n40264) );
  HS65_LH_BFX2 U24560 ( .A(n40266), .Z(n40265) );
  HS65_LH_BFX2 U24561 ( .A(n40267), .Z(n40266) );
  HS65_LH_BFX2 U24562 ( .A(n40268), .Z(n40267) );
  HS65_LH_BFX2 U24563 ( .A(n40269), .Z(n40268) );
  HS65_LH_BFX2 U24564 ( .A(n40254), .Z(n40269) );
  HS65_LH_BFX2 U24565 ( .A(n40271), .Z(n40270) );
  HS65_LH_BFX2 U24566 ( .A(n40272), .Z(n40271) );
  HS65_LH_BFX2 U24567 ( .A(n40273), .Z(n40272) );
  HS65_LH_BFX2 U24568 ( .A(n40274), .Z(n40273) );
  HS65_LH_BFX2 U24569 ( .A(n40275), .Z(n40274) );
  HS65_LH_BFX2 U24570 ( .A(n40276), .Z(n40275) );
  HS65_LH_BFX2 U24571 ( .A(n40277), .Z(n40276) );
  HS65_LH_BFX2 U24572 ( .A(n40278), .Z(n40277) );
  HS65_LH_BFX2 U24573 ( .A(n40279), .Z(n40278) );
  HS65_LH_BFX2 U24574 ( .A(n40280), .Z(n40279) );
  HS65_LH_BFX2 U24575 ( .A(n40281), .Z(n40280) );
  HS65_LH_BFX2 U24576 ( .A(n40282), .Z(n40281) );
  HS65_LH_BFX2 U24577 ( .A(n40283), .Z(n40282) );
  HS65_LH_BFX2 U24578 ( .A(n40284), .Z(n40283) );
  HS65_LH_BFX2 U24579 ( .A(n40285), .Z(n40284) );
  HS65_LH_BFX2 U24580 ( .A(n40286), .Z(n40285) );
  HS65_LH_BFX2 U24581 ( .A(n40287), .Z(n40286) );
  HS65_LH_BFX2 U24582 ( .A(n40288), .Z(n40287) );
  HS65_LH_BFX2 U24583 ( .A(n40289), .Z(n40288) );
  HS65_LH_BFX2 U24584 ( .A(n40290), .Z(n40289) );
  HS65_LH_BFX2 U24585 ( .A(n40291), .Z(n40290) );
  HS65_LH_BFX2 U24586 ( .A(n40292), .Z(n40291) );
  HS65_LH_BFX2 U24587 ( .A(n17765), .Z(n40292) );
  HS65_LH_BFX2 U24588 ( .A(n40294), .Z(n40293) );
  HS65_LH_BFX2 U24589 ( .A(n40295), .Z(n40294) );
  HS65_LH_BFX2 U24590 ( .A(n40296), .Z(n40295) );
  HS65_LH_BFX2 U24591 ( .A(n40297), .Z(n40296) );
  HS65_LH_BFX2 U24592 ( .A(n40298), .Z(n40297) );
  HS65_LH_BFX2 U24593 ( .A(n40299), .Z(n40298) );
  HS65_LH_BFX2 U24594 ( .A(n40300), .Z(n40299) );
  HS65_LH_BFX2 U24595 ( .A(n40301), .Z(n40300) );
  HS65_LH_BFX2 U24596 ( .A(n40302), .Z(n40301) );
  HS65_LH_BFX2 U24597 ( .A(n40303), .Z(n40302) );
  HS65_LH_BFX2 U24598 ( .A(n40304), .Z(n40303) );
  HS65_LH_BFX2 U24599 ( .A(n40305), .Z(n40304) );
  HS65_LH_BFX2 U24600 ( .A(n40306), .Z(n40305) );
  HS65_LH_BFX2 U24601 ( .A(n40307), .Z(n40306) );
  HS65_LH_BFX2 U24602 ( .A(n40308), .Z(n40307) );
  HS65_LH_BFX2 U24603 ( .A(n40309), .Z(n40308) );
  HS65_LH_BFX2 U24604 ( .A(n40310), .Z(n40309) );
  HS65_LH_BFX2 U24605 ( .A(n40311), .Z(n40310) );
  HS65_LH_BFX2 U24606 ( .A(n40312), .Z(n40311) );
  HS65_LH_BFX2 U24607 ( .A(n40313), .Z(n40312) );
  HS65_LH_BFX2 U24608 ( .A(n40314), .Z(n40313) );
  HS65_LH_BFX2 U24609 ( .A(n40315), .Z(n40314) );
  HS65_LH_BFX2 U24610 ( .A(n17767), .Z(n40315) );
  HS65_LH_BFX2 U24611 ( .A(n40317), .Z(n40316) );
  HS65_LH_BFX2 U24612 ( .A(n40318), .Z(n40317) );
  HS65_LH_BFX2 U24613 ( .A(n40319), .Z(n40318) );
  HS65_LH_BFX2 U24614 ( .A(n40320), .Z(n40319) );
  HS65_LH_BFX2 U24615 ( .A(n40321), .Z(n40320) );
  HS65_LH_BFX2 U24616 ( .A(n40322), .Z(n40321) );
  HS65_LH_BFX2 U24617 ( .A(n40323), .Z(n40322) );
  HS65_LH_BFX2 U24618 ( .A(n40324), .Z(n40323) );
  HS65_LH_BFX2 U24619 ( .A(n40325), .Z(n40324) );
  HS65_LH_BFX2 U24620 ( .A(n40326), .Z(n40325) );
  HS65_LH_BFX2 U24621 ( .A(n40327), .Z(n40326) );
  HS65_LH_BFX2 U24622 ( .A(n40328), .Z(n40327) );
  HS65_LH_BFX2 U24623 ( .A(n40329), .Z(n40328) );
  HS65_LH_BFX2 U24624 ( .A(n40330), .Z(n40329) );
  HS65_LH_BFX2 U24625 ( .A(n40331), .Z(n40330) );
  HS65_LH_BFX2 U24626 ( .A(n40332), .Z(n40331) );
  HS65_LH_BFX2 U24627 ( .A(n40333), .Z(n40332) );
  HS65_LH_BFX2 U24628 ( .A(n40334), .Z(n40333) );
  HS65_LH_BFX2 U24629 ( .A(n40335), .Z(n40334) );
  HS65_LH_BFX2 U24630 ( .A(n40336), .Z(n40335) );
  HS65_LH_BFX2 U24631 ( .A(n40337), .Z(n40336) );
  HS65_LH_BFX2 U24632 ( .A(n40338), .Z(n40337) );
  HS65_LH_BFX2 U24633 ( .A(n17952), .Z(n40338) );
  HS65_LH_BFX2 U24634 ( .A(n40340), .Z(n40339) );
  HS65_LH_BFX2 U24635 ( .A(n40341), .Z(n40340) );
  HS65_LH_BFX2 U24636 ( .A(n40342), .Z(n40341) );
  HS65_LH_BFX2 U24637 ( .A(n40343), .Z(n40342) );
  HS65_LH_BFX2 U24638 ( .A(n40344), .Z(n40343) );
  HS65_LH_BFX2 U24639 ( .A(n40345), .Z(n40344) );
  HS65_LH_BFX2 U24640 ( .A(n40346), .Z(n40345) );
  HS65_LH_BFX2 U24641 ( .A(n40347), .Z(n40346) );
  HS65_LH_BFX2 U24642 ( .A(n40348), .Z(n40347) );
  HS65_LH_BFX2 U24643 ( .A(n40349), .Z(n40348) );
  HS65_LH_BFX2 U24644 ( .A(n40350), .Z(n40349) );
  HS65_LH_BFX2 U24645 ( .A(n40351), .Z(n40350) );
  HS65_LH_BFX2 U24646 ( .A(n40352), .Z(n40351) );
  HS65_LH_BFX2 U24647 ( .A(n40353), .Z(n40352) );
  HS65_LH_BFX2 U24648 ( .A(n40354), .Z(n40353) );
  HS65_LH_BFX2 U24649 ( .A(n40355), .Z(n40354) );
  HS65_LH_BFX2 U24650 ( .A(n40356), .Z(n40355) );
  HS65_LH_BFX2 U24651 ( .A(n40357), .Z(n40356) );
  HS65_LH_BFX2 U24652 ( .A(n40358), .Z(n40357) );
  HS65_LH_BFX2 U24653 ( .A(n40359), .Z(n40358) );
  HS65_LH_BFX2 U24654 ( .A(n40360), .Z(n40359) );
  HS65_LH_BFX2 U24655 ( .A(n40361), .Z(n40360) );
  HS65_LH_BFX2 U24656 ( .A(n17939), .Z(n40361) );
  HS65_LH_BFX2 U24657 ( .A(n40363), .Z(n40362) );
  HS65_LH_BFX2 U24658 ( .A(n40364), .Z(n40363) );
  HS65_LH_BFX2 U24659 ( .A(n40365), .Z(n40364) );
  HS65_LH_BFX2 U24660 ( .A(n40366), .Z(n40365) );
  HS65_LH_BFX2 U24661 ( .A(n40367), .Z(n40366) );
  HS65_LH_BFX2 U24662 ( .A(n40368), .Z(n40367) );
  HS65_LH_BFX2 U24663 ( .A(n40369), .Z(n40368) );
  HS65_LH_BFX2 U24664 ( .A(n40370), .Z(n40369) );
  HS65_LH_BFX2 U24665 ( .A(n40371), .Z(n40370) );
  HS65_LH_BFX2 U24666 ( .A(n40372), .Z(n40371) );
  HS65_LH_BFX2 U24667 ( .A(n40373), .Z(n40372) );
  HS65_LH_BFX2 U24668 ( .A(n40374), .Z(n40373) );
  HS65_LH_BFX2 U24669 ( .A(n40375), .Z(n40374) );
  HS65_LH_BFX2 U24670 ( .A(n40376), .Z(n40375) );
  HS65_LH_BFX2 U24671 ( .A(n40377), .Z(n40376) );
  HS65_LH_BFX2 U24672 ( .A(n40378), .Z(n40377) );
  HS65_LH_BFX2 U24673 ( .A(n40379), .Z(n40378) );
  HS65_LH_BFX2 U24674 ( .A(n40380), .Z(n40379) );
  HS65_LH_BFX2 U24675 ( .A(n40381), .Z(n40380) );
  HS65_LH_BFX2 U24676 ( .A(n40382), .Z(n40381) );
  HS65_LH_BFX2 U24677 ( .A(n40383), .Z(n40382) );
  HS65_LH_BFX2 U24678 ( .A(n40384), .Z(n40383) );
  HS65_LH_BFX2 U24679 ( .A(n17962), .Z(n40384) );
  HS65_LH_BFX2 U24680 ( .A(n40386), .Z(n40385) );
  HS65_LH_BFX2 U24681 ( .A(n40387), .Z(n40386) );
  HS65_LH_BFX2 U24682 ( .A(n40388), .Z(n40387) );
  HS65_LH_BFX2 U24683 ( .A(n40389), .Z(n40388) );
  HS65_LH_BFX2 U24684 ( .A(n40390), .Z(n40389) );
  HS65_LH_BFX2 U24685 ( .A(n40391), .Z(n40390) );
  HS65_LH_BFX2 U24686 ( .A(n40392), .Z(n40391) );
  HS65_LH_BFX2 U24687 ( .A(n40393), .Z(n40392) );
  HS65_LH_BFX2 U24688 ( .A(n40394), .Z(n40393) );
  HS65_LH_BFX2 U24689 ( .A(n40395), .Z(n40394) );
  HS65_LH_BFX2 U24690 ( .A(n40396), .Z(n40395) );
  HS65_LH_BFX2 U24691 ( .A(n40397), .Z(n40396) );
  HS65_LH_BFX2 U24693 ( .A(n40398), .Z(n40397) );
  HS65_LH_BFX2 U24694 ( .A(n40399), .Z(n40398) );
  HS65_LH_BFX2 U24695 ( .A(n40400), .Z(n40399) );
  HS65_LH_BFX2 U24696 ( .A(n40401), .Z(n40400) );
  HS65_LH_BFX2 U24697 ( .A(n40402), .Z(n40401) );
  HS65_LH_BFX2 U24698 ( .A(n40403), .Z(n40402) );
  HS65_LH_BFX2 U24699 ( .A(n40404), .Z(n40403) );
  HS65_LH_BFX2 U24700 ( .A(n40405), .Z(n40404) );
  HS65_LH_BFX2 U24701 ( .A(n40406), .Z(n40405) );
  HS65_LH_BFX2 U24702 ( .A(n40407), .Z(n40406) );
  HS65_LH_BFX2 U24703 ( .A(n17913), .Z(n40407) );
  HS65_LH_BFX2 U24704 ( .A(n40409), .Z(n40408) );
  HS65_LH_BFX2 U24705 ( .A(n40410), .Z(n40409) );
  HS65_LH_BFX2 U24706 ( .A(n40411), .Z(n40410) );
  HS65_LH_BFX2 U24707 ( .A(n40412), .Z(n40411) );
  HS65_LH_BFX2 U24708 ( .A(n40413), .Z(n40412) );
  HS65_LH_BFX2 U24709 ( .A(n40414), .Z(n40413) );
  HS65_LH_BFX2 U24710 ( .A(n40415), .Z(n40414) );
  HS65_LH_BFX2 U24711 ( .A(n40416), .Z(n40415) );
  HS65_LH_BFX2 U24712 ( .A(n40417), .Z(n40416) );
  HS65_LH_BFX2 U24713 ( .A(n40418), .Z(n40417) );
  HS65_LH_BFX2 U24714 ( .A(n40419), .Z(n40418) );
  HS65_LH_BFX2 U24715 ( .A(n40420), .Z(n40419) );
  HS65_LH_BFX2 U24716 ( .A(n40421), .Z(n40420) );
  HS65_LH_BFX2 U24717 ( .A(n40422), .Z(n40421) );
  HS65_LH_BFX2 U24718 ( .A(n40423), .Z(n40422) );
  HS65_LH_BFX2 U24719 ( .A(n40424), .Z(n40423) );
  HS65_LH_BFX2 U24720 ( .A(n40425), .Z(n40424) );
  HS65_LH_BFX2 U24721 ( .A(n40426), .Z(n40425) );
  HS65_LH_BFX2 U24722 ( .A(n40427), .Z(n40426) );
  HS65_LH_BFX2 U24723 ( .A(n40428), .Z(n40427) );
  HS65_LH_BFX2 U24724 ( .A(n40429), .Z(n40428) );
  HS65_LH_BFX2 U24725 ( .A(n40430), .Z(n40429) );
  HS65_LH_BFX2 U24726 ( .A(n17994), .Z(n40430) );
  HS65_LH_BFX2 U24727 ( .A(n17583), .Z(n40431) );
  HS65_LH_BFX2 U24728 ( .A(n40431), .Z(n40432) );
  HS65_LH_BFX2 U24729 ( .A(n40432), .Z(n40433) );
  HS65_LH_BFX2 U24730 ( .A(n40433), .Z(n40434) );
  HS65_LH_BFX2 U24731 ( .A(n40434), .Z(n40435) );
  HS65_LH_BFX2 U24732 ( .A(n40435), .Z(n40436) );
  HS65_LH_BFX2 U24733 ( .A(n40436), .Z(n40437) );
  HS65_LH_BFX2 U24734 ( .A(n40437), .Z(n40438) );
  HS65_LH_BFX2 U24735 ( .A(n40438), .Z(n40439) );
  HS65_LH_BFX2 U24736 ( .A(n40441), .Z(n40440) );
  HS65_LH_BFX2 U24737 ( .A(n40442), .Z(n40441) );
  HS65_LH_BFX2 U24738 ( .A(n40443), .Z(n40442) );
  HS65_LH_BFX2 U24739 ( .A(n40444), .Z(n40443) );
  HS65_LH_BFX2 U24740 ( .A(n40445), .Z(n40444) );
  HS65_LH_BFX2 U24741 ( .A(n40446), .Z(n40445) );
  HS65_LH_BFX2 U24742 ( .A(n40447), .Z(n40446) );
  HS65_LH_BFX2 U24743 ( .A(n40448), .Z(n40447) );
  HS65_LH_BFX2 U24744 ( .A(n40449), .Z(n40448) );
  HS65_LH_BFX2 U24745 ( .A(n40450), .Z(n40449) );
  HS65_LH_BFX2 U24746 ( .A(n40451), .Z(n40450) );
  HS65_LH_BFX2 U24747 ( .A(n40439), .Z(n40451) );
  HS65_LH_BFX2 U24748 ( .A(n40453), .Z(n40452) );
  HS65_LH_BFX2 U24749 ( .A(n40454), .Z(n40453) );
  HS65_LH_BFX2 U24750 ( .A(n40455), .Z(n40454) );
  HS65_LH_BFX2 U24751 ( .A(n40456), .Z(n40455) );
  HS65_LH_BFX2 U24752 ( .A(n40457), .Z(n40456) );
  HS65_LH_BFX2 U24753 ( .A(n40458), .Z(n40457) );
  HS65_LH_BFX2 U24754 ( .A(n40459), .Z(n40458) );
  HS65_LH_BFX2 U24755 ( .A(n40460), .Z(n40459) );
  HS65_LH_BFX2 U24756 ( .A(n40461), .Z(n40460) );
  HS65_LH_BFX2 U24757 ( .A(n40462), .Z(n40461) );
  HS65_LH_BFX2 U24758 ( .A(n40463), .Z(n40462) );
  HS65_LH_BFX2 U24759 ( .A(n40464), .Z(n40463) );
  HS65_LH_BFX2 U24760 ( .A(n40465), .Z(n40464) );
  HS65_LH_BFX2 U24761 ( .A(n40466), .Z(n40465) );
  HS65_LH_BFX2 U24762 ( .A(n40467), .Z(n40466) );
  HS65_LH_BFX2 U24763 ( .A(n40468), .Z(n40467) );
  HS65_LH_BFX2 U24764 ( .A(n40469), .Z(n40468) );
  HS65_LH_BFX2 U24765 ( .A(n40470), .Z(n40469) );
  HS65_LH_BFX2 U24766 ( .A(n40471), .Z(n40470) );
  HS65_LH_BFX2 U24767 ( .A(n14300), .Z(n40471) );
  HS65_LH_BFX2 U24768 ( .A(n40473), .Z(n40472) );
  HS65_LH_BFX2 U24769 ( .A(n17593), .Z(n40473) );
  HS65_LH_BFX2 U24770 ( .A(n40477), .Z(n40474) );
  HS65_LH_BFX2 U24771 ( .A(n40479), .Z(n40475) );
  HS65_LH_IVX2 U24772 ( .A(n40606), .Z(n40476) );
  HS65_LH_IVX2 U24773 ( .A(n40476), .Z(n40477) );
  HS65_LH_IVX2 U24774 ( .A(n40480), .Z(n40478) );
  HS65_LH_IVX2 U24775 ( .A(n40478), .Z(n40479) );
  HS65_LH_BFX2 U24776 ( .A(n40715), .Z(n40480) );
  HS65_LH_BFX2 U24777 ( .A(n40713), .Z(n40481) );
  HS65_LH_BFX2 U24778 ( .A(n40483), .Z(n40482) );
  HS65_LH_BFX2 U24779 ( .A(n40484), .Z(n40483) );
  HS65_LH_BFX2 U24780 ( .A(n40485), .Z(n40484) );
  HS65_LH_BFX2 U24781 ( .A(n40486), .Z(n40485) );
  HS65_LH_BFX2 U24782 ( .A(n40487), .Z(n40486) );
  HS65_LH_BFX2 U24783 ( .A(n40488), .Z(n40487) );
  HS65_LH_BFX2 U24784 ( .A(n40489), .Z(n40488) );
  HS65_LH_BFX2 U24785 ( .A(n40490), .Z(n40489) );
  HS65_LH_BFX2 U24786 ( .A(n40491), .Z(n40490) );
  HS65_LH_BFX2 U24787 ( .A(n40492), .Z(n40491) );
  HS65_LH_BFX2 U24788 ( .A(n40493), .Z(n40492) );
  HS65_LH_BFX2 U24789 ( .A(n40494), .Z(n40493) );
  HS65_LH_BFX2 U24790 ( .A(n40495), .Z(n40494) );
  HS65_LH_BFX2 U24791 ( .A(n40496), .Z(n40495) );
  HS65_LH_BFX2 U24792 ( .A(n40497), .Z(n40496) );
  HS65_LH_BFX2 U24793 ( .A(n40498), .Z(n40497) );
  HS65_LH_BFX2 U24794 ( .A(n40499), .Z(n40498) );
  HS65_LH_BFX2 U24795 ( .A(n40500), .Z(n40499) );
  HS65_LH_BFX2 U24796 ( .A(n40501), .Z(n40500) );
  HS65_LH_BFX2 U24797 ( .A(n40502), .Z(n40501) );
  HS65_LH_BFX2 U24798 ( .A(n17811), .Z(n40502) );
  HS65_LH_BFX2 U24799 ( .A(n40504), .Z(n40503) );
  HS65_LH_BFX2 U24800 ( .A(n40505), .Z(n40504) );
  HS65_LH_BFX2 U24801 ( .A(n40506), .Z(n40505) );
  HS65_LH_BFX2 U24802 ( .A(n40507), .Z(n40506) );
  HS65_LH_BFX2 U24803 ( .A(n40508), .Z(n40507) );
  HS65_LH_BFX2 U24804 ( .A(n40509), .Z(n40508) );
  HS65_LH_BFX2 U24805 ( .A(n40510), .Z(n40509) );
  HS65_LH_BFX2 U24806 ( .A(n40511), .Z(n40510) );
  HS65_LH_BFX2 U24807 ( .A(n40512), .Z(n40511) );
  HS65_LH_BFX2 U24808 ( .A(n40513), .Z(n40512) );
  HS65_LH_BFX2 U24809 ( .A(n40514), .Z(n40513) );
  HS65_LH_BFX2 U24810 ( .A(n40515), .Z(n40514) );
  HS65_LH_BFX2 U24811 ( .A(n40516), .Z(n40515) );
  HS65_LH_BFX2 U24812 ( .A(n40517), .Z(n40516) );
  HS65_LH_BFX2 U24813 ( .A(n40518), .Z(n40517) );
  HS65_LH_BFX2 U24814 ( .A(n40519), .Z(n40518) );
  HS65_LH_BFX2 U24815 ( .A(n40520), .Z(n40519) );
  HS65_LH_BFX2 U24816 ( .A(n40521), .Z(n40520) );
  HS65_LH_BFX2 U24817 ( .A(n40522), .Z(n40521) );
  HS65_LH_BFX2 U24818 ( .A(n40523), .Z(n40522) );
  HS65_LH_BFX2 U24819 ( .A(n17815), .Z(n40523) );
  HS65_LH_BFX2 U24820 ( .A(n40525), .Z(n40524) );
  HS65_LH_BFX2 U24821 ( .A(n40526), .Z(n40525) );
  HS65_LH_BFX2 U24822 ( .A(n40527), .Z(n40526) );
  HS65_LH_BFX2 U24823 ( .A(n40528), .Z(n40527) );
  HS65_LH_BFX2 U24824 ( .A(n40529), .Z(n40528) );
  HS65_LH_BFX2 U24825 ( .A(n40530), .Z(n40529) );
  HS65_LH_BFX2 U24826 ( .A(n40531), .Z(n40530) );
  HS65_LH_BFX2 U24827 ( .A(n40532), .Z(n40531) );
  HS65_LH_BFX2 U24828 ( .A(n40533), .Z(n40532) );
  HS65_LH_BFX2 U24829 ( .A(n40534), .Z(n40533) );
  HS65_LH_BFX2 U24830 ( .A(n40535), .Z(n40534) );
  HS65_LH_BFX2 U24831 ( .A(n40536), .Z(n40535) );
  HS65_LH_BFX2 U24832 ( .A(n40537), .Z(n40536) );
  HS65_LH_BFX2 U24833 ( .A(n40538), .Z(n40537) );
  HS65_LH_BFX2 U24834 ( .A(n40539), .Z(n40538) );
  HS65_LH_BFX2 U24835 ( .A(n40540), .Z(n40539) );
  HS65_LH_BFX2 U24836 ( .A(n40541), .Z(n40540) );
  HS65_LH_BFX2 U24837 ( .A(n40542), .Z(n40541) );
  HS65_LH_BFX2 U24838 ( .A(n40543), .Z(n40542) );
  HS65_LH_BFX2 U24839 ( .A(n17571), .Z(n40543) );
  HS65_LH_BFX2 U24840 ( .A(n40545), .Z(n40544) );
  HS65_LH_BFX2 U24841 ( .A(n40546), .Z(n40545) );
  HS65_LH_BFX2 U24842 ( .A(n40547), .Z(n40546) );
  HS65_LH_BFX2 U24843 ( .A(n40548), .Z(n40547) );
  HS65_LH_BFX2 U24844 ( .A(n40549), .Z(n40548) );
  HS65_LH_BFX2 U24845 ( .A(n40550), .Z(n40549) );
  HS65_LH_BFX2 U24846 ( .A(n40551), .Z(n40550) );
  HS65_LH_BFX2 U24847 ( .A(n40552), .Z(n40551) );
  HS65_LH_BFX2 U24848 ( .A(n40553), .Z(n40552) );
  HS65_LH_BFX2 U24849 ( .A(n40554), .Z(n40553) );
  HS65_LH_BFX2 U24850 ( .A(n40555), .Z(n40554) );
  HS65_LH_BFX2 U24851 ( .A(n40556), .Z(n40555) );
  HS65_LH_BFX2 U24852 ( .A(n40557), .Z(n40556) );
  HS65_LH_BFX2 U24853 ( .A(n15200), .Z(n40557) );
  HS65_LH_BFX2 U24854 ( .A(n40559), .Z(n40558) );
  HS65_LH_BFX2 U24855 ( .A(n14511), .Z(n40559) );
  HS65_LH_BFX2 U24856 ( .A(n15396), .Z(n40560) );
  HS65_LH_BFX2 U24857 ( .A(n40562), .Z(n40561) );
  HS65_LH_BFX2 U24858 ( .A(n40563), .Z(n40562) );
  HS65_LH_BFX2 U24859 ( .A(n40564), .Z(n40563) );
  HS65_LH_BFX2 U24860 ( .A(n40565), .Z(n40564) );
  HS65_LH_BFX2 U24861 ( .A(n40566), .Z(n40565) );
  HS65_LH_BFX2 U24862 ( .A(n40567), .Z(n40566) );
  HS65_LH_BFX2 U24863 ( .A(n40568), .Z(n40567) );
  HS65_LH_BFX2 U24864 ( .A(n40569), .Z(n40568) );
  HS65_LH_BFX2 U24865 ( .A(n40570), .Z(n40569) );
  HS65_LH_BFX2 U24866 ( .A(n40571), .Z(n40570) );
  HS65_LH_BFX2 U24867 ( .A(n40572), .Z(n40571) );
  HS65_LH_BFX2 U24868 ( .A(n40573), .Z(n40572) );
  HS65_LH_BFX2 U24869 ( .A(n40574), .Z(n40573) );
  HS65_LH_BFX2 U24870 ( .A(n40575), .Z(n40574) );
  HS65_LH_BFX2 U24871 ( .A(n40576), .Z(n40575) );
  HS65_LH_BFX2 U24872 ( .A(n40577), .Z(n40576) );
  HS65_LH_BFX2 U24873 ( .A(n40578), .Z(n40577) );
  HS65_LH_BFX2 U24874 ( .A(n40579), .Z(n40578) );
  HS65_LH_BFX2 U24875 ( .A(n40580), .Z(n40579) );
  HS65_LH_BFX2 U24876 ( .A(n17755), .Z(n40580) );
  HS65_LH_BFX2 U24877 ( .A(n40582), .Z(n40581) );
  HS65_LH_BFX2 U24878 ( .A(n40583), .Z(n40582) );
  HS65_LH_BFX2 U24879 ( .A(n40584), .Z(n40583) );
  HS65_LH_BFX2 U24880 ( .A(n40585), .Z(n40584) );
  HS65_LH_BFX2 U24881 ( .A(n40586), .Z(n40585) );
  HS65_LH_BFX2 U24882 ( .A(n40587), .Z(n40586) );
  HS65_LH_BFX2 U24883 ( .A(n40588), .Z(n40587) );
  HS65_LH_BFX2 U24884 ( .A(n40589), .Z(n40588) );
  HS65_LH_BFX2 U24885 ( .A(n40590), .Z(n40589) );
  HS65_LH_BFX2 U24886 ( .A(n40591), .Z(n40590) );
  HS65_LH_BFX2 U24887 ( .A(n40592), .Z(n40591) );
  HS65_LH_BFX2 U24888 ( .A(n40593), .Z(n40592) );
  HS65_LH_BFX2 U24889 ( .A(n40594), .Z(n40593) );
  HS65_LH_BFX2 U24890 ( .A(n40595), .Z(n40594) );
  HS65_LH_BFX2 U24891 ( .A(n40596), .Z(n40595) );
  HS65_LH_BFX2 U24892 ( .A(n40597), .Z(n40596) );
  HS65_LH_BFX2 U24893 ( .A(n40598), .Z(n40597) );
  HS65_LH_BFX2 U24894 ( .A(n40599), .Z(n40598) );
  HS65_LH_BFX2 U24895 ( .A(n40600), .Z(n40599) );
  HS65_LH_BFX2 U24896 ( .A(n40601), .Z(n40600) );
  HS65_LH_BFX2 U24897 ( .A(n14876), .Z(n40601) );
  HS65_LH_BFX2 U24898 ( .A(n40615), .Z(n40602) );
  HS65_LH_BFX2 U24899 ( .A(n40605), .Z(n40603) );
  HS65_LH_BFX2 U24900 ( .A(n40612), .Z(n40604) );
  HS65_LH_BFX2 U24901 ( .A(n40717), .Z(n40605) );
  HS65_LH_BFX2 U24902 ( .A(n40609), .Z(n40606) );
  HS65_LH_BFX2 U24903 ( .A(n40611), .Z(n40607) );
  HS65_LH_IVX2 U24904 ( .A(n40722), .Z(n40608) );
  HS65_LH_IVX2 U24905 ( .A(n40608), .Z(n40609) );
  HS65_LH_IVX2 U24906 ( .A(n40716), .Z(n40610) );
  HS65_LH_IVX2 U24907 ( .A(n40610), .Z(n40611) );
  HS65_LH_BFX2 U24908 ( .A(n40613), .Z(n40612) );
  HS65_LH_BFX2 U24909 ( .A(n40614), .Z(n40613) );
  HS65_LH_BFX2 U24910 ( .A(n40714), .Z(n40614) );
  HS65_LH_BFX2 U24911 ( .A(n40616), .Z(n40615) );
  HS65_LH_BFX2 U24912 ( .A(n40617), .Z(n40616) );
  HS65_LH_BFX2 U24913 ( .A(n40618), .Z(n40617) );
  HS65_LH_BFX2 U24914 ( .A(n40619), .Z(n40618) );
  HS65_LH_BFX2 U24915 ( .A(n40620), .Z(n40619) );
  HS65_LH_BFX2 U24916 ( .A(n40621), .Z(n40620) );
  HS65_LH_BFX2 U24917 ( .A(n40622), .Z(n40621) );
  HS65_LH_BFX2 U24918 ( .A(n40623), .Z(n40622) );
  HS65_LH_BFX2 U24919 ( .A(n40624), .Z(n40623) );
  HS65_LH_BFX2 U24920 ( .A(n40625), .Z(n40624) );
  HS65_LH_BFX2 U24921 ( .A(n40626), .Z(n40625) );
  HS65_LH_BFX2 U24922 ( .A(n40627), .Z(n40626) );
  HS65_LH_BFX2 U24923 ( .A(n40628), .Z(n40627) );
  HS65_LH_BFX2 U24924 ( .A(n40629), .Z(n40628) );
  HS65_LH_BFX2 U24925 ( .A(n17625), .Z(n40629) );
  HS65_LH_BFX2 U24926 ( .A(n40631), .Z(n40630) );
  HS65_LH_BFX2 U24927 ( .A(n40632), .Z(n40631) );
  HS65_LH_BFX2 U24928 ( .A(n40633), .Z(n40632) );
  HS65_LH_BFX2 U24929 ( .A(n40634), .Z(n40633) );
  HS65_LH_BFX2 U24930 ( .A(n40635), .Z(n40634) );
  HS65_LH_BFX2 U24931 ( .A(n40636), .Z(n40635) );
  HS65_LH_BFX2 U24932 ( .A(n40637), .Z(n40636) );
  HS65_LH_BFX2 U24933 ( .A(n40638), .Z(n40637) );
  HS65_LH_BFX2 U24934 ( .A(n40639), .Z(n40638) );
  HS65_LH_BFX2 U24936 ( .A(n40640), .Z(n40639) );
  HS65_LH_BFX2 U24937 ( .A(n40641), .Z(n40640) );
  HS65_LH_BFX2 U24938 ( .A(n40642), .Z(n40641) );
  HS65_LH_BFX2 U24939 ( .A(n40643), .Z(n40642) );
  HS65_LH_BFX2 U24940 ( .A(n40644), .Z(n40643) );
  HS65_LH_BFX2 U24941 ( .A(n40645), .Z(n40644) );
  HS65_LH_BFX2 U24942 ( .A(n40646), .Z(n40645) );
  HS65_LH_BFX2 U24943 ( .A(n40647), .Z(n40646) );
  HS65_LH_BFX2 U24944 ( .A(n40648), .Z(n40647) );
  HS65_LH_BFX2 U24945 ( .A(n40649), .Z(n40648) );
  HS65_LH_BFX2 U24946 ( .A(n14656), .Z(n40649) );
  HS65_LH_BFX2 U24947 ( .A(n40651), .Z(n40650) );
  HS65_LH_BFX2 U24948 ( .A(n17589), .Z(n40651) );
  HS65_LH_BFX2 U24949 ( .A(n40655), .Z(n40652) );
  HS65_LH_BFX2 U24950 ( .A(n40656), .Z(n40653) );
  HS65_LH_BFX2 U24951 ( .A(n17779), .Z(n40654) );
  HS65_LH_BFX2 U24952 ( .A(n40658), .Z(n40655) );
  HS65_LH_BFX2 U24953 ( .A(n40659), .Z(n40656) );
  HS65_LH_BFX2 U24954 ( .A(n40654), .Z(n40657) );
  HS65_LH_BFX2 U24955 ( .A(n40661), .Z(n40658) );
  HS65_LH_BFX2 U24956 ( .A(n40662), .Z(n40659) );
  HS65_LH_BFX2 U24957 ( .A(n40657), .Z(n40660) );
  HS65_LH_BFX2 U24958 ( .A(n40664), .Z(n40661) );
  HS65_LH_BFX2 U24959 ( .A(n40665), .Z(n40662) );
  HS65_LH_BFX2 U24960 ( .A(n40660), .Z(n40663) );
  HS65_LH_BFX2 U24961 ( .A(n40667), .Z(n40664) );
  HS65_LH_BFX2 U24962 ( .A(n40668), .Z(n40665) );
  HS65_LH_BFX2 U24963 ( .A(n40663), .Z(n40666) );
  HS65_LH_BFX2 U24964 ( .A(n40670), .Z(n40667) );
  HS65_LH_BFX2 U24965 ( .A(n40671), .Z(n40668) );
  HS65_LH_BFX2 U24966 ( .A(n40666), .Z(n40669) );
  HS65_LH_BFX2 U24967 ( .A(n40673), .Z(n40670) );
  HS65_LH_BFX2 U24968 ( .A(n40674), .Z(n40671) );
  HS65_LH_BFX2 U24969 ( .A(n40669), .Z(n40672) );
  HS65_LH_BFX2 U24970 ( .A(n40676), .Z(n40673) );
  HS65_LH_BFX2 U24971 ( .A(n40677), .Z(n40674) );
  HS65_LH_BFX2 U24972 ( .A(n40672), .Z(n40675) );
  HS65_LH_BFX2 U24973 ( .A(n40679), .Z(n40676) );
  HS65_LH_BFX2 U24974 ( .A(n40680), .Z(n40677) );
  HS65_LH_BFX2 U24975 ( .A(n40675), .Z(n40678) );
  HS65_LH_BFX2 U24976 ( .A(n40682), .Z(n40679) );
  HS65_LH_BFX2 U24977 ( .A(n40683), .Z(n40680) );
  HS65_LH_BFX2 U24978 ( .A(n40678), .Z(n40681) );
  HS65_LH_BFX2 U24979 ( .A(n40685), .Z(n40682) );
  HS65_LH_BFX2 U24980 ( .A(n40686), .Z(n40683) );
  HS65_LH_BFX2 U24981 ( .A(n40681), .Z(n40684) );
  HS65_LH_BFX2 U24982 ( .A(n40688), .Z(n40685) );
  HS65_LH_BFX2 U24983 ( .A(n40689), .Z(n40686) );
  HS65_LH_BFX2 U24984 ( .A(n40684), .Z(n40687) );
  HS65_LH_BFX2 U24985 ( .A(n40691), .Z(n40688) );
  HS65_LH_BFX2 U24986 ( .A(n40692), .Z(n40689) );
  HS65_LH_BFX2 U24987 ( .A(n40687), .Z(n40690) );
  HS65_LH_BFX2 U24988 ( .A(n40694), .Z(n40691) );
  HS65_LH_BFX2 U24989 ( .A(n40695), .Z(n40692) );
  HS65_LH_BFX2 U24990 ( .A(n40690), .Z(n40693) );
  HS65_LH_BFX2 U24991 ( .A(n40697), .Z(n40694) );
  HS65_LH_BFX2 U24992 ( .A(n40698), .Z(n40695) );
  HS65_LH_BFX2 U24993 ( .A(n40693), .Z(n40696) );
  HS65_LH_BFX2 U24994 ( .A(n40700), .Z(n40697) );
  HS65_LH_BFX2 U24995 ( .A(n40701), .Z(n40698) );
  HS65_LH_BFX2 U24996 ( .A(n40696), .Z(n40699) );
  HS65_LH_BFX2 U24997 ( .A(n40703), .Z(n40700) );
  HS65_LH_BFX2 U24998 ( .A(n40704), .Z(n40701) );
  HS65_LH_BFX2 U24999 ( .A(n40699), .Z(n40702) );
  HS65_LH_BFX2 U25000 ( .A(n40706), .Z(n40703) );
  HS65_LH_BFX2 U25001 ( .A(n40707), .Z(n40704) );
  HS65_LH_BFX2 U25002 ( .A(n40702), .Z(n40705) );
  HS65_LH_BFX2 U25003 ( .A(n17754), .Z(n40706) );
  HS65_LH_BFX2 U25004 ( .A(n40710), .Z(n40707) );
  HS65_LH_BFX2 U25005 ( .A(n40705), .Z(n40708) );
  HS65_LH_IVX2 U25006 ( .A(n17877), .Z(n40709) );
  HS65_LH_IVX2 U25007 ( .A(n40709), .Z(n40710) );
  HS65_LH_IVX2 U25008 ( .A(n40708), .Z(n40711) );
  HS65_LH_IVX2 U25009 ( .A(n40711), .Z(n40712) );
  HS65_LH_BFX2 U25010 ( .A(n40719), .Z(n40713) );
  HS65_LH_BFX2 U25011 ( .A(n40720), .Z(n40714) );
  HS65_LH_BFX2 U25012 ( .A(n40721), .Z(n40715) );
  HS65_LH_BFX2 U25013 ( .A(n40723), .Z(n40716) );
  HS65_LH_BFX2 U25014 ( .A(n40724), .Z(n40717) );
  HS65_LH_BFX2 U25015 ( .A(n40725), .Z(n40718) );
  HS65_LH_BFX2 U25016 ( .A(n40726), .Z(n40719) );
  HS65_LH_BFX2 U25017 ( .A(n40727), .Z(n40720) );
  HS65_LH_BFX2 U25018 ( .A(n40728), .Z(n40721) );
  HS65_LH_BFX2 U25019 ( .A(n40729), .Z(n40722) );
  HS65_LH_BFX2 U25020 ( .A(n40730), .Z(n40723) );
  HS65_LH_BFX2 U25021 ( .A(n40731), .Z(n40724) );
  HS65_LH_BFX2 U25022 ( .A(n40732), .Z(n40725) );
  HS65_LH_BFX2 U25023 ( .A(n40733), .Z(n40726) );
  HS65_LH_BFX2 U25024 ( .A(n40734), .Z(n40727) );
  HS65_LH_BFX2 U25025 ( .A(n40735), .Z(n40728) );
  HS65_LH_BFX2 U25026 ( .A(n40736), .Z(n40729) );
  HS65_LH_BFX2 U25027 ( .A(n40737), .Z(n40730) );
  HS65_LH_BFX2 U25028 ( .A(n40738), .Z(n40731) );
  HS65_LH_BFX2 U25029 ( .A(n40739), .Z(n40732) );
  HS65_LH_BFX2 U25030 ( .A(n40740), .Z(n40733) );
  HS65_LH_BFX2 U25031 ( .A(n40741), .Z(n40734) );
  HS65_LH_BFX2 U25032 ( .A(n40742), .Z(n40735) );
  HS65_LH_BFX2 U25033 ( .A(n40743), .Z(n40736) );
  HS65_LH_BFX2 U25034 ( .A(n40744), .Z(n40737) );
  HS65_LH_BFX2 U25035 ( .A(n40745), .Z(n40738) );
  HS65_LH_BFX2 U25036 ( .A(n40746), .Z(n40739) );
  HS65_LH_BFX2 U25037 ( .A(n40747), .Z(n40740) );
  HS65_LH_BFX2 U25038 ( .A(n40748), .Z(n40741) );
  HS65_LH_BFX2 U25039 ( .A(n40749), .Z(n40742) );
  HS65_LH_BFX2 U25040 ( .A(n40750), .Z(n40743) );
  HS65_LH_BFX2 U25041 ( .A(n40751), .Z(n40744) );
  HS65_LH_BFX2 U25042 ( .A(n40752), .Z(n40745) );
  HS65_LH_BFX2 U25043 ( .A(n40753), .Z(n40746) );
  HS65_LH_BFX2 U25044 ( .A(n40754), .Z(n40747) );
  HS65_LH_BFX2 U25045 ( .A(n40755), .Z(n40748) );
  HS65_LH_BFX2 U25046 ( .A(n40756), .Z(n40749) );
  HS65_LH_BFX2 U25047 ( .A(n40757), .Z(n40750) );
  HS65_LH_BFX2 U25048 ( .A(n40758), .Z(n40751) );
  HS65_LH_BFX2 U25049 ( .A(n40759), .Z(n40752) );
  HS65_LH_BFX2 U25050 ( .A(n40760), .Z(n40753) );
  HS65_LH_BFX2 U25051 ( .A(n40761), .Z(n40754) );
  HS65_LH_BFX2 U25052 ( .A(n40762), .Z(n40755) );
  HS65_LH_BFX2 U25053 ( .A(n40763), .Z(n40756) );
  HS65_LH_BFX2 U25054 ( .A(n40764), .Z(n40757) );
  HS65_LH_BFX2 U25055 ( .A(n40765), .Z(n40758) );
  HS65_LH_BFX2 U25056 ( .A(n40766), .Z(n40759) );
  HS65_LH_BFX2 U25057 ( .A(n40767), .Z(n40760) );
  HS65_LH_BFX2 U25058 ( .A(n40768), .Z(n40761) );
  HS65_LH_BFX2 U25059 ( .A(n40769), .Z(n40762) );
  HS65_LH_BFX2 U25060 ( .A(n40770), .Z(n40763) );
  HS65_LH_BFX2 U25061 ( .A(n40771), .Z(n40764) );
  HS65_LH_BFX2 U25062 ( .A(n40772), .Z(n40765) );
  HS65_LH_BFX2 U25063 ( .A(n40773), .Z(n40766) );
  HS65_LH_BFX2 U25064 ( .A(n40774), .Z(n40767) );
  HS65_LH_BFX2 U25065 ( .A(n40775), .Z(n40768) );
  HS65_LH_BFX2 U25066 ( .A(n40776), .Z(n40769) );
  HS65_LH_BFX2 U25067 ( .A(n40777), .Z(n40770) );
  HS65_LH_BFX2 U25068 ( .A(n40778), .Z(n40771) );
  HS65_LH_BFX2 U25069 ( .A(n40779), .Z(n40772) );
  HS65_LH_BFX2 U25070 ( .A(n40780), .Z(n40773) );
  HS65_LH_BFX2 U25071 ( .A(n40781), .Z(n40774) );
  HS65_LH_BFX2 U25072 ( .A(n40782), .Z(n40775) );
  HS65_LH_BFX2 U25073 ( .A(n40783), .Z(n40776) );
  HS65_LH_BFX2 U25074 ( .A(n40784), .Z(n40777) );
  HS65_LH_BFX2 U25075 ( .A(n40785), .Z(n40778) );
  HS65_LH_BFX2 U25076 ( .A(n40786), .Z(n40779) );
  HS65_LH_BFX2 U25077 ( .A(n40787), .Z(n40780) );
  HS65_LH_BFX2 U25078 ( .A(n40788), .Z(n40781) );
  HS65_LH_BFX2 U25079 ( .A(n40789), .Z(n40782) );
  HS65_LH_BFX2 U25080 ( .A(n40790), .Z(n40783) );
  HS65_LH_BFX2 U25081 ( .A(n40791), .Z(n40784) );
  HS65_LH_BFX2 U25082 ( .A(n40792), .Z(n40785) );
  HS65_LH_BFX2 U25083 ( .A(n40793), .Z(n40786) );
  HS65_LH_BFX2 U25084 ( .A(n40794), .Z(n40787) );
  HS65_LH_BFX2 U25085 ( .A(n40795), .Z(n40788) );
  HS65_LH_BFX2 U25086 ( .A(n40796), .Z(n40789) );
  HS65_LH_BFX2 U25087 ( .A(n40797), .Z(n40790) );
  HS65_LH_BFX2 U25088 ( .A(n40798), .Z(n40791) );
  HS65_LH_BFX2 U25089 ( .A(n40799), .Z(n40792) );
  HS65_LH_BFX2 U25090 ( .A(n40800), .Z(n40793) );
  HS65_LH_BFX2 U25091 ( .A(n40801), .Z(n40794) );
  HS65_LH_BFX2 U25092 ( .A(n40802), .Z(n40795) );
  HS65_LH_BFX2 U25093 ( .A(n40803), .Z(n40796) );
  HS65_LH_BFX2 U25094 ( .A(n40804), .Z(n40797) );
  HS65_LH_BFX2 U25095 ( .A(n40805), .Z(n40798) );
  HS65_LH_BFX2 U25096 ( .A(n40806), .Z(n40799) );
  HS65_LH_BFX2 U25097 ( .A(n40807), .Z(n40800) );
  HS65_LH_BFX2 U25098 ( .A(n40808), .Z(n40801) );
  HS65_LH_BFX2 U25099 ( .A(n40809), .Z(n40802) );
  HS65_LH_BFX2 U25100 ( .A(n40810), .Z(n40803) );
  HS65_LH_BFX2 U25101 ( .A(n40811), .Z(n40804) );
  HS65_LH_BFX2 U25102 ( .A(n40812), .Z(n40805) );
  HS65_LH_BFX2 U25103 ( .A(n40813), .Z(n40806) );
  HS65_LH_BFX2 U25104 ( .A(n40814), .Z(n40807) );
  HS65_LH_BFX2 U25105 ( .A(n40815), .Z(n40808) );
  HS65_LH_BFX2 U25106 ( .A(n40816), .Z(n40809) );
  HS65_LH_BFX2 U25107 ( .A(n40817), .Z(n40810) );
  HS65_LH_BFX2 U25108 ( .A(n40818), .Z(n40811) );
  HS65_LH_BFX2 U25109 ( .A(n40819), .Z(n40812) );
  HS65_LH_BFX2 U25110 ( .A(n40820), .Z(n40813) );
  HS65_LH_BFX2 U25111 ( .A(n40821), .Z(n40814) );
  HS65_LH_BFX2 U25112 ( .A(n40822), .Z(n40815) );
  HS65_LH_BFX2 U25113 ( .A(n40823), .Z(n40816) );
  HS65_LH_BFX2 U25114 ( .A(n40824), .Z(n40817) );
  HS65_LH_BFX2 U25115 ( .A(n40825), .Z(n40818) );
  HS65_LH_BFX2 U25116 ( .A(n40826), .Z(n40819) );
  HS65_LH_BFX2 U25117 ( .A(n40827), .Z(n40820) );
  HS65_LH_BFX2 U25118 ( .A(n40828), .Z(n40821) );
  HS65_LH_BFX2 U25119 ( .A(n40831), .Z(n40822) );
  HS65_LH_BFX2 U25120 ( .A(n40832), .Z(n40823) );
  HS65_LH_BFX2 U25121 ( .A(n40833), .Z(n40824) );
  HS65_LH_BFX2 U25122 ( .A(n17836), .Z(n40825) );
  HS65_LH_BFX2 U25123 ( .A(n40830), .Z(n40826) );
  HS65_LH_BFX2 U25124 ( .A(n40834), .Z(n40827) );
  HS65_LH_BFX2 U25125 ( .A(n40835), .Z(n40828) );
  HS65_LH_IVX2 U25126 ( .A(n17833), .Z(n40829) );
  HS65_LH_IVX2 U25127 ( .A(n40829), .Z(n40830) );
  HS65_LH_BFX2 U25128 ( .A(n40836), .Z(n40831) );
  HS65_LH_BFX2 U25129 ( .A(n40837), .Z(n40832) );
  HS65_LH_BFX2 U25130 ( .A(n40838), .Z(n40833) );
  HS65_LH_BFX2 U25131 ( .A(n17846), .Z(n40834) );
  HS65_LH_BFX2 U25132 ( .A(n17842), .Z(n40835) );
  HS65_LH_BFX2 U25133 ( .A(n17839), .Z(n40836) );
  HS65_LH_BFX2 U25134 ( .A(n40839), .Z(n40837) );
  HS65_LH_BFX2 U25135 ( .A(n17793), .Z(n40838) );
  HS65_LH_BFX2 U25136 ( .A(n17753), .Z(n40839) );
  HS65_LH_BFX2 U25137 ( .A(n40842), .Z(n40840) );
  HS65_LH_IVX2 U25138 ( .A(n40843), .Z(n40841) );
  HS65_LH_IVX2 U25139 ( .A(n40841), .Z(n40842) );
  HS65_LH_BFX2 U25140 ( .A(n40844), .Z(n40843) );
  HS65_LH_BFX2 U25141 ( .A(n40845), .Z(n40844) );
  HS65_LH_BFX2 U25142 ( .A(n40846), .Z(n40845) );
  HS65_LH_BFX2 U25143 ( .A(n40847), .Z(n40846) );
  HS65_LH_BFX2 U25144 ( .A(n40848), .Z(n40847) );
  HS65_LH_BFX2 U25145 ( .A(n40849), .Z(n40848) );
  HS65_LH_BFX2 U25146 ( .A(n40850), .Z(n40849) );
  HS65_LH_BFX2 U25147 ( .A(n40851), .Z(n40850) );
  HS65_LH_BFX2 U25148 ( .A(n40852), .Z(n40851) );
  HS65_LH_BFX2 U25149 ( .A(n40853), .Z(n40852) );
  HS65_LH_BFX2 U25150 ( .A(n40854), .Z(n40853) );
  HS65_LH_BFX2 U25151 ( .A(n40855), .Z(n40854) );
  HS65_LH_BFX2 U25152 ( .A(n40856), .Z(n40855) );
  HS65_LH_BFX2 U25153 ( .A(n40857), .Z(n40856) );
  HS65_LH_BFX2 U25154 ( .A(n40858), .Z(n40857) );
  HS65_LH_BFX2 U25155 ( .A(n40859), .Z(n40858) );
  HS65_LH_BFX2 U25156 ( .A(n40860), .Z(n40859) );
  HS65_LH_BFX2 U25157 ( .A(n40861), .Z(n40860) );
  HS65_LH_BFX2 U25158 ( .A(n14510), .Z(n40861) );
  HS65_LH_BFX2 U25159 ( .A(n40863), .Z(n40862) );
  HS65_LH_BFX2 U25160 ( .A(n40864), .Z(n40863) );
  HS65_LH_BFX2 U25161 ( .A(n40865), .Z(n40864) );
  HS65_LH_BFX2 U25162 ( .A(n40866), .Z(n40865) );
  HS65_LH_BFX2 U25163 ( .A(n40867), .Z(n40866) );
  HS65_LH_BFX2 U25164 ( .A(n40868), .Z(n40867) );
  HS65_LH_BFX2 U25165 ( .A(n40869), .Z(n40868) );
  HS65_LH_BFX2 U25166 ( .A(n40870), .Z(n40869) );
  HS65_LH_BFX2 U25167 ( .A(n40871), .Z(n40870) );
  HS65_LH_BFX2 U25168 ( .A(n40872), .Z(n40871) );
  HS65_LH_BFX2 U25169 ( .A(n40873), .Z(n40872) );
  HS65_LH_BFX2 U25170 ( .A(n40874), .Z(n40873) );
  HS65_LH_BFX2 U25171 ( .A(n40875), .Z(n40874) );
  HS65_LH_BFX2 U25172 ( .A(n40876), .Z(n40875) );
  HS65_LH_BFX2 U25173 ( .A(n40877), .Z(n40876) );
  HS65_LH_BFX2 U25174 ( .A(n40878), .Z(n40877) );
  HS65_LH_BFX2 U25175 ( .A(n40879), .Z(n40878) );
  HS65_LH_BFX2 U25176 ( .A(n40880), .Z(n40879) );
  HS65_LH_BFX2 U25177 ( .A(n40881), .Z(n40880) );
  HS65_LH_BFX2 U25178 ( .A(n17600), .Z(n40881) );
  HS65_LH_BFX2 U25179 ( .A(n40885), .Z(n40882) );
  HS65_LH_BFX2 U25180 ( .A(n40888), .Z(n40883) );
  HS65_LH_IVX2 U25181 ( .A(n40892), .Z(n40884) );
  HS65_LH_IVX2 U25182 ( .A(n40884), .Z(n40885) );
  HS65_LH_BFX2 U25183 ( .A(n1150), .Z(n40886) );
  HS65_LH_IVX2 U25184 ( .A(n40897), .Z(n40887) );
  HS65_LH_IVX2 U25185 ( .A(n40887), .Z(n40888) );
  HS65_LH_BFX2 U25186 ( .A(n40907), .Z(n40889) );
  HS65_LH_BFX2 U25187 ( .A(n40886), .Z(n40890) );
  HS65_LH_IVX2 U25188 ( .A(n40900), .Z(n40891) );
  HS65_LH_IVX2 U25189 ( .A(n40891), .Z(n40892) );
  HS65_LH_BFX2 U25190 ( .A(n40986), .Z(n40893) );
  HS65_LH_IVX2 U25191 ( .A(n40902), .Z(n40894) );
  HS65_LH_IVX2 U25192 ( .A(n40894), .Z(n40895) );
  HS65_LH_IVX2 U25193 ( .A(n40904), .Z(n40896) );
  HS65_LH_IVX2 U25194 ( .A(n40896), .Z(n40897) );
  HS65_LH_BFX2 U25195 ( .A(n40893), .Z(n40898) );
  HS65_LH_IVX2 U25196 ( .A(n40909), .Z(n40899) );
  HS65_LH_IVX2 U25197 ( .A(n40899), .Z(n40900) );
  HS65_LH_IVX2 U25198 ( .A(n40911), .Z(n40901) );
  HS65_LH_IVX2 U25199 ( .A(n40901), .Z(n40902) );
  HS65_LH_IVX2 U25200 ( .A(n40913), .Z(n40903) );
  HS65_LH_IVX2 U25201 ( .A(n40903), .Z(n40904) );
  HS65_LH_BFX2 U25202 ( .A(n40898), .Z(n40905) );
  HS65_LH_IVX2 U25203 ( .A(n40915), .Z(n40906) );
  HS65_LH_IVX2 U25204 ( .A(n40906), .Z(n40907) );
  HS65_LH_IVX2 U25205 ( .A(n40917), .Z(n40908) );
  HS65_LH_IVX2 U25206 ( .A(n40908), .Z(n40909) );
  HS65_LH_IVX2 U25207 ( .A(n40919), .Z(n40910) );
  HS65_LH_IVX2 U25208 ( .A(n40910), .Z(n40911) );
  HS65_LH_IVX2 U25209 ( .A(n40921), .Z(n40912) );
  HS65_LH_IVX2 U25210 ( .A(n40912), .Z(n40913) );
  HS65_LH_IVX2 U25211 ( .A(n40923), .Z(n40914) );
  HS65_LH_IVX2 U25212 ( .A(n40914), .Z(n40915) );
  HS65_LH_IVX2 U25213 ( .A(n40925), .Z(n40916) );
  HS65_LH_IVX2 U25214 ( .A(n40916), .Z(n40917) );
  HS65_LH_IVX2 U25215 ( .A(n40927), .Z(n40918) );
  HS65_LH_IVX2 U25216 ( .A(n40918), .Z(n40919) );
  HS65_LH_IVX2 U25217 ( .A(n40929), .Z(n40920) );
  HS65_LH_IVX2 U25218 ( .A(n40920), .Z(n40921) );
  HS65_LH_IVX2 U25219 ( .A(n40936), .Z(n40922) );
  HS65_LH_IVX2 U25220 ( .A(n40922), .Z(n40923) );
  HS65_LH_IVX2 U25221 ( .A(n40931), .Z(n40924) );
  HS65_LH_IVX2 U25222 ( .A(n40924), .Z(n40925) );
  HS65_LH_IVX2 U25223 ( .A(n40933), .Z(n40926) );
  HS65_LH_IVX2 U25224 ( .A(n40926), .Z(n40927) );
  HS65_LH_IVX2 U25225 ( .A(n40935), .Z(n40928) );
  HS65_LH_IVX2 U25226 ( .A(n40928), .Z(n40929) );
  HS65_LH_IVX2 U25227 ( .A(n40938), .Z(n40930) );
  HS65_LH_IVX2 U25228 ( .A(n40930), .Z(n40931) );
  HS65_LH_IVX2 U25229 ( .A(n40940), .Z(n40932) );
  HS65_LH_IVX2 U25230 ( .A(n40932), .Z(n40933) );
  HS65_LH_IVX2 U25231 ( .A(n40942), .Z(n40934) );
  HS65_LH_IVX2 U25232 ( .A(n40934), .Z(n40935) );
  HS65_LH_BFX2 U25234 ( .A(n40943), .Z(n40936) );
  HS65_LH_IVX2 U25235 ( .A(n40945), .Z(n40937) );
  HS65_LH_IVX2 U25236 ( .A(n40937), .Z(n40938) );
  HS65_LH_IVX2 U25237 ( .A(n40947), .Z(n40939) );
  HS65_LH_IVX2 U25238 ( .A(n40939), .Z(n40940) );
  HS65_LH_IVX2 U25239 ( .A(n40949), .Z(n40941) );
  HS65_LH_IVX2 U25240 ( .A(n40941), .Z(n40942) );
  HS65_LH_BFX2 U25242 ( .A(n40950), .Z(n40943) );
  HS65_LH_IVX2 U25243 ( .A(n40952), .Z(n40944) );
  HS65_LH_IVX2 U25244 ( .A(n40944), .Z(n40945) );
  HS65_LH_IVX2 U25245 ( .A(n40954), .Z(n40946) );
  HS65_LH_IVX2 U25246 ( .A(n40946), .Z(n40947) );
  HS65_LH_IVX2 U25248 ( .A(n40956), .Z(n40948) );
  HS65_LH_IVX2 U25251 ( .A(n40948), .Z(n40949) );
  HS65_LH_BFX2 U25252 ( .A(n40957), .Z(n40950) );
  HS65_LH_IVX2 U25253 ( .A(n40959), .Z(n40951) );
  HS65_LH_IVX2 U25254 ( .A(n40951), .Z(n40952) );
  HS65_LH_IVX2 U25255 ( .A(n40961), .Z(n40953) );
  HS65_LH_IVX2 U25256 ( .A(n40953), .Z(n40954) );
  HS65_LH_IVX2 U25257 ( .A(n40963), .Z(n40955) );
  HS65_LH_IVX2 U25259 ( .A(n40955), .Z(n40956) );
  HS65_LH_BFX2 U25260 ( .A(n21117), .Z(n40957) );
  HS65_LH_IVX2 U25261 ( .A(n40968), .Z(n40958) );
  HS65_LH_IVX2 U25262 ( .A(n40958), .Z(n40959) );
  HS65_LH_IVX2 U25263 ( .A(n40965), .Z(n40960) );
  HS65_LH_IVX2 U25264 ( .A(n40960), .Z(n40961) );
  HS65_LH_IVX2 U25265 ( .A(n40967), .Z(n40962) );
  HS65_LH_IVX2 U25266 ( .A(n40962), .Z(n40963) );
  HS65_LH_IVX2 U25267 ( .A(n40970), .Z(n40964) );
  HS65_LH_IVX2 U25268 ( .A(n40964), .Z(n40965) );
  HS65_LH_IVX2 U25269 ( .A(n40972), .Z(n40966) );
  HS65_LH_IVX2 U25270 ( .A(n40966), .Z(n40967) );
  HS65_LH_BFX2 U25271 ( .A(n40973), .Z(n40968) );
  HS65_LH_IVX2 U25272 ( .A(n40980), .Z(n40969) );
  HS65_LH_IVX2 U25273 ( .A(n40969), .Z(n40970) );
  HS65_LH_IVX2 U25274 ( .A(n40975), .Z(n40971) );
  HS65_LH_IVX2 U25275 ( .A(n40971), .Z(n40972) );
  HS65_LH_BFX2 U25276 ( .A(n40977), .Z(n40973) );
  HS65_LH_IVX2 U25277 ( .A(n1151), .Z(n40974) );
  HS65_LH_IVX2 U25278 ( .A(n40974), .Z(n40975) );
  HS65_LH_BFX2 U25279 ( .A(n17168), .Z(n40976) );
  HS65_LH_BFX2 U25280 ( .A(n40979), .Z(n40977) );
  HS65_LH_IVX2 U25281 ( .A(n40981), .Z(n40978) );
  HS65_LH_IVX2 U25282 ( .A(n40978), .Z(n40979) );
  HS65_LH_BFX2 U25283 ( .A(n40890), .Z(n40980) );
  HS65_LH_BFX2 U25284 ( .A(n40982), .Z(n40981) );
  HS65_LH_BFX2 U25285 ( .A(n40983), .Z(n40982) );
  HS65_LH_BFX2 U25286 ( .A(n40984), .Z(n40983) );
  HS65_LH_BFX2 U25287 ( .A(n17845), .Z(n40984) );
  HS65_LH_IVX18 U25288 ( .A(n17489), .Z(n29653) );
  HS65_LH_IVX18 U25289 ( .A(n18140), .Z(n29655) );
  HS65_LH_IVX18 U25290 ( .A(n18141), .Z(n29657) );
  HS65_LH_IVX18 U25291 ( .A(n18142), .Z(n29659) );
  HS65_LH_IVX18 U25292 ( .A(n18143), .Z(n29661) );
  HS65_LH_IVX18 U25293 ( .A(n18144), .Z(n29663) );
  HS65_LH_IVX18 U25294 ( .A(n18145), .Z(n29665) );
  HS65_LH_IVX18 U25295 ( .A(n18146), .Z(n29667) );
  HS65_LH_IVX18 U25296 ( .A(n18132), .Z(n29669) );
  HS65_LH_IVX18 U25297 ( .A(n18135), .Z(n29671) );
  HS65_LH_IVX18 U25298 ( .A(n17459), .Z(n29673) );
  HS65_LH_IVX18 U25299 ( .A(n18133), .Z(n29675) );
  HS65_LH_IVX18 U25300 ( .A(n18128), .Z(n29677) );
  HS65_LH_IVX18 U25301 ( .A(n18129), .Z(n29679) );
  HS65_LH_IVX18 U25302 ( .A(n18134), .Z(n29681) );
  HS65_LH_IVX18 U25303 ( .A(n18130), .Z(n29683) );
  HS65_LH_IVX18 U25304 ( .A(n18131), .Z(n29685) );
  HS65_LH_IVX18 U25305 ( .A(n17490), .Z(n29687) );
  HS65_LH_IVX18 U25306 ( .A(n17627), .Z(n29689) );
  HS65_LH_MUXI21X5 U25307 ( .D0(n32068), .D1(n17609), .S0(n17528), .Z(n15341)
         );
  HS65_LH_IVX18 U25308 ( .A(n40999), .Z(n29694) );
  HS65_LH_IVX9 U25309 ( .A(n14218), .Z(n14226) );
  HS65_LH_OAI212X3 U25310 ( .A(n17480), .B(n17698), .C(n17613), .D(n17586), 
        .E(n15175), .Z(n40986) );
  HS65_LH_AOI22X1 U25311 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][17] ), .B(n17121), .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][17] ), .D(n17403), 
        .Z(n40987) );
  HS65_LH_AOI22X1 U25312 ( .A(n17420), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][31] ), .C(n16446), 
        .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][31] ), .Z(
        n40988) );
  HS65_LH_NAND2X2 U25313 ( .A(n16674), .B(n16673), .Z(n40989) );
  HS65_LH_AOI21X2 U25314 ( .A(n15754), .B(n37070), .C(n24656), .Z(n40990) );
  HS65_LH_AOI21X2 U25315 ( .A(n17305), .B(n17446), .C(n17267), .Z(n40991) );
  HS65_LH_BFX2 U25316 ( .A(n17410), .Z(n40993) );
  HS65_LH_BFX2 U25317 ( .A(n17408), .Z(n40994) );
  HS65_LH_BFX2 U25318 ( .A(n17417), .Z(n40995) );
  HS65_LH_NOR2X5 U25319 ( .A(n15341), .B(n15500), .Z(n14218) );
  HS65_LH_IVX2 U25320 ( .A(n17245), .Z(n40996) );
  HS65_LH_IVX2 U25321 ( .A(n40996), .Z(n40997) );
  HS65_LH_IVX2 U25322 ( .A(n40996), .Z(n40998) );
  HS65_LH_IVX2 U25323 ( .A(n40996), .Z(n40999) );
  HS65_LH_IVX2 U25324 ( .A(n40996), .Z(n41000) );
  HS65_LH_IVX4 U25325 ( .A(n29694), .Z(n29651) );
endmodule

