--------------------------------------------------------------------------------
-- Decode Unit
-- This unit implements the decode unit. Sub-units which are contained are:
--  - Hazard Detection Unit
--   - Register File
--  - Sign-Extension
--  - Extender
--  - Mux Stall
--------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use work.globals.all;

--------------------------------------------------------------------------------
--------------------------------------------------------------------------------

entity decode_unit is
  port (
    -- INPUTS
    address_write          : in std_logic_vector(4 downto 0);                         -- register address that should be written
    data_write             : in std_logic_vector(31 downto 0);                        -- data to be written in the reg file
    pc_4_from_dec          : in std_logic_vector(31 downto 0);                        -- Program counter incremented by 4
    instruction            : in std_logic_vector(31 downto 0);                        -- instruction fetched
    idex_rt                : in std_logic_vector(4 downto 0);                         -- Rt register coming from the ex stage
    clk                    : in std_logic;                                            -- global clock
    rst                    : in std_logic;                                            -- global reset signal
    reg_write              : in std_logic;                                            -- Reg Write signal to enable the write operation
    idex_mem_read          : in std_logic_vector(3 downto 0);                         -- control signals for Mem Read (lb,lhu, lw, lbu)
    cw                     : in std_logic_vector((CW_SIZE+ALUOP_SIZE)-1 downto 0);    -- control word + alu operation produced by the CU
    -- OUTPUTS
    cw_to_ex               : out std_logic_vector((CW_SIZE+ALUOP_SIZE)-2 downto 0);   -- control word + alu operation for the ex stage (-2 since unsigned control signal used i the decode stage)
    jump_address           : out std_logic_vector(31 downto 0);                       -- jump address sign-extended
    pc_4_to_ex             : out std_logic_vector(31 downto 0);                       -- Program counter incremented by 4 directed to the ex stage
    data_read_1            : out std_logic_vector(31 downto 0);                       -- Output of read port 1 of reg file
    data_read_2            : out std_logic_vector(31 downto 0);                       -- Output of read port 2 of reg file
    immediate_ext          : out std_logic_vector(31 downto 0);                       -- Immediate field signe-exntended
    immediate              : out std_logic_vector(15 downto 0);                       -- Immediate filed not sign extended (for LUI instruction)
    rt                     : out std_logic_Vector(4 downto 0);                        -- rt address (instruction 20-16)
    rd                     : out std_logic_vector(4 downto 0);                        -- rd address (instruction 15-11)
    rs                     : out std_logic_vector(4 downto 0);                        -- rs address (instruction 25-21)
    opcode                 : out std_logic_vector(OPCODE_SIZE-1 downto 0);            -- opcode for the CU, instruction (31-26)
    func                   : out std_logic_vector(FUNC_SIZE-1 downto 0);              -- func field of instruction (10-0) to the CU
    pcwrite                : out std_logic;                                           -- write enable generated by the Hazard Detection Unit for the PC
    ifid_write             : out std_logic                                            -- write enable generated by the Hazard Detection Unit for the IF/ID pipeline register
    );
end decode_unit;


--------------------------------------------------------------------------------
--------------------------------------------------------------------------------

architecture structural of decode_unit is

-- Component Declarations
component reg_file is
  port (
    -- INPUTS
    read_address_1   : in std_logic_vector(4 downto 0);   -- address of reg 1 to be read(instruction 25-21)
    read_address_2   : in std_logic_vector(4 downto 0);   -- address of reg 2 to be read(instruction 20-16)
    write_address    : in std_logic_vector(4 downto 0);   -- address of reg to be written
    write_data       : in std_logic_vector(31 downto 0);  -- data to be written at the address specified in wirte_address
    reg_write        : in std_logic;
    rst              : in std_logic;
    -- OUTPUTS
    data_reg_1       : out std_logic_vector(31 downto 0);  -- data from read port 1
    data_reg_2       : out std_logic_vector(31 downto 0)   -- data from read port 2
    );
end component;


component extender is
  port (
    -- INPUTS
    immediate      : in std_logic_vector(15 downto 0);    -- immediate filed (instruction 15 -0)
    unsigned_value : in std_logic;                        -- control signal generated by the CU
    -- OUTPUTS
    extended       : out std_logic_vector(31 downto 0)    -- extended value
    );
end component;


component sign_extender is
  port (
    -- INPUTS
    immediate_jump   : in std_logic_vector(25 downto 0);  -- instructon (25-0)
    -- OUTPUTS
    extended_jump    : out std_logic_vector(31 downto 0)  -- sign-extended jump immediate
    );
end component;

component mux_stall is
  port (
    -- INPUTS
    cw_from_cu    : in std_logic_vector((CW_SIZE + ALUOP_SIZE)-1 downto 0);      -- control word produced by the CU
    mux_op        : in std_logic;                                                -- control signal produced by the hazard detection unit
    -- OUTPUTS
    cw_from_mux   : out std_logic_vector((CW_SIZE+ALUOP_SIZE)-1 downto 0)        -- control word produced by the mux
    );
end component;


component hdu is
  port (
    -- INPUTS
    clk             : in std_logic;                           -- global clock signal
    rst             : in std_logic;                           -- global reset signal
    idex_mem_read   : in std_logic_vector(3 downto 0);        -- ID/EX MemRead control signals (lbu, lw, lhu, lb)
    idex_rt         : in std_logic_vector(4 downto 0);        -- ID/EX Rt address
    rs              : in std_logic_vector(4 downto 0);        -- Rs address instruction (25-21)
    rt              : in std_logic_vector(4 downto 0);        -- Rt address instruction (20-16)
    -- OUTPUTS
    pcwrite         : out std_logic;                          -- control signal write enable for the PC register
    ifidwrite       : out std_logic;                          -- control signal write enable for the pipeline register IF/ID
    mux_op          : out std_logic                           -- control signal directed to the mux stall
    );
end component;

-- Internal Signals
signal unsigned_value_i  : std_logic;
signal cw_i              : std_logic_vector((CW_SIZE+ALUOP_SIZE)-1 downto 0);
signal mux_op_i          : std_logic;

begin

  -- Cuncurrent statements

  -- Extract from the control word the unsigned control signal and re-arrenge the Cw itself
  cw_to_ex           <= cw_i((CW_SIZE+ALUOP_SIZE)-1) & cw_i((CW_SIZE+ALUOP_SIZE)-3 downto 0);
  unsigned_value_i   <= cw_i((CW_SIZE+ALUOP_SIZE)-2);

  -- Output assignmet
  opcode       <= instruction(31 downto 26);
  func         <= instruction(10 downto 0);
  pc_4_to_ex   <= pc_4_from_dec;
  immediate    <= instruction(15 downto 0);
  rt           <= instruction(20 downto 16);
  rd           <= instruction(15 downto 11);
  rs           <= instruction(25 downto 21);

  -- Components instantiation
  hdu_0: hdu port map (
        clk             => clk,
        rst             => rst,
        idex_mem_read   => idex_mem_read,
        idex_rt         => idex_rt,
        rs              => instruction(25 downto 21),
        rt              => instruction(20 downto 16),
        pcwrite         => pcwrite,
        ifidwrite       => ifid_write,
        mux_op          => mux_op_i
        );

  mux_stall0: mux_stall port map(
          cw_from_cu    => cw,
          mux_op        => mux_op_i,
          cw_from_mux   => cw_i
          );

  sign_extender0: sign_extender port map(
            immediate_jump => instruction(25 downto 0),
            extended_jump  => jump_address
            );

  extender0: extender port map (
          immediate       => instruction(15 downto 0),
          unsigned_value  => unsigned_value_i,
          extended        => immediate_ext
          );

  reg_file0: reg_file port map (
          read_address_1   => instruction(25 downto 21),
          read_address_2   => instruction(20 downto 16),
          write_address    => address_write,
          write_data       => data_write,
          reg_write        => reg_write,
          rst              => rst,
          data_reg_1       => data_read_1,
          data_reg_2       => data_read_2
          );




end structural;
